module basic_500_3000_500_3_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_273,In_206);
nand U1 (N_1,In_87,In_484);
nand U2 (N_2,In_132,In_18);
nand U3 (N_3,In_212,In_51);
and U4 (N_4,In_357,In_328);
and U5 (N_5,In_445,In_78);
and U6 (N_6,In_415,In_184);
or U7 (N_7,In_83,In_279);
nand U8 (N_8,In_320,In_193);
or U9 (N_9,In_53,In_365);
and U10 (N_10,In_351,In_135);
and U11 (N_11,In_225,In_61);
and U12 (N_12,In_466,In_438);
xor U13 (N_13,In_324,In_491);
or U14 (N_14,In_75,In_158);
xnor U15 (N_15,In_182,In_373);
or U16 (N_16,In_290,In_370);
xor U17 (N_17,In_272,In_405);
nand U18 (N_18,In_67,In_307);
and U19 (N_19,In_34,In_82);
xnor U20 (N_20,In_6,In_3);
xnor U21 (N_21,In_295,In_248);
nand U22 (N_22,In_462,In_460);
or U23 (N_23,In_452,In_44);
nor U24 (N_24,In_123,In_227);
nor U25 (N_25,In_162,In_362);
or U26 (N_26,In_113,In_404);
nand U27 (N_27,In_38,In_299);
or U28 (N_28,In_15,In_310);
nand U29 (N_29,In_104,In_128);
and U30 (N_30,In_375,In_169);
xnor U31 (N_31,In_165,In_497);
xor U32 (N_32,In_60,In_24);
or U33 (N_33,In_140,In_309);
nand U34 (N_34,In_346,In_489);
xnor U35 (N_35,In_455,In_122);
and U36 (N_36,In_407,In_349);
or U37 (N_37,In_444,In_447);
nand U38 (N_38,In_190,In_396);
nand U39 (N_39,In_347,In_402);
nand U40 (N_40,In_353,In_474);
or U41 (N_41,In_263,In_427);
and U42 (N_42,In_418,In_383);
or U43 (N_43,In_26,In_260);
or U44 (N_44,In_208,In_361);
or U45 (N_45,In_437,In_251);
nand U46 (N_46,In_339,In_315);
and U47 (N_47,In_245,In_194);
nor U48 (N_48,In_145,In_183);
xnor U49 (N_49,In_33,In_226);
nand U50 (N_50,In_237,In_12);
or U51 (N_51,In_446,In_468);
xnor U52 (N_52,In_48,In_35);
or U53 (N_53,In_143,In_285);
and U54 (N_54,In_72,In_178);
and U55 (N_55,In_477,In_413);
or U56 (N_56,In_441,In_392);
and U57 (N_57,In_327,In_464);
and U58 (N_58,In_220,In_216);
nor U59 (N_59,In_68,In_157);
nand U60 (N_60,In_319,In_287);
and U61 (N_61,In_175,In_229);
nor U62 (N_62,In_329,In_449);
nand U63 (N_63,In_435,In_210);
or U64 (N_64,In_440,In_160);
xor U65 (N_65,In_282,In_298);
xnor U66 (N_66,In_79,In_371);
or U67 (N_67,In_63,In_431);
nor U68 (N_68,In_207,In_28);
nor U69 (N_69,In_341,In_246);
xnor U70 (N_70,In_55,In_19);
or U71 (N_71,In_163,In_377);
nor U72 (N_72,In_267,In_133);
or U73 (N_73,In_231,In_101);
nor U74 (N_74,In_265,In_81);
nand U75 (N_75,In_335,In_17);
nor U76 (N_76,In_120,In_368);
and U77 (N_77,In_271,In_420);
nor U78 (N_78,In_98,In_172);
or U79 (N_79,In_149,In_49);
nor U80 (N_80,In_451,In_280);
nand U81 (N_81,In_344,In_322);
or U82 (N_82,In_269,In_209);
or U83 (N_83,In_25,In_180);
or U84 (N_84,In_286,In_323);
and U85 (N_85,In_142,In_257);
or U86 (N_86,In_302,In_264);
and U87 (N_87,In_16,In_196);
nor U88 (N_88,In_36,In_458);
nor U89 (N_89,In_105,In_480);
xor U90 (N_90,In_116,In_54);
and U91 (N_91,In_150,In_296);
and U92 (N_92,In_117,In_159);
xor U93 (N_93,In_359,In_41);
nand U94 (N_94,In_469,In_52);
and U95 (N_95,In_258,In_125);
xor U96 (N_96,In_121,In_381);
or U97 (N_97,In_379,In_382);
nand U98 (N_98,In_131,In_270);
nor U99 (N_99,In_336,In_367);
xnor U100 (N_100,In_118,In_201);
or U101 (N_101,In_119,In_65);
and U102 (N_102,In_204,In_40);
and U103 (N_103,In_283,In_86);
xor U104 (N_104,In_337,In_102);
and U105 (N_105,In_23,In_84);
and U106 (N_106,In_443,In_192);
xnor U107 (N_107,In_199,In_250);
and U108 (N_108,In_423,In_403);
nand U109 (N_109,In_168,In_334);
or U110 (N_110,In_228,In_454);
and U111 (N_111,In_151,In_369);
xnor U112 (N_112,In_64,In_235);
nand U113 (N_113,In_146,In_74);
nand U114 (N_114,In_316,In_236);
or U115 (N_115,In_358,In_218);
or U116 (N_116,In_90,In_417);
and U117 (N_117,In_30,In_0);
xor U118 (N_118,In_161,In_170);
xor U119 (N_119,In_380,In_166);
nand U120 (N_120,In_37,In_378);
nand U121 (N_121,In_171,In_490);
nor U122 (N_122,In_400,In_342);
and U123 (N_123,In_465,In_495);
nor U124 (N_124,In_253,In_385);
and U125 (N_125,In_191,In_202);
or U126 (N_126,In_434,In_419);
nand U127 (N_127,In_111,In_356);
or U128 (N_128,In_97,In_92);
xnor U129 (N_129,In_408,In_252);
nor U130 (N_130,In_56,In_412);
and U131 (N_131,In_69,In_401);
nor U132 (N_132,In_376,In_360);
and U133 (N_133,In_5,In_481);
or U134 (N_134,In_141,In_390);
xnor U135 (N_135,In_42,In_374);
nand U136 (N_136,In_148,In_115);
or U137 (N_137,In_313,In_200);
xor U138 (N_138,In_453,In_241);
nor U139 (N_139,In_487,In_494);
xor U140 (N_140,In_106,In_303);
nor U141 (N_141,In_174,In_177);
xnor U142 (N_142,In_234,In_467);
and U143 (N_143,In_372,In_486);
nor U144 (N_144,In_317,In_197);
or U145 (N_145,In_305,In_22);
and U146 (N_146,In_364,In_99);
xor U147 (N_147,In_66,In_232);
nor U148 (N_148,In_21,In_278);
and U149 (N_149,In_31,In_259);
nand U150 (N_150,In_243,In_11);
nor U151 (N_151,In_397,In_414);
nor U152 (N_152,In_155,In_488);
and U153 (N_153,In_139,In_409);
nand U154 (N_154,In_219,In_185);
and U155 (N_155,In_222,In_448);
or U156 (N_156,In_406,In_43);
xor U157 (N_157,In_103,In_181);
and U158 (N_158,In_95,In_483);
xnor U159 (N_159,In_217,In_492);
and U160 (N_160,In_325,In_77);
nor U161 (N_161,In_1,In_136);
nor U162 (N_162,In_421,In_108);
nor U163 (N_163,In_152,In_274);
nor U164 (N_164,In_138,In_312);
nand U165 (N_165,In_112,In_398);
and U166 (N_166,In_354,In_70);
and U167 (N_167,In_189,In_58);
or U168 (N_168,In_13,In_126);
nand U169 (N_169,In_442,In_333);
nand U170 (N_170,In_110,In_129);
or U171 (N_171,In_297,In_394);
and U172 (N_172,In_188,In_304);
nor U173 (N_173,In_153,In_88);
nand U174 (N_174,In_355,In_473);
nand U175 (N_175,In_345,In_255);
and U176 (N_176,In_164,In_485);
nor U177 (N_177,In_395,In_284);
or U178 (N_178,In_130,In_478);
or U179 (N_179,In_173,In_433);
nor U180 (N_180,In_213,In_456);
xnor U181 (N_181,In_156,In_463);
xor U182 (N_182,In_91,In_50);
nor U183 (N_183,In_47,In_27);
or U184 (N_184,In_124,In_71);
or U185 (N_185,In_144,In_242);
and U186 (N_186,In_186,In_176);
nor U187 (N_187,In_73,In_247);
and U188 (N_188,In_471,In_428);
or U189 (N_189,In_80,In_343);
nor U190 (N_190,In_389,In_100);
nand U191 (N_191,In_300,In_308);
nand U192 (N_192,In_340,In_20);
nor U193 (N_193,In_425,In_457);
xnor U194 (N_194,In_230,In_472);
nand U195 (N_195,In_461,In_107);
or U196 (N_196,In_261,In_14);
nor U197 (N_197,In_256,In_85);
and U198 (N_198,In_432,In_332);
or U199 (N_199,In_59,In_391);
xor U200 (N_200,In_89,In_393);
nor U201 (N_201,In_331,In_294);
nor U202 (N_202,In_76,In_238);
xor U203 (N_203,In_8,In_496);
nand U204 (N_204,In_326,In_45);
nand U205 (N_205,In_470,In_187);
xor U206 (N_206,In_223,In_224);
and U207 (N_207,In_276,In_4);
nor U208 (N_208,In_482,In_262);
nand U209 (N_209,In_9,In_363);
and U210 (N_210,In_277,In_147);
and U211 (N_211,In_288,In_399);
nor U212 (N_212,In_93,In_211);
xnor U213 (N_213,In_7,In_475);
and U214 (N_214,In_94,In_459);
nand U215 (N_215,In_289,In_429);
or U216 (N_216,In_114,In_62);
nand U217 (N_217,In_411,In_293);
and U218 (N_218,In_127,In_306);
nand U219 (N_219,In_249,In_318);
nor U220 (N_220,In_281,In_424);
xnor U221 (N_221,In_350,In_314);
nand U222 (N_222,In_439,In_410);
nand U223 (N_223,In_254,In_215);
xor U224 (N_224,In_426,In_436);
and U225 (N_225,In_57,In_321);
nand U226 (N_226,In_291,In_195);
or U227 (N_227,In_244,In_137);
and U228 (N_228,In_198,In_266);
xor U229 (N_229,In_338,In_301);
and U230 (N_230,In_388,In_352);
xnor U231 (N_231,In_476,In_416);
nand U232 (N_232,In_450,In_330);
nor U233 (N_233,In_10,In_134);
or U234 (N_234,In_240,In_214);
or U235 (N_235,In_2,In_29);
or U236 (N_236,In_39,In_239);
or U237 (N_237,In_96,In_479);
and U238 (N_238,In_233,In_221);
or U239 (N_239,In_498,In_292);
and U240 (N_240,In_109,In_422);
and U241 (N_241,In_366,In_32);
nand U242 (N_242,In_205,In_167);
nor U243 (N_243,In_311,In_348);
and U244 (N_244,In_387,In_268);
nor U245 (N_245,In_386,In_275);
and U246 (N_246,In_179,In_493);
nor U247 (N_247,In_499,In_46);
xnor U248 (N_248,In_430,In_384);
and U249 (N_249,In_154,In_203);
nor U250 (N_250,In_458,In_61);
nand U251 (N_251,In_182,In_45);
nand U252 (N_252,In_397,In_130);
nand U253 (N_253,In_34,In_472);
and U254 (N_254,In_468,In_301);
nor U255 (N_255,In_164,In_295);
nand U256 (N_256,In_242,In_383);
and U257 (N_257,In_317,In_281);
and U258 (N_258,In_256,In_372);
or U259 (N_259,In_174,In_349);
xor U260 (N_260,In_234,In_55);
and U261 (N_261,In_117,In_424);
xnor U262 (N_262,In_218,In_397);
or U263 (N_263,In_47,In_89);
or U264 (N_264,In_217,In_348);
nor U265 (N_265,In_497,In_380);
and U266 (N_266,In_130,In_324);
xor U267 (N_267,In_10,In_149);
nand U268 (N_268,In_334,In_213);
xor U269 (N_269,In_76,In_28);
and U270 (N_270,In_313,In_407);
nor U271 (N_271,In_450,In_219);
xor U272 (N_272,In_431,In_249);
xnor U273 (N_273,In_213,In_132);
nand U274 (N_274,In_80,In_13);
or U275 (N_275,In_340,In_466);
xnor U276 (N_276,In_101,In_225);
and U277 (N_277,In_339,In_121);
nor U278 (N_278,In_114,In_370);
nand U279 (N_279,In_238,In_467);
nand U280 (N_280,In_351,In_387);
nor U281 (N_281,In_323,In_300);
and U282 (N_282,In_148,In_450);
and U283 (N_283,In_161,In_147);
and U284 (N_284,In_25,In_372);
or U285 (N_285,In_108,In_167);
xor U286 (N_286,In_202,In_479);
xor U287 (N_287,In_70,In_38);
nor U288 (N_288,In_276,In_243);
xnor U289 (N_289,In_499,In_266);
xnor U290 (N_290,In_220,In_472);
nor U291 (N_291,In_34,In_150);
and U292 (N_292,In_465,In_356);
xnor U293 (N_293,In_371,In_372);
xnor U294 (N_294,In_72,In_27);
xnor U295 (N_295,In_483,In_305);
nand U296 (N_296,In_351,In_315);
and U297 (N_297,In_409,In_94);
nor U298 (N_298,In_65,In_290);
xor U299 (N_299,In_27,In_103);
nand U300 (N_300,In_463,In_159);
or U301 (N_301,In_350,In_166);
nand U302 (N_302,In_21,In_292);
xnor U303 (N_303,In_228,In_248);
nand U304 (N_304,In_240,In_187);
xnor U305 (N_305,In_39,In_190);
xnor U306 (N_306,In_152,In_463);
or U307 (N_307,In_216,In_55);
nand U308 (N_308,In_291,In_473);
or U309 (N_309,In_424,In_377);
or U310 (N_310,In_366,In_114);
or U311 (N_311,In_51,In_223);
xor U312 (N_312,In_66,In_249);
xor U313 (N_313,In_127,In_359);
nor U314 (N_314,In_442,In_399);
nor U315 (N_315,In_278,In_257);
or U316 (N_316,In_23,In_56);
or U317 (N_317,In_499,In_131);
nor U318 (N_318,In_415,In_103);
or U319 (N_319,In_402,In_322);
nor U320 (N_320,In_144,In_11);
nor U321 (N_321,In_94,In_327);
or U322 (N_322,In_471,In_236);
nor U323 (N_323,In_232,In_325);
nand U324 (N_324,In_147,In_95);
or U325 (N_325,In_383,In_271);
nor U326 (N_326,In_30,In_67);
xor U327 (N_327,In_282,In_214);
and U328 (N_328,In_334,In_283);
nand U329 (N_329,In_249,In_10);
and U330 (N_330,In_440,In_251);
or U331 (N_331,In_286,In_460);
xor U332 (N_332,In_484,In_156);
or U333 (N_333,In_214,In_441);
nand U334 (N_334,In_297,In_290);
nor U335 (N_335,In_447,In_94);
nor U336 (N_336,In_286,In_357);
and U337 (N_337,In_441,In_191);
nor U338 (N_338,In_364,In_348);
xor U339 (N_339,In_67,In_383);
nor U340 (N_340,In_375,In_237);
xor U341 (N_341,In_145,In_141);
and U342 (N_342,In_254,In_157);
and U343 (N_343,In_25,In_352);
xnor U344 (N_344,In_137,In_363);
and U345 (N_345,In_255,In_109);
or U346 (N_346,In_212,In_149);
nand U347 (N_347,In_497,In_292);
or U348 (N_348,In_148,In_262);
nand U349 (N_349,In_480,In_117);
or U350 (N_350,In_362,In_325);
nor U351 (N_351,In_107,In_469);
or U352 (N_352,In_396,In_18);
xor U353 (N_353,In_130,In_301);
and U354 (N_354,In_408,In_304);
nand U355 (N_355,In_49,In_350);
or U356 (N_356,In_127,In_351);
nor U357 (N_357,In_382,In_190);
nor U358 (N_358,In_494,In_143);
or U359 (N_359,In_349,In_262);
or U360 (N_360,In_150,In_429);
nand U361 (N_361,In_209,In_17);
or U362 (N_362,In_477,In_452);
and U363 (N_363,In_111,In_26);
nand U364 (N_364,In_354,In_458);
or U365 (N_365,In_428,In_258);
or U366 (N_366,In_275,In_277);
nand U367 (N_367,In_69,In_218);
xor U368 (N_368,In_78,In_154);
and U369 (N_369,In_452,In_227);
or U370 (N_370,In_313,In_213);
and U371 (N_371,In_109,In_214);
and U372 (N_372,In_441,In_315);
nand U373 (N_373,In_117,In_324);
nor U374 (N_374,In_427,In_391);
xor U375 (N_375,In_317,In_375);
nor U376 (N_376,In_272,In_341);
nand U377 (N_377,In_423,In_28);
xor U378 (N_378,In_64,In_54);
and U379 (N_379,In_110,In_441);
xnor U380 (N_380,In_231,In_106);
or U381 (N_381,In_27,In_145);
and U382 (N_382,In_357,In_352);
nor U383 (N_383,In_458,In_83);
nand U384 (N_384,In_322,In_25);
xnor U385 (N_385,In_24,In_102);
and U386 (N_386,In_269,In_127);
or U387 (N_387,In_329,In_498);
nor U388 (N_388,In_0,In_434);
nor U389 (N_389,In_286,In_224);
or U390 (N_390,In_316,In_286);
xor U391 (N_391,In_455,In_266);
nor U392 (N_392,In_82,In_134);
and U393 (N_393,In_440,In_282);
and U394 (N_394,In_215,In_29);
nor U395 (N_395,In_459,In_323);
and U396 (N_396,In_114,In_308);
nor U397 (N_397,In_71,In_144);
nor U398 (N_398,In_76,In_346);
xnor U399 (N_399,In_148,In_390);
or U400 (N_400,In_267,In_132);
or U401 (N_401,In_199,In_467);
and U402 (N_402,In_324,In_327);
and U403 (N_403,In_256,In_150);
nand U404 (N_404,In_44,In_429);
xnor U405 (N_405,In_86,In_231);
xor U406 (N_406,In_427,In_416);
or U407 (N_407,In_281,In_270);
or U408 (N_408,In_495,In_202);
and U409 (N_409,In_135,In_339);
or U410 (N_410,In_324,In_497);
xnor U411 (N_411,In_338,In_169);
nor U412 (N_412,In_90,In_43);
nor U413 (N_413,In_256,In_140);
or U414 (N_414,In_288,In_403);
nor U415 (N_415,In_350,In_57);
xnor U416 (N_416,In_460,In_390);
xor U417 (N_417,In_97,In_446);
and U418 (N_418,In_488,In_234);
nand U419 (N_419,In_223,In_370);
xor U420 (N_420,In_281,In_77);
nand U421 (N_421,In_406,In_245);
nor U422 (N_422,In_260,In_318);
or U423 (N_423,In_376,In_318);
nor U424 (N_424,In_434,In_354);
or U425 (N_425,In_73,In_314);
nand U426 (N_426,In_259,In_427);
nand U427 (N_427,In_465,In_27);
nand U428 (N_428,In_332,In_169);
or U429 (N_429,In_253,In_278);
or U430 (N_430,In_402,In_204);
xor U431 (N_431,In_467,In_339);
xor U432 (N_432,In_455,In_250);
nor U433 (N_433,In_494,In_373);
or U434 (N_434,In_276,In_138);
nor U435 (N_435,In_67,In_304);
or U436 (N_436,In_65,In_71);
or U437 (N_437,In_367,In_490);
nand U438 (N_438,In_60,In_150);
nor U439 (N_439,In_142,In_253);
nand U440 (N_440,In_477,In_327);
nor U441 (N_441,In_100,In_331);
nand U442 (N_442,In_384,In_276);
nand U443 (N_443,In_151,In_426);
or U444 (N_444,In_27,In_116);
xnor U445 (N_445,In_229,In_15);
xor U446 (N_446,In_124,In_111);
xnor U447 (N_447,In_264,In_361);
xor U448 (N_448,In_153,In_298);
nand U449 (N_449,In_347,In_204);
or U450 (N_450,In_2,In_341);
and U451 (N_451,In_286,In_137);
xnor U452 (N_452,In_392,In_292);
and U453 (N_453,In_350,In_35);
xnor U454 (N_454,In_0,In_215);
nand U455 (N_455,In_422,In_91);
xnor U456 (N_456,In_350,In_393);
or U457 (N_457,In_483,In_492);
or U458 (N_458,In_232,In_130);
nand U459 (N_459,In_383,In_54);
and U460 (N_460,In_282,In_202);
nor U461 (N_461,In_218,In_142);
nand U462 (N_462,In_8,In_375);
nor U463 (N_463,In_138,In_149);
nor U464 (N_464,In_230,In_388);
nand U465 (N_465,In_1,In_490);
xor U466 (N_466,In_108,In_74);
nor U467 (N_467,In_75,In_281);
nor U468 (N_468,In_408,In_211);
nor U469 (N_469,In_228,In_40);
and U470 (N_470,In_400,In_242);
nand U471 (N_471,In_19,In_229);
xnor U472 (N_472,In_229,In_319);
nor U473 (N_473,In_203,In_200);
nand U474 (N_474,In_34,In_387);
xnor U475 (N_475,In_397,In_323);
nor U476 (N_476,In_291,In_125);
nand U477 (N_477,In_188,In_463);
or U478 (N_478,In_356,In_181);
xor U479 (N_479,In_103,In_78);
and U480 (N_480,In_117,In_376);
nor U481 (N_481,In_326,In_24);
nand U482 (N_482,In_92,In_31);
xor U483 (N_483,In_9,In_137);
xor U484 (N_484,In_154,In_290);
xnor U485 (N_485,In_260,In_334);
and U486 (N_486,In_427,In_405);
xor U487 (N_487,In_70,In_464);
nand U488 (N_488,In_488,In_151);
or U489 (N_489,In_368,In_461);
nand U490 (N_490,In_122,In_357);
nand U491 (N_491,In_62,In_146);
nor U492 (N_492,In_175,In_402);
and U493 (N_493,In_168,In_335);
nand U494 (N_494,In_286,In_354);
nand U495 (N_495,In_188,In_402);
nand U496 (N_496,In_8,In_428);
xnor U497 (N_497,In_101,In_191);
or U498 (N_498,In_26,In_421);
and U499 (N_499,In_208,In_459);
nor U500 (N_500,In_255,In_269);
or U501 (N_501,In_58,In_195);
and U502 (N_502,In_124,In_338);
and U503 (N_503,In_98,In_185);
nor U504 (N_504,In_418,In_335);
and U505 (N_505,In_224,In_212);
nand U506 (N_506,In_334,In_296);
or U507 (N_507,In_416,In_72);
nand U508 (N_508,In_159,In_292);
or U509 (N_509,In_199,In_427);
and U510 (N_510,In_247,In_310);
or U511 (N_511,In_347,In_261);
and U512 (N_512,In_73,In_174);
or U513 (N_513,In_27,In_401);
xor U514 (N_514,In_278,In_231);
nor U515 (N_515,In_104,In_26);
and U516 (N_516,In_217,In_391);
nor U517 (N_517,In_144,In_305);
or U518 (N_518,In_443,In_6);
and U519 (N_519,In_158,In_119);
or U520 (N_520,In_449,In_334);
nand U521 (N_521,In_215,In_453);
and U522 (N_522,In_443,In_277);
and U523 (N_523,In_113,In_308);
xnor U524 (N_524,In_277,In_314);
xor U525 (N_525,In_393,In_41);
or U526 (N_526,In_188,In_439);
nor U527 (N_527,In_199,In_70);
nand U528 (N_528,In_479,In_197);
xnor U529 (N_529,In_470,In_14);
and U530 (N_530,In_237,In_64);
nor U531 (N_531,In_107,In_225);
nand U532 (N_532,In_244,In_94);
or U533 (N_533,In_146,In_186);
nand U534 (N_534,In_359,In_268);
xor U535 (N_535,In_373,In_376);
nor U536 (N_536,In_234,In_228);
nor U537 (N_537,In_465,In_6);
and U538 (N_538,In_249,In_305);
or U539 (N_539,In_493,In_264);
and U540 (N_540,In_67,In_487);
or U541 (N_541,In_450,In_122);
and U542 (N_542,In_324,In_45);
and U543 (N_543,In_452,In_141);
and U544 (N_544,In_330,In_426);
and U545 (N_545,In_157,In_173);
xor U546 (N_546,In_248,In_272);
and U547 (N_547,In_276,In_385);
and U548 (N_548,In_461,In_283);
nor U549 (N_549,In_135,In_300);
or U550 (N_550,In_230,In_315);
nor U551 (N_551,In_121,In_379);
xnor U552 (N_552,In_196,In_8);
and U553 (N_553,In_428,In_3);
nand U554 (N_554,In_25,In_48);
xnor U555 (N_555,In_293,In_326);
and U556 (N_556,In_170,In_23);
and U557 (N_557,In_344,In_40);
nand U558 (N_558,In_225,In_252);
nor U559 (N_559,In_375,In_234);
and U560 (N_560,In_141,In_427);
or U561 (N_561,In_334,In_219);
xnor U562 (N_562,In_109,In_348);
xor U563 (N_563,In_157,In_134);
and U564 (N_564,In_170,In_402);
nand U565 (N_565,In_237,In_177);
and U566 (N_566,In_145,In_438);
xor U567 (N_567,In_398,In_423);
and U568 (N_568,In_296,In_241);
nor U569 (N_569,In_46,In_297);
and U570 (N_570,In_123,In_365);
nor U571 (N_571,In_252,In_77);
nand U572 (N_572,In_380,In_381);
or U573 (N_573,In_338,In_112);
nand U574 (N_574,In_491,In_86);
nand U575 (N_575,In_322,In_491);
xnor U576 (N_576,In_426,In_371);
and U577 (N_577,In_258,In_36);
xor U578 (N_578,In_234,In_74);
or U579 (N_579,In_448,In_163);
nand U580 (N_580,In_324,In_67);
xnor U581 (N_581,In_18,In_127);
nor U582 (N_582,In_76,In_498);
or U583 (N_583,In_111,In_224);
xnor U584 (N_584,In_67,In_342);
nor U585 (N_585,In_448,In_78);
or U586 (N_586,In_495,In_75);
or U587 (N_587,In_414,In_140);
or U588 (N_588,In_496,In_365);
nor U589 (N_589,In_0,In_196);
and U590 (N_590,In_394,In_449);
nand U591 (N_591,In_114,In_22);
or U592 (N_592,In_66,In_465);
and U593 (N_593,In_51,In_105);
nor U594 (N_594,In_183,In_467);
nor U595 (N_595,In_170,In_39);
or U596 (N_596,In_298,In_10);
or U597 (N_597,In_314,In_51);
or U598 (N_598,In_196,In_350);
or U599 (N_599,In_345,In_18);
and U600 (N_600,In_82,In_259);
and U601 (N_601,In_191,In_367);
nor U602 (N_602,In_175,In_202);
or U603 (N_603,In_382,In_54);
and U604 (N_604,In_73,In_220);
and U605 (N_605,In_28,In_201);
nand U606 (N_606,In_373,In_157);
and U607 (N_607,In_415,In_292);
or U608 (N_608,In_295,In_242);
or U609 (N_609,In_105,In_415);
and U610 (N_610,In_186,In_286);
or U611 (N_611,In_376,In_363);
nor U612 (N_612,In_261,In_265);
nor U613 (N_613,In_301,In_494);
and U614 (N_614,In_384,In_299);
and U615 (N_615,In_401,In_441);
and U616 (N_616,In_423,In_466);
and U617 (N_617,In_240,In_110);
nor U618 (N_618,In_440,In_352);
nand U619 (N_619,In_248,In_58);
nand U620 (N_620,In_433,In_298);
nand U621 (N_621,In_471,In_481);
nand U622 (N_622,In_358,In_200);
or U623 (N_623,In_240,In_400);
nor U624 (N_624,In_309,In_341);
nor U625 (N_625,In_441,In_102);
nor U626 (N_626,In_241,In_416);
and U627 (N_627,In_14,In_116);
nand U628 (N_628,In_355,In_369);
nand U629 (N_629,In_216,In_127);
or U630 (N_630,In_178,In_286);
nor U631 (N_631,In_443,In_362);
nand U632 (N_632,In_363,In_473);
nand U633 (N_633,In_441,In_370);
nor U634 (N_634,In_453,In_82);
nor U635 (N_635,In_423,In_81);
nor U636 (N_636,In_417,In_229);
nor U637 (N_637,In_477,In_16);
nand U638 (N_638,In_71,In_132);
and U639 (N_639,In_231,In_219);
or U640 (N_640,In_239,In_281);
or U641 (N_641,In_312,In_404);
nor U642 (N_642,In_468,In_109);
xnor U643 (N_643,In_44,In_438);
nand U644 (N_644,In_174,In_118);
xnor U645 (N_645,In_51,In_268);
nor U646 (N_646,In_344,In_239);
nor U647 (N_647,In_7,In_237);
nand U648 (N_648,In_210,In_473);
and U649 (N_649,In_357,In_3);
or U650 (N_650,In_368,In_489);
xor U651 (N_651,In_157,In_191);
nor U652 (N_652,In_287,In_443);
nor U653 (N_653,In_51,In_118);
and U654 (N_654,In_444,In_411);
xor U655 (N_655,In_158,In_243);
xnor U656 (N_656,In_105,In_222);
nand U657 (N_657,In_209,In_454);
and U658 (N_658,In_497,In_5);
nor U659 (N_659,In_234,In_240);
nand U660 (N_660,In_223,In_470);
and U661 (N_661,In_87,In_123);
and U662 (N_662,In_381,In_365);
and U663 (N_663,In_144,In_207);
or U664 (N_664,In_297,In_72);
and U665 (N_665,In_134,In_17);
or U666 (N_666,In_72,In_475);
xnor U667 (N_667,In_61,In_377);
and U668 (N_668,In_472,In_479);
or U669 (N_669,In_163,In_105);
or U670 (N_670,In_184,In_249);
nor U671 (N_671,In_223,In_290);
nor U672 (N_672,In_19,In_310);
or U673 (N_673,In_483,In_422);
nand U674 (N_674,In_463,In_441);
xnor U675 (N_675,In_29,In_390);
and U676 (N_676,In_272,In_251);
nor U677 (N_677,In_365,In_357);
xnor U678 (N_678,In_299,In_262);
and U679 (N_679,In_106,In_305);
nor U680 (N_680,In_221,In_242);
nand U681 (N_681,In_404,In_328);
xnor U682 (N_682,In_154,In_271);
nor U683 (N_683,In_433,In_148);
and U684 (N_684,In_195,In_200);
or U685 (N_685,In_464,In_359);
and U686 (N_686,In_339,In_421);
and U687 (N_687,In_323,In_60);
or U688 (N_688,In_231,In_58);
xnor U689 (N_689,In_446,In_284);
nand U690 (N_690,In_332,In_207);
and U691 (N_691,In_127,In_145);
xnor U692 (N_692,In_144,In_313);
or U693 (N_693,In_413,In_52);
or U694 (N_694,In_96,In_480);
xor U695 (N_695,In_328,In_158);
nand U696 (N_696,In_465,In_72);
or U697 (N_697,In_92,In_379);
and U698 (N_698,In_8,In_429);
xnor U699 (N_699,In_148,In_472);
nand U700 (N_700,In_37,In_178);
xor U701 (N_701,In_453,In_221);
nor U702 (N_702,In_419,In_128);
xnor U703 (N_703,In_491,In_194);
and U704 (N_704,In_339,In_272);
or U705 (N_705,In_163,In_98);
nor U706 (N_706,In_26,In_171);
nor U707 (N_707,In_337,In_219);
and U708 (N_708,In_331,In_265);
or U709 (N_709,In_116,In_287);
nand U710 (N_710,In_77,In_328);
nand U711 (N_711,In_24,In_142);
xnor U712 (N_712,In_350,In_342);
and U713 (N_713,In_137,In_153);
and U714 (N_714,In_111,In_395);
xnor U715 (N_715,In_366,In_414);
xor U716 (N_716,In_17,In_475);
and U717 (N_717,In_374,In_307);
nand U718 (N_718,In_440,In_78);
or U719 (N_719,In_205,In_380);
nor U720 (N_720,In_27,In_44);
xor U721 (N_721,In_21,In_497);
xnor U722 (N_722,In_488,In_168);
nor U723 (N_723,In_115,In_488);
xor U724 (N_724,In_418,In_389);
nor U725 (N_725,In_32,In_320);
nand U726 (N_726,In_144,In_223);
nor U727 (N_727,In_317,In_0);
or U728 (N_728,In_353,In_144);
or U729 (N_729,In_230,In_349);
and U730 (N_730,In_432,In_228);
xnor U731 (N_731,In_53,In_454);
and U732 (N_732,In_300,In_0);
nor U733 (N_733,In_315,In_0);
nor U734 (N_734,In_310,In_381);
nand U735 (N_735,In_69,In_369);
and U736 (N_736,In_201,In_356);
or U737 (N_737,In_131,In_464);
or U738 (N_738,In_37,In_157);
xnor U739 (N_739,In_312,In_155);
nand U740 (N_740,In_240,In_45);
nand U741 (N_741,In_201,In_419);
xnor U742 (N_742,In_240,In_58);
nand U743 (N_743,In_352,In_312);
and U744 (N_744,In_6,In_234);
nand U745 (N_745,In_329,In_14);
nor U746 (N_746,In_81,In_394);
or U747 (N_747,In_173,In_440);
nor U748 (N_748,In_152,In_273);
and U749 (N_749,In_59,In_111);
xnor U750 (N_750,In_355,In_50);
xnor U751 (N_751,In_426,In_255);
xor U752 (N_752,In_154,In_305);
xor U753 (N_753,In_256,In_105);
or U754 (N_754,In_413,In_67);
or U755 (N_755,In_90,In_58);
nand U756 (N_756,In_76,In_264);
nor U757 (N_757,In_469,In_352);
nor U758 (N_758,In_253,In_99);
or U759 (N_759,In_237,In_65);
nor U760 (N_760,In_270,In_205);
nor U761 (N_761,In_476,In_301);
and U762 (N_762,In_240,In_303);
and U763 (N_763,In_449,In_84);
or U764 (N_764,In_375,In_413);
xnor U765 (N_765,In_48,In_108);
xor U766 (N_766,In_127,In_38);
and U767 (N_767,In_379,In_261);
nor U768 (N_768,In_41,In_277);
nand U769 (N_769,In_349,In_290);
xor U770 (N_770,In_342,In_185);
nand U771 (N_771,In_441,In_273);
nand U772 (N_772,In_18,In_82);
or U773 (N_773,In_3,In_225);
xnor U774 (N_774,In_86,In_311);
nand U775 (N_775,In_480,In_237);
or U776 (N_776,In_424,In_3);
or U777 (N_777,In_152,In_383);
and U778 (N_778,In_126,In_37);
nor U779 (N_779,In_414,In_136);
nand U780 (N_780,In_326,In_11);
nor U781 (N_781,In_205,In_404);
nor U782 (N_782,In_210,In_79);
and U783 (N_783,In_294,In_330);
xnor U784 (N_784,In_73,In_282);
nand U785 (N_785,In_471,In_462);
nor U786 (N_786,In_400,In_382);
nor U787 (N_787,In_494,In_380);
nand U788 (N_788,In_277,In_144);
xor U789 (N_789,In_308,In_242);
nand U790 (N_790,In_408,In_346);
xnor U791 (N_791,In_335,In_401);
nor U792 (N_792,In_104,In_168);
nor U793 (N_793,In_75,In_29);
or U794 (N_794,In_308,In_161);
or U795 (N_795,In_110,In_497);
xor U796 (N_796,In_98,In_271);
or U797 (N_797,In_370,In_442);
nand U798 (N_798,In_302,In_488);
and U799 (N_799,In_138,In_69);
xor U800 (N_800,In_185,In_439);
xor U801 (N_801,In_256,In_458);
nand U802 (N_802,In_169,In_347);
xnor U803 (N_803,In_246,In_291);
xnor U804 (N_804,In_229,In_199);
and U805 (N_805,In_108,In_462);
and U806 (N_806,In_86,In_193);
and U807 (N_807,In_379,In_489);
xor U808 (N_808,In_496,In_397);
nor U809 (N_809,In_407,In_204);
xor U810 (N_810,In_116,In_344);
and U811 (N_811,In_119,In_310);
nor U812 (N_812,In_21,In_291);
xnor U813 (N_813,In_498,In_282);
and U814 (N_814,In_392,In_433);
or U815 (N_815,In_170,In_47);
nand U816 (N_816,In_468,In_345);
xnor U817 (N_817,In_429,In_4);
nand U818 (N_818,In_14,In_31);
nand U819 (N_819,In_123,In_336);
xor U820 (N_820,In_498,In_320);
and U821 (N_821,In_131,In_497);
and U822 (N_822,In_30,In_219);
or U823 (N_823,In_30,In_255);
or U824 (N_824,In_468,In_412);
nor U825 (N_825,In_191,In_358);
or U826 (N_826,In_191,In_280);
nand U827 (N_827,In_251,In_54);
nor U828 (N_828,In_9,In_47);
nor U829 (N_829,In_101,In_338);
nor U830 (N_830,In_422,In_323);
and U831 (N_831,In_353,In_70);
xnor U832 (N_832,In_139,In_442);
xor U833 (N_833,In_403,In_326);
nor U834 (N_834,In_294,In_354);
xor U835 (N_835,In_287,In_217);
nand U836 (N_836,In_447,In_327);
nor U837 (N_837,In_42,In_182);
nor U838 (N_838,In_423,In_347);
nand U839 (N_839,In_487,In_215);
or U840 (N_840,In_251,In_451);
nor U841 (N_841,In_364,In_350);
and U842 (N_842,In_50,In_320);
nand U843 (N_843,In_219,In_43);
and U844 (N_844,In_16,In_367);
or U845 (N_845,In_499,In_488);
or U846 (N_846,In_176,In_370);
nor U847 (N_847,In_190,In_424);
nor U848 (N_848,In_102,In_139);
and U849 (N_849,In_141,In_68);
nand U850 (N_850,In_395,In_381);
nor U851 (N_851,In_46,In_74);
or U852 (N_852,In_308,In_177);
xnor U853 (N_853,In_301,In_341);
and U854 (N_854,In_181,In_264);
nor U855 (N_855,In_149,In_477);
or U856 (N_856,In_145,In_471);
and U857 (N_857,In_26,In_450);
or U858 (N_858,In_119,In_74);
and U859 (N_859,In_477,In_390);
and U860 (N_860,In_99,In_343);
xnor U861 (N_861,In_499,In_7);
xor U862 (N_862,In_475,In_5);
nand U863 (N_863,In_442,In_369);
or U864 (N_864,In_85,In_5);
and U865 (N_865,In_476,In_302);
nor U866 (N_866,In_225,In_433);
nand U867 (N_867,In_101,In_79);
nand U868 (N_868,In_20,In_381);
and U869 (N_869,In_380,In_73);
or U870 (N_870,In_165,In_305);
or U871 (N_871,In_371,In_59);
nor U872 (N_872,In_356,In_486);
xnor U873 (N_873,In_213,In_419);
nand U874 (N_874,In_12,In_267);
and U875 (N_875,In_230,In_132);
and U876 (N_876,In_280,In_113);
or U877 (N_877,In_372,In_147);
xnor U878 (N_878,In_384,In_233);
xor U879 (N_879,In_97,In_160);
and U880 (N_880,In_152,In_11);
nor U881 (N_881,In_356,In_454);
nor U882 (N_882,In_318,In_10);
and U883 (N_883,In_381,In_384);
and U884 (N_884,In_111,In_191);
and U885 (N_885,In_353,In_483);
and U886 (N_886,In_431,In_489);
and U887 (N_887,In_73,In_221);
nand U888 (N_888,In_225,In_333);
nand U889 (N_889,In_374,In_391);
xor U890 (N_890,In_146,In_429);
or U891 (N_891,In_119,In_268);
or U892 (N_892,In_327,In_211);
xnor U893 (N_893,In_3,In_212);
nand U894 (N_894,In_308,In_427);
nor U895 (N_895,In_172,In_258);
nand U896 (N_896,In_112,In_418);
nand U897 (N_897,In_79,In_290);
and U898 (N_898,In_431,In_271);
or U899 (N_899,In_465,In_94);
or U900 (N_900,In_291,In_279);
and U901 (N_901,In_450,In_238);
xnor U902 (N_902,In_346,In_331);
nor U903 (N_903,In_290,In_486);
nand U904 (N_904,In_170,In_85);
nor U905 (N_905,In_269,In_433);
xor U906 (N_906,In_177,In_424);
and U907 (N_907,In_447,In_365);
nor U908 (N_908,In_158,In_44);
nor U909 (N_909,In_466,In_333);
xor U910 (N_910,In_262,In_216);
xnor U911 (N_911,In_12,In_328);
or U912 (N_912,In_57,In_55);
nor U913 (N_913,In_419,In_126);
nand U914 (N_914,In_381,In_192);
and U915 (N_915,In_6,In_125);
nor U916 (N_916,In_430,In_174);
or U917 (N_917,In_205,In_334);
nor U918 (N_918,In_90,In_83);
and U919 (N_919,In_145,In_130);
or U920 (N_920,In_481,In_316);
and U921 (N_921,In_237,In_305);
nor U922 (N_922,In_483,In_6);
or U923 (N_923,In_251,In_5);
xor U924 (N_924,In_187,In_339);
or U925 (N_925,In_128,In_153);
xor U926 (N_926,In_158,In_312);
nor U927 (N_927,In_493,In_356);
nor U928 (N_928,In_398,In_386);
xnor U929 (N_929,In_282,In_454);
and U930 (N_930,In_328,In_120);
and U931 (N_931,In_382,In_250);
nor U932 (N_932,In_13,In_228);
nand U933 (N_933,In_415,In_192);
nor U934 (N_934,In_282,In_89);
xor U935 (N_935,In_165,In_148);
nor U936 (N_936,In_196,In_374);
xor U937 (N_937,In_219,In_152);
and U938 (N_938,In_437,In_74);
xor U939 (N_939,In_430,In_18);
or U940 (N_940,In_232,In_4);
or U941 (N_941,In_60,In_313);
nor U942 (N_942,In_492,In_355);
nor U943 (N_943,In_339,In_52);
nor U944 (N_944,In_285,In_306);
xor U945 (N_945,In_10,In_346);
nand U946 (N_946,In_276,In_338);
xor U947 (N_947,In_81,In_93);
xnor U948 (N_948,In_5,In_169);
and U949 (N_949,In_144,In_408);
or U950 (N_950,In_15,In_284);
nand U951 (N_951,In_285,In_311);
and U952 (N_952,In_31,In_322);
nor U953 (N_953,In_94,In_485);
nand U954 (N_954,In_206,In_496);
and U955 (N_955,In_386,In_408);
nor U956 (N_956,In_123,In_90);
xor U957 (N_957,In_20,In_7);
xor U958 (N_958,In_213,In_144);
or U959 (N_959,In_340,In_190);
nand U960 (N_960,In_375,In_123);
xor U961 (N_961,In_47,In_382);
nor U962 (N_962,In_432,In_66);
nor U963 (N_963,In_285,In_325);
or U964 (N_964,In_75,In_333);
nor U965 (N_965,In_330,In_335);
nand U966 (N_966,In_131,In_445);
nand U967 (N_967,In_316,In_59);
xnor U968 (N_968,In_261,In_248);
and U969 (N_969,In_12,In_248);
nor U970 (N_970,In_397,In_314);
nor U971 (N_971,In_307,In_340);
nor U972 (N_972,In_360,In_297);
nor U973 (N_973,In_330,In_298);
and U974 (N_974,In_363,In_303);
nand U975 (N_975,In_426,In_396);
nor U976 (N_976,In_405,In_408);
or U977 (N_977,In_53,In_119);
nor U978 (N_978,In_296,In_468);
and U979 (N_979,In_409,In_227);
and U980 (N_980,In_244,In_324);
xnor U981 (N_981,In_450,In_123);
nand U982 (N_982,In_194,In_451);
nor U983 (N_983,In_183,In_68);
and U984 (N_984,In_90,In_231);
or U985 (N_985,In_328,In_85);
nor U986 (N_986,In_473,In_165);
xor U987 (N_987,In_33,In_36);
nor U988 (N_988,In_102,In_223);
or U989 (N_989,In_386,In_251);
or U990 (N_990,In_251,In_498);
nor U991 (N_991,In_232,In_112);
or U992 (N_992,In_31,In_493);
or U993 (N_993,In_486,In_105);
nor U994 (N_994,In_171,In_16);
xor U995 (N_995,In_125,In_410);
nor U996 (N_996,In_28,In_316);
or U997 (N_997,In_455,In_300);
xor U998 (N_998,In_192,In_167);
xor U999 (N_999,In_7,In_66);
or U1000 (N_1000,N_532,N_166);
and U1001 (N_1001,N_117,N_867);
xor U1002 (N_1002,N_839,N_374);
xnor U1003 (N_1003,N_292,N_649);
or U1004 (N_1004,N_865,N_610);
nor U1005 (N_1005,N_35,N_660);
or U1006 (N_1006,N_54,N_555);
or U1007 (N_1007,N_545,N_114);
xnor U1008 (N_1008,N_92,N_999);
nand U1009 (N_1009,N_133,N_709);
nor U1010 (N_1010,N_426,N_457);
nand U1011 (N_1011,N_352,N_847);
and U1012 (N_1012,N_978,N_364);
or U1013 (N_1013,N_681,N_155);
or U1014 (N_1014,N_105,N_298);
and U1015 (N_1015,N_198,N_517);
and U1016 (N_1016,N_349,N_551);
xor U1017 (N_1017,N_849,N_227);
nand U1018 (N_1018,N_486,N_738);
nand U1019 (N_1019,N_110,N_537);
xor U1020 (N_1020,N_548,N_846);
nand U1021 (N_1021,N_553,N_630);
nor U1022 (N_1022,N_52,N_47);
or U1023 (N_1023,N_936,N_496);
nand U1024 (N_1024,N_890,N_515);
nand U1025 (N_1025,N_564,N_115);
and U1026 (N_1026,N_26,N_225);
or U1027 (N_1027,N_309,N_642);
and U1028 (N_1028,N_279,N_324);
xor U1029 (N_1029,N_747,N_346);
nand U1030 (N_1030,N_932,N_192);
nand U1031 (N_1031,N_565,N_882);
or U1032 (N_1032,N_245,N_488);
or U1033 (N_1033,N_519,N_755);
xnor U1034 (N_1034,N_69,N_211);
xnor U1035 (N_1035,N_434,N_123);
nor U1036 (N_1036,N_692,N_990);
and U1037 (N_1037,N_577,N_760);
nand U1038 (N_1038,N_857,N_881);
or U1039 (N_1039,N_343,N_247);
nor U1040 (N_1040,N_575,N_776);
nand U1041 (N_1041,N_726,N_810);
nor U1042 (N_1042,N_106,N_684);
or U1043 (N_1043,N_243,N_480);
nor U1044 (N_1044,N_419,N_764);
xnor U1045 (N_1045,N_39,N_199);
nor U1046 (N_1046,N_997,N_23);
nor U1047 (N_1047,N_955,N_395);
or U1048 (N_1048,N_204,N_58);
nand U1049 (N_1049,N_369,N_396);
and U1050 (N_1050,N_896,N_503);
nor U1051 (N_1051,N_912,N_840);
xor U1052 (N_1052,N_914,N_948);
nor U1053 (N_1053,N_898,N_843);
nor U1054 (N_1054,N_841,N_613);
xnor U1055 (N_1055,N_66,N_705);
nand U1056 (N_1056,N_32,N_916);
nand U1057 (N_1057,N_530,N_987);
and U1058 (N_1058,N_191,N_94);
nor U1059 (N_1059,N_226,N_716);
or U1060 (N_1060,N_802,N_653);
or U1061 (N_1061,N_72,N_677);
nand U1062 (N_1062,N_327,N_145);
nor U1063 (N_1063,N_976,N_41);
and U1064 (N_1064,N_656,N_201);
xnor U1065 (N_1065,N_73,N_304);
xor U1066 (N_1066,N_528,N_661);
and U1067 (N_1067,N_177,N_989);
and U1068 (N_1068,N_576,N_290);
nor U1069 (N_1069,N_627,N_38);
xnor U1070 (N_1070,N_391,N_638);
nor U1071 (N_1071,N_70,N_864);
xor U1072 (N_1072,N_959,N_996);
and U1073 (N_1073,N_13,N_446);
and U1074 (N_1074,N_650,N_734);
xnor U1075 (N_1075,N_658,N_621);
or U1076 (N_1076,N_383,N_8);
and U1077 (N_1077,N_851,N_569);
and U1078 (N_1078,N_558,N_877);
or U1079 (N_1079,N_467,N_652);
nand U1080 (N_1080,N_824,N_90);
nand U1081 (N_1081,N_906,N_602);
xor U1082 (N_1082,N_688,N_823);
or U1083 (N_1083,N_521,N_982);
nor U1084 (N_1084,N_580,N_965);
or U1085 (N_1085,N_63,N_272);
nand U1086 (N_1086,N_100,N_56);
xnor U1087 (N_1087,N_617,N_927);
xor U1088 (N_1088,N_572,N_379);
nand U1089 (N_1089,N_428,N_282);
nor U1090 (N_1090,N_414,N_445);
and U1091 (N_1091,N_132,N_510);
or U1092 (N_1092,N_808,N_502);
and U1093 (N_1093,N_326,N_274);
or U1094 (N_1094,N_745,N_728);
nand U1095 (N_1095,N_703,N_669);
and U1096 (N_1096,N_368,N_281);
or U1097 (N_1097,N_601,N_471);
and U1098 (N_1098,N_163,N_271);
nand U1099 (N_1099,N_303,N_422);
nor U1100 (N_1100,N_819,N_888);
nor U1101 (N_1101,N_934,N_77);
xnor U1102 (N_1102,N_233,N_71);
and U1103 (N_1103,N_562,N_981);
nor U1104 (N_1104,N_401,N_345);
or U1105 (N_1105,N_970,N_767);
or U1106 (N_1106,N_98,N_875);
xor U1107 (N_1107,N_822,N_796);
or U1108 (N_1108,N_746,N_501);
and U1109 (N_1109,N_311,N_659);
nand U1110 (N_1110,N_871,N_852);
nor U1111 (N_1111,N_625,N_672);
and U1112 (N_1112,N_818,N_620);
and U1113 (N_1113,N_607,N_180);
nand U1114 (N_1114,N_64,N_963);
nor U1115 (N_1115,N_557,N_430);
or U1116 (N_1116,N_128,N_778);
nand U1117 (N_1117,N_112,N_167);
and U1118 (N_1118,N_244,N_826);
or U1119 (N_1119,N_219,N_79);
and U1120 (N_1120,N_749,N_696);
xnor U1121 (N_1121,N_868,N_20);
and U1122 (N_1122,N_968,N_68);
and U1123 (N_1123,N_24,N_312);
or U1124 (N_1124,N_992,N_10);
or U1125 (N_1125,N_803,N_933);
nand U1126 (N_1126,N_240,N_332);
nand U1127 (N_1127,N_831,N_78);
or U1128 (N_1128,N_65,N_122);
and U1129 (N_1129,N_435,N_815);
or U1130 (N_1130,N_774,N_61);
xor U1131 (N_1131,N_724,N_231);
nand U1132 (N_1132,N_769,N_581);
and U1133 (N_1133,N_685,N_319);
and U1134 (N_1134,N_483,N_805);
nor U1135 (N_1135,N_433,N_397);
nor U1136 (N_1136,N_950,N_450);
xnor U1137 (N_1137,N_585,N_60);
or U1138 (N_1138,N_59,N_615);
or U1139 (N_1139,N_269,N_179);
or U1140 (N_1140,N_478,N_729);
nor U1141 (N_1141,N_855,N_498);
nand U1142 (N_1142,N_294,N_30);
nand U1143 (N_1143,N_152,N_811);
xnor U1144 (N_1144,N_783,N_333);
or U1145 (N_1145,N_468,N_238);
or U1146 (N_1146,N_829,N_230);
or U1147 (N_1147,N_215,N_624);
xor U1148 (N_1148,N_402,N_842);
nand U1149 (N_1149,N_780,N_858);
nor U1150 (N_1150,N_5,N_883);
and U1151 (N_1151,N_276,N_908);
and U1152 (N_1152,N_812,N_917);
and U1153 (N_1153,N_40,N_209);
xnor U1154 (N_1154,N_463,N_506);
or U1155 (N_1155,N_554,N_474);
or U1156 (N_1156,N_361,N_736);
or U1157 (N_1157,N_331,N_687);
or U1158 (N_1158,N_801,N_925);
nor U1159 (N_1159,N_157,N_140);
and U1160 (N_1160,N_214,N_598);
xor U1161 (N_1161,N_340,N_360);
and U1162 (N_1162,N_451,N_619);
or U1163 (N_1163,N_33,N_208);
nand U1164 (N_1164,N_777,N_880);
nor U1165 (N_1165,N_249,N_389);
nand U1166 (N_1166,N_759,N_991);
nand U1167 (N_1167,N_228,N_588);
xnor U1168 (N_1168,N_518,N_377);
xor U1169 (N_1169,N_953,N_178);
xnor U1170 (N_1170,N_590,N_974);
and U1171 (N_1171,N_522,N_482);
nor U1172 (N_1172,N_499,N_629);
and U1173 (N_1173,N_646,N_194);
nor U1174 (N_1174,N_935,N_512);
nand U1175 (N_1175,N_641,N_334);
xor U1176 (N_1176,N_489,N_221);
nand U1177 (N_1177,N_437,N_96);
or U1178 (N_1178,N_816,N_946);
or U1179 (N_1179,N_97,N_570);
nand U1180 (N_1180,N_504,N_727);
nor U1181 (N_1181,N_126,N_16);
nand U1182 (N_1182,N_797,N_51);
nor U1183 (N_1183,N_689,N_479);
or U1184 (N_1184,N_994,N_534);
nor U1185 (N_1185,N_121,N_573);
nor U1186 (N_1186,N_862,N_931);
xnor U1187 (N_1187,N_578,N_310);
nor U1188 (N_1188,N_961,N_359);
or U1189 (N_1189,N_807,N_357);
and U1190 (N_1190,N_144,N_36);
or U1191 (N_1191,N_623,N_164);
nand U1192 (N_1192,N_901,N_938);
and U1193 (N_1193,N_964,N_930);
or U1194 (N_1194,N_984,N_275);
or U1195 (N_1195,N_835,N_266);
nor U1196 (N_1196,N_207,N_306);
nor U1197 (N_1197,N_365,N_142);
xor U1198 (N_1198,N_469,N_22);
nor U1199 (N_1199,N_323,N_866);
xor U1200 (N_1200,N_655,N_265);
or U1201 (N_1201,N_514,N_213);
nand U1202 (N_1202,N_109,N_466);
or U1203 (N_1203,N_337,N_693);
and U1204 (N_1204,N_717,N_859);
and U1205 (N_1205,N_43,N_427);
nand U1206 (N_1206,N_257,N_611);
nor U1207 (N_1207,N_785,N_605);
or U1208 (N_1208,N_270,N_295);
or U1209 (N_1209,N_246,N_465);
xor U1210 (N_1210,N_205,N_367);
nand U1211 (N_1211,N_113,N_600);
xor U1212 (N_1212,N_436,N_967);
or U1213 (N_1213,N_62,N_863);
nand U1214 (N_1214,N_673,N_386);
nor U1215 (N_1215,N_339,N_186);
nand U1216 (N_1216,N_739,N_477);
and U1217 (N_1217,N_766,N_520);
nand U1218 (N_1218,N_637,N_644);
nor U1219 (N_1219,N_668,N_907);
nor U1220 (N_1220,N_293,N_256);
nor U1221 (N_1221,N_143,N_657);
xnor U1222 (N_1222,N_160,N_595);
and U1223 (N_1223,N_348,N_790);
xnor U1224 (N_1224,N_666,N_779);
nor U1225 (N_1225,N_516,N_542);
nand U1226 (N_1226,N_103,N_330);
or U1227 (N_1227,N_886,N_95);
nor U1228 (N_1228,N_174,N_161);
nor U1229 (N_1229,N_549,N_329);
or U1230 (N_1230,N_561,N_772);
xor U1231 (N_1231,N_552,N_318);
nand U1232 (N_1232,N_720,N_476);
and U1233 (N_1233,N_472,N_628);
nand U1234 (N_1234,N_686,N_314);
or U1235 (N_1235,N_118,N_381);
xor U1236 (N_1236,N_57,N_743);
xor U1237 (N_1237,N_193,N_492);
nand U1238 (N_1238,N_945,N_757);
or U1239 (N_1239,N_44,N_850);
xnor U1240 (N_1240,N_500,N_497);
xor U1241 (N_1241,N_37,N_836);
nor U1242 (N_1242,N_455,N_511);
nand U1243 (N_1243,N_399,N_612);
or U1244 (N_1244,N_975,N_574);
or U1245 (N_1245,N_320,N_284);
nor U1246 (N_1246,N_242,N_74);
nor U1247 (N_1247,N_694,N_176);
xor U1248 (N_1248,N_550,N_280);
or U1249 (N_1249,N_583,N_639);
or U1250 (N_1250,N_988,N_856);
nand U1251 (N_1251,N_929,N_892);
nand U1252 (N_1252,N_973,N_131);
and U1253 (N_1253,N_338,N_756);
xnor U1254 (N_1254,N_305,N_385);
nor U1255 (N_1255,N_321,N_387);
or U1256 (N_1256,N_150,N_316);
nor U1257 (N_1257,N_217,N_845);
xor U1258 (N_1258,N_972,N_640);
xor U1259 (N_1259,N_232,N_29);
or U1260 (N_1260,N_116,N_363);
nand U1261 (N_1261,N_636,N_546);
nand U1262 (N_1262,N_34,N_526);
or U1263 (N_1263,N_667,N_18);
or U1264 (N_1264,N_366,N_529);
xnor U1265 (N_1265,N_248,N_586);
xnor U1266 (N_1266,N_335,N_301);
and U1267 (N_1267,N_782,N_513);
nor U1268 (N_1268,N_151,N_926);
nand U1269 (N_1269,N_631,N_136);
nor U1270 (N_1270,N_42,N_962);
nor U1271 (N_1271,N_531,N_909);
and U1272 (N_1272,N_108,N_358);
or U1273 (N_1273,N_210,N_336);
nand U1274 (N_1274,N_791,N_887);
xor U1275 (N_1275,N_168,N_566);
nand U1276 (N_1276,N_559,N_375);
xor U1277 (N_1277,N_853,N_287);
xnor U1278 (N_1278,N_919,N_543);
and U1279 (N_1279,N_317,N_922);
nor U1280 (N_1280,N_2,N_99);
or U1281 (N_1281,N_879,N_770);
and U1282 (N_1282,N_763,N_353);
nand U1283 (N_1283,N_708,N_394);
nand U1284 (N_1284,N_920,N_942);
nor U1285 (N_1285,N_789,N_203);
nand U1286 (N_1286,N_404,N_407);
nand U1287 (N_1287,N_643,N_216);
nor U1288 (N_1288,N_1,N_45);
or U1289 (N_1289,N_674,N_408);
nand U1290 (N_1290,N_351,N_443);
nor U1291 (N_1291,N_158,N_682);
and U1292 (N_1292,N_960,N_251);
nor U1293 (N_1293,N_834,N_737);
nand U1294 (N_1294,N_91,N_568);
nor U1295 (N_1295,N_169,N_165);
nor U1296 (N_1296,N_966,N_718);
xor U1297 (N_1297,N_4,N_184);
or U1298 (N_1298,N_795,N_277);
xor U1299 (N_1299,N_495,N_609);
and U1300 (N_1300,N_732,N_135);
nand U1301 (N_1301,N_21,N_170);
nand U1302 (N_1302,N_715,N_924);
and U1303 (N_1303,N_254,N_187);
xor U1304 (N_1304,N_538,N_129);
xnor U1305 (N_1305,N_236,N_260);
nand U1306 (N_1306,N_183,N_125);
xnor U1307 (N_1307,N_384,N_263);
xnor U1308 (N_1308,N_372,N_665);
and U1309 (N_1309,N_189,N_382);
nand U1310 (N_1310,N_172,N_235);
nand U1311 (N_1311,N_758,N_241);
or U1312 (N_1312,N_910,N_154);
or U1313 (N_1313,N_252,N_804);
and U1314 (N_1314,N_897,N_809);
or U1315 (N_1315,N_596,N_119);
xnor U1316 (N_1316,N_944,N_438);
nand U1317 (N_1317,N_484,N_239);
nand U1318 (N_1318,N_765,N_149);
nand U1319 (N_1319,N_535,N_283);
or U1320 (N_1320,N_902,N_400);
nor U1321 (N_1321,N_458,N_706);
xor U1322 (N_1322,N_828,N_89);
or U1323 (N_1323,N_711,N_918);
xor U1324 (N_1324,N_899,N_632);
and U1325 (N_1325,N_147,N_723);
and U1326 (N_1326,N_606,N_420);
nor U1327 (N_1327,N_761,N_49);
nand U1328 (N_1328,N_262,N_313);
and U1329 (N_1329,N_876,N_127);
or U1330 (N_1330,N_784,N_196);
and U1331 (N_1331,N_411,N_76);
nand U1332 (N_1332,N_947,N_7);
xor U1333 (N_1333,N_181,N_456);
nor U1334 (N_1334,N_481,N_376);
or U1335 (N_1335,N_579,N_825);
xnor U1336 (N_1336,N_680,N_224);
or U1337 (N_1337,N_28,N_425);
and U1338 (N_1338,N_921,N_884);
nor U1339 (N_1339,N_714,N_173);
nand U1340 (N_1340,N_775,N_951);
nand U1341 (N_1341,N_218,N_793);
and U1342 (N_1342,N_81,N_995);
xnor U1343 (N_1343,N_285,N_648);
xor U1344 (N_1344,N_905,N_593);
or U1345 (N_1345,N_261,N_302);
nor U1346 (N_1346,N_403,N_900);
nand U1347 (N_1347,N_740,N_751);
and U1348 (N_1348,N_915,N_447);
nor U1349 (N_1349,N_423,N_893);
nor U1350 (N_1350,N_487,N_683);
nor U1351 (N_1351,N_453,N_985);
nor U1352 (N_1352,N_297,N_874);
nor U1353 (N_1353,N_195,N_440);
and U1354 (N_1354,N_539,N_398);
xor U1355 (N_1355,N_124,N_373);
or U1356 (N_1356,N_787,N_750);
nor U1357 (N_1357,N_589,N_413);
xnor U1358 (N_1358,N_444,N_928);
or U1359 (N_1359,N_730,N_977);
xnor U1360 (N_1360,N_162,N_786);
nand U1361 (N_1361,N_702,N_75);
or U1362 (N_1362,N_664,N_25);
xnor U1363 (N_1363,N_773,N_536);
or U1364 (N_1364,N_837,N_663);
nand U1365 (N_1365,N_541,N_53);
or U1366 (N_1366,N_820,N_547);
and U1367 (N_1367,N_821,N_197);
nor U1368 (N_1368,N_212,N_85);
nor U1369 (N_1369,N_355,N_200);
nor U1370 (N_1370,N_182,N_651);
xnor U1371 (N_1371,N_523,N_344);
nor U1372 (N_1372,N_993,N_412);
nand U1373 (N_1373,N_223,N_634);
or U1374 (N_1374,N_84,N_31);
or U1375 (N_1375,N_255,N_137);
xor U1376 (N_1376,N_153,N_234);
nor U1377 (N_1377,N_647,N_699);
and U1378 (N_1378,N_584,N_80);
and U1379 (N_1379,N_540,N_998);
nor U1380 (N_1380,N_788,N_409);
nand U1381 (N_1381,N_690,N_87);
nor U1382 (N_1382,N_278,N_139);
xnor U1383 (N_1383,N_417,N_104);
or U1384 (N_1384,N_697,N_582);
and U1385 (N_1385,N_464,N_347);
and U1386 (N_1386,N_618,N_286);
nand U1387 (N_1387,N_870,N_792);
and U1388 (N_1388,N_253,N_671);
nor U1389 (N_1389,N_833,N_291);
xor U1390 (N_1390,N_55,N_645);
and U1391 (N_1391,N_806,N_459);
or U1392 (N_1392,N_9,N_670);
nor U1393 (N_1393,N_980,N_952);
nand U1394 (N_1394,N_662,N_762);
xor U1395 (N_1395,N_567,N_415);
or U1396 (N_1396,N_533,N_442);
nand U1397 (N_1397,N_861,N_679);
xor U1398 (N_1398,N_120,N_721);
nand U1399 (N_1399,N_698,N_141);
and U1400 (N_1400,N_872,N_904);
nand U1401 (N_1401,N_603,N_350);
and U1402 (N_1402,N_704,N_431);
nand U1403 (N_1403,N_695,N_494);
nand U1404 (N_1404,N_490,N_911);
xnor U1405 (N_1405,N_111,N_700);
xnor U1406 (N_1406,N_88,N_691);
or U1407 (N_1407,N_941,N_50);
nor U1408 (N_1408,N_885,N_838);
nor U1409 (N_1409,N_869,N_707);
or U1410 (N_1410,N_712,N_940);
or U1411 (N_1411,N_958,N_626);
or U1412 (N_1412,N_429,N_903);
xor U1413 (N_1413,N_814,N_470);
nor U1414 (N_1414,N_6,N_722);
or U1415 (N_1415,N_393,N_300);
or U1416 (N_1416,N_509,N_571);
nand U1417 (N_1417,N_424,N_986);
or U1418 (N_1418,N_406,N_273);
or U1419 (N_1419,N_923,N_594);
and U1420 (N_1420,N_800,N_388);
xor U1421 (N_1421,N_954,N_956);
nand U1422 (N_1422,N_969,N_701);
nand U1423 (N_1423,N_156,N_449);
and U1424 (N_1424,N_622,N_979);
and U1425 (N_1425,N_591,N_308);
or U1426 (N_1426,N_202,N_735);
nand U1427 (N_1427,N_83,N_138);
and U1428 (N_1428,N_485,N_493);
xnor U1429 (N_1429,N_86,N_432);
nor U1430 (N_1430,N_159,N_93);
xnor U1431 (N_1431,N_741,N_148);
nand U1432 (N_1432,N_744,N_604);
or U1433 (N_1433,N_416,N_676);
and U1434 (N_1434,N_742,N_894);
and U1435 (N_1435,N_370,N_421);
nand U1436 (N_1436,N_354,N_616);
or U1437 (N_1437,N_889,N_848);
nand U1438 (N_1438,N_380,N_556);
nor U1439 (N_1439,N_250,N_710);
or U1440 (N_1440,N_527,N_713);
nor U1441 (N_1441,N_798,N_983);
nor U1442 (N_1442,N_19,N_794);
and U1443 (N_1443,N_371,N_27);
xnor U1444 (N_1444,N_102,N_971);
nor U1445 (N_1445,N_461,N_299);
nand U1446 (N_1446,N_362,N_264);
xor U1447 (N_1447,N_752,N_525);
or U1448 (N_1448,N_258,N_462);
xnor U1449 (N_1449,N_448,N_654);
or U1450 (N_1450,N_608,N_441);
xor U1451 (N_1451,N_597,N_943);
nand U1452 (N_1452,N_15,N_17);
nor U1453 (N_1453,N_222,N_799);
nor U1454 (N_1454,N_322,N_67);
xor U1455 (N_1455,N_827,N_505);
xnor U1456 (N_1456,N_508,N_259);
or U1457 (N_1457,N_206,N_830);
nand U1458 (N_1458,N_325,N_46);
or U1459 (N_1459,N_635,N_587);
xnor U1460 (N_1460,N_733,N_939);
and U1461 (N_1461,N_719,N_891);
or U1462 (N_1462,N_267,N_190);
nor U1463 (N_1463,N_289,N_753);
and U1464 (N_1464,N_560,N_817);
and U1465 (N_1465,N_48,N_229);
xnor U1466 (N_1466,N_12,N_268);
xor U1467 (N_1467,N_768,N_452);
nor U1468 (N_1468,N_475,N_11);
xnor U1469 (N_1469,N_957,N_771);
nor U1470 (N_1470,N_725,N_592);
and U1471 (N_1471,N_220,N_748);
nand U1472 (N_1472,N_832,N_844);
xnor U1473 (N_1473,N_288,N_524);
nor U1474 (N_1474,N_675,N_873);
or U1475 (N_1475,N_473,N_563);
or U1476 (N_1476,N_754,N_405);
xor U1477 (N_1477,N_307,N_3);
or U1478 (N_1478,N_860,N_439);
nor U1479 (N_1479,N_378,N_813);
xor U1480 (N_1480,N_175,N_296);
nand U1481 (N_1481,N_544,N_491);
nor U1482 (N_1482,N_101,N_878);
or U1483 (N_1483,N_82,N_731);
nand U1484 (N_1484,N_678,N_14);
and U1485 (N_1485,N_460,N_781);
and U1486 (N_1486,N_315,N_237);
or U1487 (N_1487,N_895,N_418);
and U1488 (N_1488,N_356,N_146);
nand U1489 (N_1489,N_0,N_341);
nand U1490 (N_1490,N_410,N_188);
or U1491 (N_1491,N_599,N_171);
nand U1492 (N_1492,N_342,N_854);
or U1493 (N_1493,N_633,N_454);
nor U1494 (N_1494,N_614,N_390);
or U1495 (N_1495,N_949,N_107);
nor U1496 (N_1496,N_328,N_130);
nor U1497 (N_1497,N_913,N_134);
nor U1498 (N_1498,N_507,N_185);
xor U1499 (N_1499,N_937,N_392);
nor U1500 (N_1500,N_9,N_743);
or U1501 (N_1501,N_844,N_872);
or U1502 (N_1502,N_834,N_871);
xnor U1503 (N_1503,N_447,N_118);
nand U1504 (N_1504,N_576,N_822);
xnor U1505 (N_1505,N_392,N_146);
or U1506 (N_1506,N_497,N_224);
nor U1507 (N_1507,N_428,N_564);
nor U1508 (N_1508,N_305,N_687);
nor U1509 (N_1509,N_40,N_916);
or U1510 (N_1510,N_873,N_724);
and U1511 (N_1511,N_463,N_141);
nor U1512 (N_1512,N_672,N_542);
nor U1513 (N_1513,N_253,N_132);
xor U1514 (N_1514,N_170,N_715);
and U1515 (N_1515,N_533,N_853);
or U1516 (N_1516,N_511,N_92);
nor U1517 (N_1517,N_249,N_917);
nor U1518 (N_1518,N_792,N_229);
nand U1519 (N_1519,N_463,N_833);
or U1520 (N_1520,N_902,N_355);
xor U1521 (N_1521,N_24,N_539);
nand U1522 (N_1522,N_100,N_646);
or U1523 (N_1523,N_796,N_700);
xnor U1524 (N_1524,N_627,N_540);
nor U1525 (N_1525,N_910,N_713);
or U1526 (N_1526,N_810,N_106);
or U1527 (N_1527,N_750,N_517);
nand U1528 (N_1528,N_128,N_213);
nand U1529 (N_1529,N_877,N_120);
or U1530 (N_1530,N_514,N_281);
xor U1531 (N_1531,N_258,N_528);
xor U1532 (N_1532,N_262,N_500);
or U1533 (N_1533,N_62,N_488);
and U1534 (N_1534,N_853,N_345);
xnor U1535 (N_1535,N_290,N_297);
or U1536 (N_1536,N_889,N_716);
or U1537 (N_1537,N_133,N_303);
nand U1538 (N_1538,N_327,N_59);
or U1539 (N_1539,N_590,N_379);
nand U1540 (N_1540,N_570,N_961);
nand U1541 (N_1541,N_210,N_884);
xor U1542 (N_1542,N_266,N_203);
xnor U1543 (N_1543,N_408,N_99);
nand U1544 (N_1544,N_80,N_137);
xnor U1545 (N_1545,N_424,N_391);
nor U1546 (N_1546,N_291,N_716);
xor U1547 (N_1547,N_730,N_426);
nand U1548 (N_1548,N_107,N_938);
or U1549 (N_1549,N_870,N_724);
xor U1550 (N_1550,N_313,N_461);
nand U1551 (N_1551,N_220,N_296);
xnor U1552 (N_1552,N_793,N_558);
nand U1553 (N_1553,N_204,N_700);
or U1554 (N_1554,N_318,N_75);
and U1555 (N_1555,N_360,N_198);
xnor U1556 (N_1556,N_851,N_464);
nand U1557 (N_1557,N_703,N_371);
xnor U1558 (N_1558,N_280,N_139);
nand U1559 (N_1559,N_297,N_113);
xor U1560 (N_1560,N_255,N_319);
nand U1561 (N_1561,N_49,N_492);
xor U1562 (N_1562,N_227,N_889);
nand U1563 (N_1563,N_86,N_470);
and U1564 (N_1564,N_296,N_132);
or U1565 (N_1565,N_759,N_828);
xnor U1566 (N_1566,N_130,N_49);
nor U1567 (N_1567,N_772,N_608);
nor U1568 (N_1568,N_201,N_912);
nand U1569 (N_1569,N_669,N_509);
nor U1570 (N_1570,N_232,N_261);
nand U1571 (N_1571,N_125,N_433);
nand U1572 (N_1572,N_926,N_953);
and U1573 (N_1573,N_563,N_859);
and U1574 (N_1574,N_383,N_748);
and U1575 (N_1575,N_545,N_169);
nand U1576 (N_1576,N_122,N_157);
and U1577 (N_1577,N_787,N_291);
nor U1578 (N_1578,N_720,N_161);
xor U1579 (N_1579,N_383,N_71);
nand U1580 (N_1580,N_606,N_823);
nand U1581 (N_1581,N_526,N_356);
nor U1582 (N_1582,N_954,N_838);
or U1583 (N_1583,N_812,N_154);
nor U1584 (N_1584,N_643,N_374);
and U1585 (N_1585,N_693,N_968);
xnor U1586 (N_1586,N_814,N_93);
nand U1587 (N_1587,N_146,N_669);
nand U1588 (N_1588,N_171,N_761);
or U1589 (N_1589,N_278,N_339);
nand U1590 (N_1590,N_136,N_687);
nor U1591 (N_1591,N_445,N_732);
and U1592 (N_1592,N_876,N_100);
xnor U1593 (N_1593,N_6,N_10);
or U1594 (N_1594,N_708,N_495);
xor U1595 (N_1595,N_701,N_347);
nand U1596 (N_1596,N_589,N_19);
xor U1597 (N_1597,N_905,N_928);
nand U1598 (N_1598,N_703,N_577);
and U1599 (N_1599,N_983,N_957);
and U1600 (N_1600,N_542,N_52);
and U1601 (N_1601,N_726,N_239);
or U1602 (N_1602,N_668,N_719);
nor U1603 (N_1603,N_55,N_843);
nor U1604 (N_1604,N_397,N_10);
nor U1605 (N_1605,N_282,N_452);
xor U1606 (N_1606,N_219,N_454);
nor U1607 (N_1607,N_999,N_285);
nor U1608 (N_1608,N_750,N_945);
nand U1609 (N_1609,N_255,N_553);
nand U1610 (N_1610,N_161,N_757);
nand U1611 (N_1611,N_561,N_524);
nor U1612 (N_1612,N_444,N_165);
or U1613 (N_1613,N_966,N_950);
nand U1614 (N_1614,N_948,N_144);
nand U1615 (N_1615,N_836,N_726);
nand U1616 (N_1616,N_499,N_641);
and U1617 (N_1617,N_859,N_472);
nor U1618 (N_1618,N_45,N_384);
and U1619 (N_1619,N_85,N_560);
and U1620 (N_1620,N_330,N_387);
nand U1621 (N_1621,N_919,N_776);
nor U1622 (N_1622,N_651,N_974);
nand U1623 (N_1623,N_95,N_122);
and U1624 (N_1624,N_219,N_743);
nor U1625 (N_1625,N_153,N_353);
and U1626 (N_1626,N_467,N_178);
and U1627 (N_1627,N_839,N_284);
and U1628 (N_1628,N_253,N_989);
or U1629 (N_1629,N_97,N_553);
nor U1630 (N_1630,N_778,N_95);
nand U1631 (N_1631,N_160,N_650);
nor U1632 (N_1632,N_369,N_657);
and U1633 (N_1633,N_148,N_590);
nand U1634 (N_1634,N_843,N_456);
and U1635 (N_1635,N_599,N_535);
nor U1636 (N_1636,N_137,N_482);
or U1637 (N_1637,N_625,N_107);
or U1638 (N_1638,N_393,N_941);
xor U1639 (N_1639,N_636,N_898);
nor U1640 (N_1640,N_920,N_518);
or U1641 (N_1641,N_289,N_109);
nor U1642 (N_1642,N_222,N_520);
xnor U1643 (N_1643,N_685,N_115);
and U1644 (N_1644,N_259,N_721);
and U1645 (N_1645,N_319,N_160);
and U1646 (N_1646,N_989,N_533);
xor U1647 (N_1647,N_221,N_189);
nand U1648 (N_1648,N_103,N_436);
nor U1649 (N_1649,N_964,N_481);
xor U1650 (N_1650,N_446,N_755);
or U1651 (N_1651,N_720,N_305);
or U1652 (N_1652,N_810,N_50);
xnor U1653 (N_1653,N_103,N_422);
xnor U1654 (N_1654,N_440,N_814);
nand U1655 (N_1655,N_445,N_114);
xor U1656 (N_1656,N_701,N_287);
nor U1657 (N_1657,N_579,N_348);
xor U1658 (N_1658,N_687,N_329);
nor U1659 (N_1659,N_548,N_406);
and U1660 (N_1660,N_539,N_113);
nand U1661 (N_1661,N_377,N_105);
nand U1662 (N_1662,N_199,N_105);
nand U1663 (N_1663,N_29,N_706);
or U1664 (N_1664,N_613,N_75);
nand U1665 (N_1665,N_851,N_740);
nor U1666 (N_1666,N_474,N_415);
nor U1667 (N_1667,N_562,N_42);
nor U1668 (N_1668,N_828,N_782);
and U1669 (N_1669,N_486,N_465);
or U1670 (N_1670,N_535,N_152);
and U1671 (N_1671,N_113,N_39);
or U1672 (N_1672,N_556,N_420);
nand U1673 (N_1673,N_861,N_959);
or U1674 (N_1674,N_613,N_451);
xor U1675 (N_1675,N_737,N_806);
nor U1676 (N_1676,N_461,N_86);
nor U1677 (N_1677,N_329,N_700);
and U1678 (N_1678,N_200,N_848);
or U1679 (N_1679,N_435,N_47);
nor U1680 (N_1680,N_136,N_37);
and U1681 (N_1681,N_808,N_642);
nand U1682 (N_1682,N_381,N_368);
nor U1683 (N_1683,N_786,N_466);
and U1684 (N_1684,N_330,N_190);
nor U1685 (N_1685,N_461,N_787);
nor U1686 (N_1686,N_132,N_881);
nand U1687 (N_1687,N_176,N_960);
or U1688 (N_1688,N_406,N_322);
nand U1689 (N_1689,N_829,N_15);
and U1690 (N_1690,N_820,N_205);
nand U1691 (N_1691,N_471,N_685);
or U1692 (N_1692,N_414,N_858);
xor U1693 (N_1693,N_821,N_142);
and U1694 (N_1694,N_138,N_0);
and U1695 (N_1695,N_859,N_707);
or U1696 (N_1696,N_657,N_821);
nor U1697 (N_1697,N_371,N_46);
nor U1698 (N_1698,N_993,N_782);
and U1699 (N_1699,N_708,N_414);
nor U1700 (N_1700,N_828,N_56);
nand U1701 (N_1701,N_106,N_792);
and U1702 (N_1702,N_381,N_575);
xor U1703 (N_1703,N_730,N_532);
nor U1704 (N_1704,N_250,N_740);
nand U1705 (N_1705,N_426,N_827);
nor U1706 (N_1706,N_118,N_545);
and U1707 (N_1707,N_603,N_731);
nor U1708 (N_1708,N_290,N_727);
nor U1709 (N_1709,N_274,N_227);
or U1710 (N_1710,N_96,N_861);
xnor U1711 (N_1711,N_388,N_530);
nand U1712 (N_1712,N_195,N_108);
or U1713 (N_1713,N_238,N_514);
nand U1714 (N_1714,N_477,N_305);
xnor U1715 (N_1715,N_485,N_161);
nand U1716 (N_1716,N_374,N_60);
or U1717 (N_1717,N_173,N_735);
and U1718 (N_1718,N_921,N_543);
or U1719 (N_1719,N_4,N_809);
nor U1720 (N_1720,N_163,N_99);
nor U1721 (N_1721,N_893,N_86);
xor U1722 (N_1722,N_757,N_437);
nand U1723 (N_1723,N_634,N_215);
nand U1724 (N_1724,N_329,N_426);
xor U1725 (N_1725,N_494,N_727);
or U1726 (N_1726,N_349,N_337);
nand U1727 (N_1727,N_471,N_721);
nor U1728 (N_1728,N_406,N_72);
xor U1729 (N_1729,N_221,N_402);
nor U1730 (N_1730,N_164,N_746);
nor U1731 (N_1731,N_826,N_780);
xor U1732 (N_1732,N_989,N_609);
and U1733 (N_1733,N_824,N_292);
or U1734 (N_1734,N_265,N_918);
xor U1735 (N_1735,N_894,N_42);
nor U1736 (N_1736,N_352,N_593);
nand U1737 (N_1737,N_194,N_784);
nor U1738 (N_1738,N_52,N_159);
nand U1739 (N_1739,N_907,N_305);
and U1740 (N_1740,N_839,N_584);
nand U1741 (N_1741,N_102,N_64);
nor U1742 (N_1742,N_904,N_258);
nor U1743 (N_1743,N_298,N_991);
nor U1744 (N_1744,N_33,N_782);
nor U1745 (N_1745,N_600,N_584);
nand U1746 (N_1746,N_392,N_498);
or U1747 (N_1747,N_629,N_615);
or U1748 (N_1748,N_612,N_484);
and U1749 (N_1749,N_948,N_990);
nor U1750 (N_1750,N_423,N_688);
or U1751 (N_1751,N_126,N_700);
or U1752 (N_1752,N_703,N_1);
and U1753 (N_1753,N_251,N_689);
nor U1754 (N_1754,N_660,N_860);
xnor U1755 (N_1755,N_96,N_204);
xor U1756 (N_1756,N_541,N_63);
or U1757 (N_1757,N_793,N_609);
nor U1758 (N_1758,N_444,N_542);
nand U1759 (N_1759,N_533,N_429);
or U1760 (N_1760,N_862,N_881);
or U1761 (N_1761,N_766,N_183);
xnor U1762 (N_1762,N_770,N_24);
xnor U1763 (N_1763,N_59,N_628);
and U1764 (N_1764,N_952,N_405);
xnor U1765 (N_1765,N_108,N_963);
or U1766 (N_1766,N_173,N_655);
and U1767 (N_1767,N_698,N_299);
xnor U1768 (N_1768,N_863,N_280);
nor U1769 (N_1769,N_727,N_811);
or U1770 (N_1770,N_263,N_961);
nand U1771 (N_1771,N_204,N_875);
and U1772 (N_1772,N_378,N_128);
and U1773 (N_1773,N_297,N_216);
nor U1774 (N_1774,N_703,N_885);
xor U1775 (N_1775,N_666,N_682);
nand U1776 (N_1776,N_31,N_686);
xnor U1777 (N_1777,N_662,N_673);
xor U1778 (N_1778,N_517,N_518);
xor U1779 (N_1779,N_124,N_491);
nor U1780 (N_1780,N_73,N_551);
or U1781 (N_1781,N_750,N_538);
or U1782 (N_1782,N_355,N_374);
nor U1783 (N_1783,N_258,N_584);
and U1784 (N_1784,N_462,N_477);
and U1785 (N_1785,N_232,N_995);
nor U1786 (N_1786,N_601,N_107);
nor U1787 (N_1787,N_842,N_339);
nor U1788 (N_1788,N_291,N_658);
and U1789 (N_1789,N_446,N_568);
nand U1790 (N_1790,N_130,N_200);
xor U1791 (N_1791,N_958,N_365);
and U1792 (N_1792,N_33,N_954);
nand U1793 (N_1793,N_392,N_455);
nand U1794 (N_1794,N_824,N_457);
or U1795 (N_1795,N_445,N_716);
nor U1796 (N_1796,N_329,N_860);
xnor U1797 (N_1797,N_958,N_369);
nor U1798 (N_1798,N_682,N_108);
nor U1799 (N_1799,N_375,N_474);
nor U1800 (N_1800,N_859,N_10);
or U1801 (N_1801,N_735,N_71);
xor U1802 (N_1802,N_358,N_730);
and U1803 (N_1803,N_266,N_865);
xnor U1804 (N_1804,N_925,N_743);
nor U1805 (N_1805,N_645,N_107);
or U1806 (N_1806,N_756,N_484);
nand U1807 (N_1807,N_663,N_156);
and U1808 (N_1808,N_430,N_822);
xnor U1809 (N_1809,N_143,N_834);
and U1810 (N_1810,N_811,N_105);
or U1811 (N_1811,N_507,N_212);
xor U1812 (N_1812,N_897,N_879);
or U1813 (N_1813,N_191,N_814);
nand U1814 (N_1814,N_576,N_712);
nor U1815 (N_1815,N_161,N_941);
and U1816 (N_1816,N_562,N_366);
or U1817 (N_1817,N_711,N_188);
or U1818 (N_1818,N_747,N_752);
nor U1819 (N_1819,N_791,N_522);
nand U1820 (N_1820,N_237,N_723);
nor U1821 (N_1821,N_195,N_263);
or U1822 (N_1822,N_829,N_569);
nand U1823 (N_1823,N_386,N_504);
nand U1824 (N_1824,N_352,N_763);
xor U1825 (N_1825,N_455,N_822);
nand U1826 (N_1826,N_288,N_907);
nand U1827 (N_1827,N_470,N_274);
or U1828 (N_1828,N_557,N_137);
and U1829 (N_1829,N_512,N_851);
nand U1830 (N_1830,N_137,N_938);
xnor U1831 (N_1831,N_215,N_284);
nor U1832 (N_1832,N_826,N_302);
and U1833 (N_1833,N_533,N_266);
xor U1834 (N_1834,N_127,N_70);
nor U1835 (N_1835,N_243,N_868);
nand U1836 (N_1836,N_355,N_718);
and U1837 (N_1837,N_578,N_738);
nand U1838 (N_1838,N_2,N_800);
nor U1839 (N_1839,N_303,N_21);
nand U1840 (N_1840,N_572,N_291);
and U1841 (N_1841,N_140,N_34);
or U1842 (N_1842,N_898,N_752);
xnor U1843 (N_1843,N_348,N_742);
and U1844 (N_1844,N_725,N_233);
nor U1845 (N_1845,N_394,N_259);
nor U1846 (N_1846,N_117,N_130);
nor U1847 (N_1847,N_463,N_651);
xor U1848 (N_1848,N_83,N_784);
nand U1849 (N_1849,N_79,N_329);
and U1850 (N_1850,N_255,N_77);
nor U1851 (N_1851,N_973,N_29);
or U1852 (N_1852,N_46,N_131);
nand U1853 (N_1853,N_616,N_756);
or U1854 (N_1854,N_207,N_2);
nor U1855 (N_1855,N_767,N_734);
nand U1856 (N_1856,N_265,N_211);
nor U1857 (N_1857,N_218,N_825);
nand U1858 (N_1858,N_28,N_397);
nand U1859 (N_1859,N_63,N_597);
xnor U1860 (N_1860,N_228,N_157);
or U1861 (N_1861,N_208,N_786);
or U1862 (N_1862,N_710,N_227);
nand U1863 (N_1863,N_32,N_470);
and U1864 (N_1864,N_826,N_558);
nor U1865 (N_1865,N_929,N_750);
nand U1866 (N_1866,N_428,N_588);
nor U1867 (N_1867,N_15,N_493);
nand U1868 (N_1868,N_730,N_51);
nand U1869 (N_1869,N_801,N_323);
nand U1870 (N_1870,N_434,N_48);
xor U1871 (N_1871,N_538,N_324);
xor U1872 (N_1872,N_317,N_835);
and U1873 (N_1873,N_190,N_707);
xnor U1874 (N_1874,N_608,N_731);
nor U1875 (N_1875,N_203,N_977);
or U1876 (N_1876,N_461,N_530);
nand U1877 (N_1877,N_80,N_106);
nor U1878 (N_1878,N_830,N_507);
nand U1879 (N_1879,N_941,N_185);
or U1880 (N_1880,N_297,N_767);
nand U1881 (N_1881,N_696,N_710);
and U1882 (N_1882,N_54,N_258);
nand U1883 (N_1883,N_321,N_144);
nor U1884 (N_1884,N_85,N_921);
nand U1885 (N_1885,N_496,N_992);
and U1886 (N_1886,N_497,N_283);
or U1887 (N_1887,N_712,N_653);
nor U1888 (N_1888,N_300,N_106);
and U1889 (N_1889,N_83,N_303);
nand U1890 (N_1890,N_889,N_634);
or U1891 (N_1891,N_927,N_742);
nor U1892 (N_1892,N_399,N_863);
and U1893 (N_1893,N_586,N_811);
or U1894 (N_1894,N_241,N_645);
nand U1895 (N_1895,N_24,N_847);
nor U1896 (N_1896,N_273,N_887);
and U1897 (N_1897,N_502,N_421);
or U1898 (N_1898,N_694,N_633);
or U1899 (N_1899,N_118,N_583);
and U1900 (N_1900,N_340,N_127);
nor U1901 (N_1901,N_662,N_428);
or U1902 (N_1902,N_189,N_840);
or U1903 (N_1903,N_200,N_121);
or U1904 (N_1904,N_152,N_837);
and U1905 (N_1905,N_722,N_403);
xnor U1906 (N_1906,N_689,N_473);
nor U1907 (N_1907,N_809,N_418);
or U1908 (N_1908,N_275,N_677);
xnor U1909 (N_1909,N_302,N_981);
nor U1910 (N_1910,N_382,N_353);
nand U1911 (N_1911,N_116,N_307);
nor U1912 (N_1912,N_804,N_10);
or U1913 (N_1913,N_544,N_419);
nor U1914 (N_1914,N_410,N_156);
xnor U1915 (N_1915,N_409,N_837);
and U1916 (N_1916,N_302,N_470);
nor U1917 (N_1917,N_493,N_229);
nand U1918 (N_1918,N_130,N_528);
and U1919 (N_1919,N_148,N_9);
nand U1920 (N_1920,N_452,N_825);
and U1921 (N_1921,N_623,N_545);
and U1922 (N_1922,N_31,N_753);
xor U1923 (N_1923,N_192,N_326);
nand U1924 (N_1924,N_50,N_235);
and U1925 (N_1925,N_816,N_664);
or U1926 (N_1926,N_942,N_623);
and U1927 (N_1927,N_424,N_174);
nor U1928 (N_1928,N_50,N_795);
nand U1929 (N_1929,N_646,N_28);
and U1930 (N_1930,N_158,N_15);
nand U1931 (N_1931,N_231,N_762);
xor U1932 (N_1932,N_448,N_406);
and U1933 (N_1933,N_143,N_366);
nand U1934 (N_1934,N_405,N_523);
xnor U1935 (N_1935,N_284,N_687);
nor U1936 (N_1936,N_583,N_946);
nor U1937 (N_1937,N_146,N_247);
or U1938 (N_1938,N_980,N_127);
and U1939 (N_1939,N_95,N_814);
xnor U1940 (N_1940,N_868,N_337);
and U1941 (N_1941,N_589,N_591);
and U1942 (N_1942,N_896,N_259);
and U1943 (N_1943,N_744,N_645);
nor U1944 (N_1944,N_97,N_409);
and U1945 (N_1945,N_186,N_304);
nor U1946 (N_1946,N_158,N_246);
nand U1947 (N_1947,N_350,N_874);
xnor U1948 (N_1948,N_501,N_688);
nor U1949 (N_1949,N_906,N_864);
or U1950 (N_1950,N_541,N_693);
and U1951 (N_1951,N_551,N_36);
or U1952 (N_1952,N_269,N_832);
or U1953 (N_1953,N_728,N_576);
xor U1954 (N_1954,N_488,N_483);
or U1955 (N_1955,N_645,N_782);
xor U1956 (N_1956,N_763,N_286);
or U1957 (N_1957,N_566,N_777);
or U1958 (N_1958,N_210,N_404);
nor U1959 (N_1959,N_965,N_588);
or U1960 (N_1960,N_432,N_887);
nand U1961 (N_1961,N_863,N_559);
or U1962 (N_1962,N_517,N_112);
or U1963 (N_1963,N_94,N_460);
nand U1964 (N_1964,N_244,N_703);
xor U1965 (N_1965,N_986,N_694);
nor U1966 (N_1966,N_60,N_850);
and U1967 (N_1967,N_697,N_993);
and U1968 (N_1968,N_702,N_40);
and U1969 (N_1969,N_348,N_513);
or U1970 (N_1970,N_631,N_347);
nor U1971 (N_1971,N_946,N_413);
nand U1972 (N_1972,N_21,N_595);
nand U1973 (N_1973,N_355,N_849);
and U1974 (N_1974,N_982,N_643);
nor U1975 (N_1975,N_914,N_231);
nor U1976 (N_1976,N_502,N_619);
or U1977 (N_1977,N_649,N_955);
or U1978 (N_1978,N_873,N_474);
nor U1979 (N_1979,N_850,N_891);
xor U1980 (N_1980,N_87,N_233);
nand U1981 (N_1981,N_832,N_290);
nand U1982 (N_1982,N_128,N_196);
and U1983 (N_1983,N_77,N_555);
nand U1984 (N_1984,N_723,N_920);
and U1985 (N_1985,N_816,N_805);
and U1986 (N_1986,N_825,N_99);
or U1987 (N_1987,N_852,N_991);
and U1988 (N_1988,N_827,N_187);
and U1989 (N_1989,N_205,N_343);
or U1990 (N_1990,N_17,N_42);
or U1991 (N_1991,N_515,N_961);
or U1992 (N_1992,N_125,N_97);
or U1993 (N_1993,N_678,N_723);
xnor U1994 (N_1994,N_22,N_177);
xnor U1995 (N_1995,N_523,N_415);
or U1996 (N_1996,N_975,N_390);
xnor U1997 (N_1997,N_196,N_890);
nand U1998 (N_1998,N_140,N_705);
nor U1999 (N_1999,N_373,N_914);
and U2000 (N_2000,N_1874,N_1420);
or U2001 (N_2001,N_1077,N_1649);
nor U2002 (N_2002,N_1114,N_1111);
and U2003 (N_2003,N_1486,N_1873);
nand U2004 (N_2004,N_1431,N_1623);
xnor U2005 (N_2005,N_1367,N_1499);
xor U2006 (N_2006,N_1476,N_1036);
nand U2007 (N_2007,N_1883,N_1277);
nor U2008 (N_2008,N_1030,N_1598);
nand U2009 (N_2009,N_1457,N_1738);
xor U2010 (N_2010,N_1854,N_1353);
nor U2011 (N_2011,N_1311,N_1388);
or U2012 (N_2012,N_1703,N_1063);
nor U2013 (N_2013,N_1797,N_1449);
xnor U2014 (N_2014,N_1684,N_1344);
or U2015 (N_2015,N_1740,N_1565);
and U2016 (N_2016,N_1328,N_1024);
nor U2017 (N_2017,N_1378,N_1671);
nor U2018 (N_2018,N_1660,N_1133);
nor U2019 (N_2019,N_1336,N_1628);
or U2020 (N_2020,N_1710,N_1257);
or U2021 (N_2021,N_1340,N_1936);
xnor U2022 (N_2022,N_1472,N_1366);
and U2023 (N_2023,N_1553,N_1548);
nand U2024 (N_2024,N_1039,N_1924);
xor U2025 (N_2025,N_1374,N_1363);
or U2026 (N_2026,N_1739,N_1821);
or U2027 (N_2027,N_1405,N_1183);
xnor U2028 (N_2028,N_1426,N_1347);
nand U2029 (N_2029,N_1653,N_1530);
nand U2030 (N_2030,N_1622,N_1935);
nand U2031 (N_2031,N_1611,N_1162);
nor U2032 (N_2032,N_1748,N_1147);
xor U2033 (N_2033,N_1569,N_1325);
or U2034 (N_2034,N_1369,N_1690);
nor U2035 (N_2035,N_1411,N_1656);
or U2036 (N_2036,N_1142,N_1828);
or U2037 (N_2037,N_1872,N_1759);
nor U2038 (N_2038,N_1349,N_1465);
xor U2039 (N_2039,N_1931,N_1364);
nand U2040 (N_2040,N_1331,N_1817);
or U2041 (N_2041,N_1721,N_1644);
xor U2042 (N_2042,N_1217,N_1758);
nor U2043 (N_2043,N_1497,N_1942);
nor U2044 (N_2044,N_1826,N_1729);
xnor U2045 (N_2045,N_1483,N_1932);
nor U2046 (N_2046,N_1238,N_1168);
xnor U2047 (N_2047,N_1899,N_1085);
and U2048 (N_2048,N_1595,N_1749);
nand U2049 (N_2049,N_1824,N_1144);
and U2050 (N_2050,N_1993,N_1679);
nand U2051 (N_2051,N_1042,N_1596);
and U2052 (N_2052,N_1626,N_1507);
and U2053 (N_2053,N_1638,N_1469);
xnor U2054 (N_2054,N_1723,N_1506);
nand U2055 (N_2055,N_1919,N_1757);
nand U2056 (N_2056,N_1037,N_1381);
xnor U2057 (N_2057,N_1475,N_1377);
and U2058 (N_2058,N_1260,N_1308);
nor U2059 (N_2059,N_1876,N_1365);
nand U2060 (N_2060,N_1953,N_1341);
nor U2061 (N_2061,N_1354,N_1053);
xnor U2062 (N_2062,N_1021,N_1323);
nand U2063 (N_2063,N_1035,N_1819);
and U2064 (N_2064,N_1445,N_1988);
nor U2065 (N_2065,N_1361,N_1470);
or U2066 (N_2066,N_1514,N_1525);
and U2067 (N_2067,N_1187,N_1337);
and U2068 (N_2068,N_1072,N_1555);
and U2069 (N_2069,N_1808,N_1359);
and U2070 (N_2070,N_1563,N_1327);
nand U2071 (N_2071,N_1098,N_1101);
and U2072 (N_2072,N_1802,N_1895);
nand U2073 (N_2073,N_1847,N_1067);
or U2074 (N_2074,N_1853,N_1273);
xor U2075 (N_2075,N_1552,N_1448);
xor U2076 (N_2076,N_1262,N_1446);
nand U2077 (N_2077,N_1214,N_1702);
xnor U2078 (N_2078,N_1040,N_1665);
nand U2079 (N_2079,N_1103,N_1813);
nor U2080 (N_2080,N_1708,N_1677);
xnor U2081 (N_2081,N_1857,N_1003);
nor U2082 (N_2082,N_1334,N_1655);
and U2083 (N_2083,N_1915,N_1652);
or U2084 (N_2084,N_1602,N_1494);
nand U2085 (N_2085,N_1706,N_1482);
xnor U2086 (N_2086,N_1265,N_1081);
or U2087 (N_2087,N_1401,N_1864);
nand U2088 (N_2088,N_1750,N_1298);
and U2089 (N_2089,N_1135,N_1699);
nor U2090 (N_2090,N_1001,N_1385);
nand U2091 (N_2091,N_1302,N_1430);
and U2092 (N_2092,N_1952,N_1523);
or U2093 (N_2093,N_1767,N_1437);
nor U2094 (N_2094,N_1458,N_1176);
nand U2095 (N_2095,N_1301,N_1267);
or U2096 (N_2096,N_1515,N_1230);
nor U2097 (N_2097,N_1734,N_1146);
nor U2098 (N_2098,N_1784,N_1222);
nor U2099 (N_2099,N_1118,N_1186);
or U2100 (N_2100,N_1989,N_1627);
or U2101 (N_2101,N_1505,N_1856);
xor U2102 (N_2102,N_1779,N_1316);
or U2103 (N_2103,N_1259,N_1068);
and U2104 (N_2104,N_1551,N_1810);
or U2105 (N_2105,N_1643,N_1544);
and U2106 (N_2106,N_1180,N_1687);
or U2107 (N_2107,N_1400,N_1827);
nor U2108 (N_2108,N_1455,N_1329);
xnor U2109 (N_2109,N_1669,N_1080);
or U2110 (N_2110,N_1194,N_1235);
and U2111 (N_2111,N_1283,N_1502);
nor U2112 (N_2112,N_1079,N_1295);
and U2113 (N_2113,N_1865,N_1519);
and U2114 (N_2114,N_1579,N_1435);
or U2115 (N_2115,N_1433,N_1124);
or U2116 (N_2116,N_1838,N_1536);
xor U2117 (N_2117,N_1674,N_1616);
or U2118 (N_2118,N_1165,N_1885);
nor U2119 (N_2119,N_1126,N_1440);
xor U2120 (N_2120,N_1982,N_1450);
xnor U2121 (N_2121,N_1913,N_1417);
xnor U2122 (N_2122,N_1140,N_1641);
or U2123 (N_2123,N_1689,N_1766);
xnor U2124 (N_2124,N_1834,N_1558);
or U2125 (N_2125,N_1120,N_1276);
or U2126 (N_2126,N_1646,N_1790);
nor U2127 (N_2127,N_1123,N_1956);
nand U2128 (N_2128,N_1585,N_1675);
nand U2129 (N_2129,N_1795,N_1383);
or U2130 (N_2130,N_1402,N_1948);
nand U2131 (N_2131,N_1460,N_1179);
and U2132 (N_2132,N_1275,N_1752);
nor U2133 (N_2133,N_1692,N_1861);
xor U2134 (N_2134,N_1593,N_1882);
or U2135 (N_2135,N_1521,N_1312);
and U2136 (N_2136,N_1203,N_1288);
nor U2137 (N_2137,N_1645,N_1540);
and U2138 (N_2138,N_1352,N_1709);
nand U2139 (N_2139,N_1228,N_1816);
or U2140 (N_2140,N_1468,N_1207);
nor U2141 (N_2141,N_1946,N_1736);
xnor U2142 (N_2142,N_1875,N_1054);
nand U2143 (N_2143,N_1326,N_1958);
and U2144 (N_2144,N_1518,N_1095);
or U2145 (N_2145,N_1831,N_1373);
or U2146 (N_2146,N_1017,N_1539);
or U2147 (N_2147,N_1389,N_1537);
nand U2148 (N_2148,N_1157,N_1822);
or U2149 (N_2149,N_1052,N_1439);
nor U2150 (N_2150,N_1412,N_1392);
nand U2151 (N_2151,N_1572,N_1108);
nand U2152 (N_2152,N_1914,N_1704);
and U2153 (N_2153,N_1282,N_1905);
and U2154 (N_2154,N_1884,N_1866);
nor U2155 (N_2155,N_1911,N_1093);
xor U2156 (N_2156,N_1076,N_1125);
nor U2157 (N_2157,N_1733,N_1934);
nand U2158 (N_2158,N_1681,N_1964);
xnor U2159 (N_2159,N_1406,N_1303);
nor U2160 (N_2160,N_1557,N_1229);
nor U2161 (N_2161,N_1529,N_1473);
nor U2162 (N_2162,N_1432,N_1787);
and U2163 (N_2163,N_1212,N_1453);
nand U2164 (N_2164,N_1169,N_1799);
nand U2165 (N_2165,N_1501,N_1517);
nor U2166 (N_2166,N_1945,N_1693);
or U2167 (N_2167,N_1160,N_1588);
or U2168 (N_2168,N_1429,N_1310);
nor U2169 (N_2169,N_1916,N_1570);
nor U2170 (N_2170,N_1741,N_1727);
or U2171 (N_2171,N_1069,N_1711);
xor U2172 (N_2172,N_1609,N_1564);
nand U2173 (N_2173,N_1726,N_1320);
xor U2174 (N_2174,N_1843,N_1143);
nand U2175 (N_2175,N_1929,N_1603);
nand U2176 (N_2176,N_1859,N_1688);
nand U2177 (N_2177,N_1754,N_1705);
nand U2178 (N_2178,N_1666,N_1744);
or U2179 (N_2179,N_1995,N_1683);
and U2180 (N_2180,N_1601,N_1906);
xor U2181 (N_2181,N_1116,N_1263);
xnor U2182 (N_2182,N_1720,N_1425);
and U2183 (N_2183,N_1503,N_1390);
nor U2184 (N_2184,N_1893,N_1663);
nor U2185 (N_2185,N_1041,N_1901);
nor U2186 (N_2186,N_1992,N_1747);
xor U2187 (N_2187,N_1015,N_1393);
xor U2188 (N_2188,N_1296,N_1031);
nand U2189 (N_2189,N_1100,N_1038);
xor U2190 (N_2190,N_1131,N_1793);
and U2191 (N_2191,N_1066,N_1490);
or U2192 (N_2192,N_1966,N_1657);
nor U2193 (N_2193,N_1957,N_1839);
and U2194 (N_2194,N_1981,N_1286);
or U2195 (N_2195,N_1300,N_1918);
nand U2196 (N_2196,N_1780,N_1044);
and U2197 (N_2197,N_1785,N_1668);
nor U2198 (N_2198,N_1962,N_1614);
nand U2199 (N_2199,N_1877,N_1809);
nor U2200 (N_2200,N_1200,N_1184);
or U2201 (N_2201,N_1737,N_1771);
nand U2202 (N_2202,N_1322,N_1315);
nor U2203 (N_2203,N_1249,N_1670);
nor U2204 (N_2204,N_1892,N_1023);
or U2205 (N_2205,N_1608,N_1535);
nor U2206 (N_2206,N_1491,N_1065);
nand U2207 (N_2207,N_1561,N_1836);
xnor U2208 (N_2208,N_1049,N_1285);
xnor U2209 (N_2209,N_1753,N_1145);
or U2210 (N_2210,N_1830,N_1567);
and U2211 (N_2211,N_1937,N_1778);
xor U2212 (N_2212,N_1951,N_1922);
xnor U2213 (N_2213,N_1156,N_1129);
nor U2214 (N_2214,N_1648,N_1208);
nand U2215 (N_2215,N_1404,N_1423);
nor U2216 (N_2216,N_1890,N_1092);
nor U2217 (N_2217,N_1541,N_1342);
or U2218 (N_2218,N_1545,N_1855);
nor U2219 (N_2219,N_1173,N_1481);
nor U2220 (N_2220,N_1421,N_1121);
and U2221 (N_2221,N_1575,N_1020);
nor U2222 (N_2222,N_1188,N_1223);
xor U2223 (N_2223,N_1474,N_1635);
nor U2224 (N_2224,N_1013,N_1731);
or U2225 (N_2225,N_1624,N_1697);
nor U2226 (N_2226,N_1636,N_1532);
and U2227 (N_2227,N_1508,N_1250);
nor U2228 (N_2228,N_1625,N_1584);
xnor U2229 (N_2229,N_1141,N_1175);
and U2230 (N_2230,N_1651,N_1968);
xor U2231 (N_2231,N_1938,N_1343);
nand U2232 (N_2232,N_1471,N_1255);
xor U2233 (N_2233,N_1464,N_1451);
and U2234 (N_2234,N_1858,N_1005);
nor U2235 (N_2235,N_1461,N_1926);
xor U2236 (N_2236,N_1027,N_1436);
nand U2237 (N_2237,N_1161,N_1048);
nor U2238 (N_2238,N_1770,N_1271);
xor U2239 (N_2239,N_1713,N_1806);
or U2240 (N_2240,N_1742,N_1008);
nor U2241 (N_2241,N_1479,N_1191);
nand U2242 (N_2242,N_1871,N_1586);
nand U2243 (N_2243,N_1197,N_1484);
nor U2244 (N_2244,N_1533,N_1985);
nand U2245 (N_2245,N_1969,N_1763);
xor U2246 (N_2246,N_1413,N_1115);
or U2247 (N_2247,N_1061,N_1820);
or U2248 (N_2248,N_1216,N_1047);
xnor U2249 (N_2249,N_1278,N_1746);
and U2250 (N_2250,N_1084,N_1456);
nand U2251 (N_2251,N_1332,N_1801);
nand U2252 (N_2252,N_1279,N_1234);
nand U2253 (N_2253,N_1415,N_1632);
or U2254 (N_2254,N_1358,N_1132);
and U2255 (N_2255,N_1304,N_1338);
and U2256 (N_2256,N_1012,N_1606);
or U2257 (N_2257,N_1199,N_1504);
nand U2258 (N_2258,N_1888,N_1137);
or U2259 (N_2259,N_1351,N_1236);
and U2260 (N_2260,N_1886,N_1438);
nor U2261 (N_2261,N_1781,N_1904);
nand U2262 (N_2262,N_1130,N_1794);
nand U2263 (N_2263,N_1983,N_1167);
and U2264 (N_2264,N_1219,N_1500);
or U2265 (N_2265,N_1324,N_1270);
nand U2266 (N_2266,N_1807,N_1833);
or U2267 (N_2267,N_1231,N_1792);
or U2268 (N_2268,N_1164,N_1357);
nand U2269 (N_2269,N_1493,N_1025);
and U2270 (N_2270,N_1512,N_1607);
nand U2271 (N_2271,N_1452,N_1835);
and U2272 (N_2272,N_1573,N_1716);
nand U2273 (N_2273,N_1202,N_1462);
xor U2274 (N_2274,N_1718,N_1695);
and U2275 (N_2275,N_1192,N_1292);
nand U2276 (N_2276,N_1016,N_1057);
or U2277 (N_2277,N_1396,N_1371);
nor U2278 (N_2278,N_1756,N_1495);
nor U2279 (N_2279,N_1158,N_1339);
and U2280 (N_2280,N_1127,N_1087);
or U2281 (N_2281,N_1391,N_1587);
or U2282 (N_2282,N_1014,N_1743);
or U2283 (N_2283,N_1676,N_1867);
and U2284 (N_2284,N_1818,N_1189);
nor U2285 (N_2285,N_1765,N_1086);
nand U2286 (N_2286,N_1549,N_1345);
or U2287 (N_2287,N_1944,N_1940);
and U2288 (N_2288,N_1496,N_1617);
xor U2289 (N_2289,N_1247,N_1590);
xor U2290 (N_2290,N_1917,N_1428);
xor U2291 (N_2291,N_1712,N_1696);
nand U2292 (N_2292,N_1583,N_1064);
or U2293 (N_2293,N_1955,N_1097);
nor U2294 (N_2294,N_1242,N_1782);
nand U2295 (N_2295,N_1463,N_1350);
nand U2296 (N_2296,N_1900,N_1399);
nand U2297 (N_2297,N_1788,N_1630);
nor U2298 (N_2298,N_1868,N_1618);
nor U2299 (N_2299,N_1928,N_1898);
and U2300 (N_2300,N_1987,N_1933);
nand U2301 (N_2301,N_1629,N_1051);
xor U2302 (N_2302,N_1775,N_1070);
nor U2303 (N_2303,N_1386,N_1485);
nor U2304 (N_2304,N_1848,N_1984);
and U2305 (N_2305,N_1408,N_1007);
nand U2306 (N_2306,N_1290,N_1999);
and U2307 (N_2307,N_1447,N_1177);
nand U2308 (N_2308,N_1730,N_1949);
xor U2309 (N_2309,N_1849,N_1119);
xor U2310 (N_2310,N_1566,N_1082);
xnor U2311 (N_2311,N_1789,N_1233);
or U2312 (N_2312,N_1978,N_1498);
nand U2313 (N_2313,N_1979,N_1812);
xnor U2314 (N_2314,N_1870,N_1961);
nand U2315 (N_2315,N_1823,N_1224);
and U2316 (N_2316,N_1409,N_1209);
and U2317 (N_2317,N_1215,N_1105);
or U2318 (N_2318,N_1043,N_1174);
and U2319 (N_2319,N_1612,N_1894);
nor U2320 (N_2320,N_1582,N_1317);
nor U2321 (N_2321,N_1193,N_1280);
or U2322 (N_2322,N_1370,N_1912);
nand U2323 (N_2323,N_1717,N_1891);
and U2324 (N_2324,N_1443,N_1434);
nor U2325 (N_2325,N_1592,N_1254);
nor U2326 (N_2326,N_1073,N_1520);
or U2327 (N_2327,N_1970,N_1467);
and U2328 (N_2328,N_1996,N_1136);
nand U2329 (N_2329,N_1634,N_1150);
xnor U2330 (N_2330,N_1029,N_1113);
nand U2331 (N_2331,N_1416,N_1246);
nor U2332 (N_2332,N_1889,N_1510);
nand U2333 (N_2333,N_1407,N_1289);
nor U2334 (N_2334,N_1805,N_1600);
xor U2335 (N_2335,N_1394,N_1783);
or U2336 (N_2336,N_1099,N_1480);
xor U2337 (N_2337,N_1562,N_1526);
nor U2338 (N_2338,N_1777,N_1967);
nand U2339 (N_2339,N_1205,N_1376);
xor U2340 (N_2340,N_1441,N_1554);
and U2341 (N_2341,N_1910,N_1550);
nand U2342 (N_2342,N_1639,N_1959);
nor U2343 (N_2343,N_1678,N_1825);
xnor U2344 (N_2344,N_1163,N_1221);
nor U2345 (N_2345,N_1045,N_1346);
nand U2346 (N_2346,N_1903,N_1897);
or U2347 (N_2347,N_1581,N_1348);
or U2348 (N_2348,N_1306,N_1239);
nor U2349 (N_2349,N_1387,N_1004);
nor U2350 (N_2350,N_1691,N_1605);
and U2351 (N_2351,N_1841,N_1640);
or U2352 (N_2352,N_1686,N_1281);
nand U2353 (N_2353,N_1963,N_1509);
nor U2354 (N_2354,N_1154,N_1800);
xnor U2355 (N_2355,N_1033,N_1002);
and U2356 (N_2356,N_1459,N_1796);
nand U2357 (N_2357,N_1355,N_1732);
or U2358 (N_2358,N_1642,N_1574);
and U2359 (N_2359,N_1769,N_1368);
xor U2360 (N_2360,N_1685,N_1925);
nor U2361 (N_2361,N_1589,N_1719);
or U2362 (N_2362,N_1975,N_1102);
nor U2363 (N_2363,N_1701,N_1577);
nor U2364 (N_2364,N_1424,N_1243);
nor U2365 (N_2365,N_1284,N_1244);
nor U2366 (N_2366,N_1735,N_1815);
and U2367 (N_2367,N_1994,N_1560);
and U2368 (N_2368,N_1965,N_1028);
nand U2369 (N_2369,N_1707,N_1990);
xnor U2370 (N_2370,N_1804,N_1226);
and U2371 (N_2371,N_1335,N_1397);
or U2372 (N_2372,N_1921,N_1106);
nor U2373 (N_2373,N_1578,N_1264);
nor U2374 (N_2374,N_1724,N_1427);
xnor U2375 (N_2375,N_1599,N_1591);
nor U2376 (N_2376,N_1321,N_1291);
nor U2377 (N_2377,N_1006,N_1211);
and U2378 (N_2378,N_1009,N_1832);
or U2379 (N_2379,N_1261,N_1682);
xnor U2380 (N_2380,N_1680,N_1330);
nor U2381 (N_2381,N_1728,N_1973);
nor U2382 (N_2382,N_1094,N_1878);
nor U2383 (N_2383,N_1151,N_1225);
nor U2384 (N_2384,N_1362,N_1232);
or U2385 (N_2385,N_1869,N_1309);
or U2386 (N_2386,N_1487,N_1516);
nor U2387 (N_2387,N_1851,N_1091);
nor U2388 (N_2388,N_1182,N_1714);
or U2389 (N_2389,N_1148,N_1220);
and U2390 (N_2390,N_1972,N_1059);
nand U2391 (N_2391,N_1814,N_1576);
nand U2392 (N_2392,N_1379,N_1803);
xor U2393 (N_2393,N_1178,N_1166);
nor U2394 (N_2394,N_1908,N_1213);
nand U2395 (N_2395,N_1319,N_1647);
or U2396 (N_2396,N_1527,N_1954);
nor U2397 (N_2397,N_1772,N_1662);
nor U2398 (N_2398,N_1542,N_1543);
nand U2399 (N_2399,N_1258,N_1032);
and U2400 (N_2400,N_1372,N_1110);
or U2401 (N_2401,N_1923,N_1986);
and U2402 (N_2402,N_1422,N_1943);
and U2403 (N_2403,N_1395,N_1997);
and U2404 (N_2404,N_1976,N_1109);
nor U2405 (N_2405,N_1088,N_1251);
or U2406 (N_2406,N_1305,N_1410);
xor U2407 (N_2407,N_1930,N_1019);
or U2408 (N_2408,N_1253,N_1297);
and U2409 (N_2409,N_1190,N_1171);
or U2410 (N_2410,N_1356,N_1907);
nand U2411 (N_2411,N_1725,N_1050);
and U2412 (N_2412,N_1844,N_1631);
nor U2413 (N_2413,N_1149,N_1773);
and U2414 (N_2414,N_1237,N_1206);
nor U2415 (N_2415,N_1571,N_1654);
xor U2416 (N_2416,N_1971,N_1248);
xor U2417 (N_2417,N_1000,N_1774);
and U2418 (N_2418,N_1768,N_1062);
nand U2419 (N_2419,N_1266,N_1980);
xor U2420 (N_2420,N_1700,N_1299);
nand U2421 (N_2421,N_1010,N_1074);
or U2422 (N_2422,N_1333,N_1418);
or U2423 (N_2423,N_1139,N_1998);
nand U2424 (N_2424,N_1947,N_1829);
nor U2425 (N_2425,N_1172,N_1538);
and U2426 (N_2426,N_1466,N_1198);
xor U2427 (N_2427,N_1667,N_1974);
nand U2428 (N_2428,N_1559,N_1185);
xor U2429 (N_2429,N_1078,N_1011);
xor U2430 (N_2430,N_1414,N_1960);
and U2431 (N_2431,N_1531,N_1477);
nand U2432 (N_2432,N_1293,N_1107);
nor U2433 (N_2433,N_1026,N_1056);
or U2434 (N_2434,N_1478,N_1977);
xor U2435 (N_2435,N_1274,N_1811);
xnor U2436 (N_2436,N_1664,N_1096);
xor U2437 (N_2437,N_1615,N_1619);
nand U2438 (N_2438,N_1715,N_1863);
nand U2439 (N_2439,N_1633,N_1318);
xnor U2440 (N_2440,N_1610,N_1384);
and U2441 (N_2441,N_1195,N_1294);
xor U2442 (N_2442,N_1661,N_1252);
xnor U2443 (N_2443,N_1227,N_1881);
xor U2444 (N_2444,N_1568,N_1360);
xor U2445 (N_2445,N_1138,N_1204);
and U2446 (N_2446,N_1240,N_1762);
nand U2447 (N_2447,N_1534,N_1950);
or U2448 (N_2448,N_1522,N_1798);
nand U2449 (N_2449,N_1307,N_1761);
nor U2450 (N_2450,N_1528,N_1659);
or U2451 (N_2451,N_1852,N_1287);
or U2452 (N_2452,N_1159,N_1313);
or U2453 (N_2453,N_1492,N_1489);
nor U2454 (N_2454,N_1419,N_1210);
and U2455 (N_2455,N_1786,N_1673);
nor U2456 (N_2456,N_1846,N_1488);
and U2457 (N_2457,N_1170,N_1071);
xnor U2458 (N_2458,N_1939,N_1860);
and U2459 (N_2459,N_1751,N_1128);
or U2460 (N_2460,N_1403,N_1850);
and U2461 (N_2461,N_1022,N_1201);
and U2462 (N_2462,N_1046,N_1060);
xor U2463 (N_2463,N_1269,N_1776);
nor U2464 (N_2464,N_1134,N_1650);
nand U2465 (N_2465,N_1546,N_1112);
nand U2466 (N_2466,N_1513,N_1941);
nand U2467 (N_2467,N_1382,N_1454);
and U2468 (N_2468,N_1837,N_1256);
xnor U2469 (N_2469,N_1694,N_1594);
xor U2470 (N_2470,N_1879,N_1845);
nand U2471 (N_2471,N_1547,N_1760);
or U2472 (N_2472,N_1055,N_1241);
nor U2473 (N_2473,N_1991,N_1380);
xor U2474 (N_2474,N_1880,N_1218);
nor U2475 (N_2475,N_1083,N_1637);
and U2476 (N_2476,N_1658,N_1613);
nand U2477 (N_2477,N_1524,N_1597);
xor U2478 (N_2478,N_1268,N_1755);
or U2479 (N_2479,N_1862,N_1920);
nor U2480 (N_2480,N_1621,N_1034);
or U2481 (N_2481,N_1117,N_1152);
or U2482 (N_2482,N_1375,N_1896);
or U2483 (N_2483,N_1196,N_1902);
nand U2484 (N_2484,N_1764,N_1089);
nand U2485 (N_2485,N_1580,N_1058);
nand U2486 (N_2486,N_1620,N_1887);
nand U2487 (N_2487,N_1604,N_1927);
nor U2488 (N_2488,N_1698,N_1075);
nand U2489 (N_2489,N_1745,N_1122);
or U2490 (N_2490,N_1090,N_1444);
and U2491 (N_2491,N_1791,N_1672);
xor U2492 (N_2492,N_1272,N_1840);
nand U2493 (N_2493,N_1155,N_1722);
xor U2494 (N_2494,N_1511,N_1181);
nand U2495 (N_2495,N_1245,N_1556);
xnor U2496 (N_2496,N_1442,N_1314);
nand U2497 (N_2497,N_1909,N_1018);
and U2498 (N_2498,N_1104,N_1153);
and U2499 (N_2499,N_1842,N_1398);
and U2500 (N_2500,N_1818,N_1597);
and U2501 (N_2501,N_1734,N_1429);
nand U2502 (N_2502,N_1795,N_1313);
nand U2503 (N_2503,N_1068,N_1410);
and U2504 (N_2504,N_1214,N_1780);
nand U2505 (N_2505,N_1068,N_1572);
xnor U2506 (N_2506,N_1791,N_1146);
xnor U2507 (N_2507,N_1519,N_1910);
or U2508 (N_2508,N_1515,N_1183);
nand U2509 (N_2509,N_1932,N_1387);
nor U2510 (N_2510,N_1160,N_1930);
or U2511 (N_2511,N_1142,N_1388);
nand U2512 (N_2512,N_1333,N_1980);
nand U2513 (N_2513,N_1068,N_1969);
or U2514 (N_2514,N_1560,N_1139);
nor U2515 (N_2515,N_1045,N_1185);
and U2516 (N_2516,N_1111,N_1809);
and U2517 (N_2517,N_1278,N_1826);
nor U2518 (N_2518,N_1423,N_1952);
and U2519 (N_2519,N_1015,N_1325);
or U2520 (N_2520,N_1958,N_1567);
xnor U2521 (N_2521,N_1054,N_1385);
xor U2522 (N_2522,N_1886,N_1851);
or U2523 (N_2523,N_1234,N_1276);
nand U2524 (N_2524,N_1970,N_1310);
nand U2525 (N_2525,N_1889,N_1506);
and U2526 (N_2526,N_1231,N_1489);
xor U2527 (N_2527,N_1533,N_1277);
and U2528 (N_2528,N_1600,N_1393);
and U2529 (N_2529,N_1015,N_1994);
nand U2530 (N_2530,N_1553,N_1277);
nand U2531 (N_2531,N_1222,N_1833);
and U2532 (N_2532,N_1727,N_1759);
xnor U2533 (N_2533,N_1028,N_1404);
xnor U2534 (N_2534,N_1724,N_1633);
and U2535 (N_2535,N_1726,N_1274);
xnor U2536 (N_2536,N_1141,N_1142);
nor U2537 (N_2537,N_1996,N_1695);
xor U2538 (N_2538,N_1128,N_1151);
or U2539 (N_2539,N_1539,N_1701);
or U2540 (N_2540,N_1934,N_1439);
nor U2541 (N_2541,N_1568,N_1071);
xor U2542 (N_2542,N_1979,N_1936);
and U2543 (N_2543,N_1015,N_1993);
nand U2544 (N_2544,N_1204,N_1524);
or U2545 (N_2545,N_1744,N_1147);
xor U2546 (N_2546,N_1244,N_1328);
or U2547 (N_2547,N_1892,N_1300);
or U2548 (N_2548,N_1109,N_1076);
xor U2549 (N_2549,N_1050,N_1849);
or U2550 (N_2550,N_1644,N_1120);
nor U2551 (N_2551,N_1233,N_1363);
nand U2552 (N_2552,N_1255,N_1869);
or U2553 (N_2553,N_1093,N_1891);
and U2554 (N_2554,N_1104,N_1226);
and U2555 (N_2555,N_1436,N_1100);
nand U2556 (N_2556,N_1088,N_1776);
xor U2557 (N_2557,N_1948,N_1972);
nor U2558 (N_2558,N_1803,N_1318);
xnor U2559 (N_2559,N_1297,N_1578);
xor U2560 (N_2560,N_1409,N_1728);
or U2561 (N_2561,N_1228,N_1245);
nand U2562 (N_2562,N_1244,N_1841);
xnor U2563 (N_2563,N_1946,N_1701);
and U2564 (N_2564,N_1366,N_1686);
nor U2565 (N_2565,N_1908,N_1551);
xor U2566 (N_2566,N_1549,N_1264);
nor U2567 (N_2567,N_1098,N_1613);
xor U2568 (N_2568,N_1787,N_1382);
and U2569 (N_2569,N_1115,N_1507);
xnor U2570 (N_2570,N_1277,N_1733);
nand U2571 (N_2571,N_1631,N_1641);
nor U2572 (N_2572,N_1942,N_1430);
or U2573 (N_2573,N_1776,N_1844);
nor U2574 (N_2574,N_1240,N_1650);
nand U2575 (N_2575,N_1370,N_1230);
nor U2576 (N_2576,N_1267,N_1181);
and U2577 (N_2577,N_1860,N_1471);
nand U2578 (N_2578,N_1121,N_1826);
nand U2579 (N_2579,N_1947,N_1683);
nand U2580 (N_2580,N_1185,N_1291);
nor U2581 (N_2581,N_1180,N_1143);
xnor U2582 (N_2582,N_1398,N_1504);
nand U2583 (N_2583,N_1220,N_1072);
and U2584 (N_2584,N_1101,N_1543);
or U2585 (N_2585,N_1391,N_1845);
nor U2586 (N_2586,N_1604,N_1898);
and U2587 (N_2587,N_1603,N_1200);
xnor U2588 (N_2588,N_1744,N_1938);
nor U2589 (N_2589,N_1211,N_1625);
or U2590 (N_2590,N_1722,N_1807);
nand U2591 (N_2591,N_1287,N_1631);
xor U2592 (N_2592,N_1830,N_1307);
nand U2593 (N_2593,N_1919,N_1230);
or U2594 (N_2594,N_1607,N_1931);
and U2595 (N_2595,N_1675,N_1674);
nor U2596 (N_2596,N_1401,N_1676);
or U2597 (N_2597,N_1995,N_1717);
and U2598 (N_2598,N_1580,N_1994);
or U2599 (N_2599,N_1400,N_1863);
xnor U2600 (N_2600,N_1689,N_1531);
xnor U2601 (N_2601,N_1439,N_1111);
and U2602 (N_2602,N_1337,N_1450);
nand U2603 (N_2603,N_1539,N_1506);
nand U2604 (N_2604,N_1844,N_1887);
nand U2605 (N_2605,N_1574,N_1379);
and U2606 (N_2606,N_1298,N_1973);
nor U2607 (N_2607,N_1032,N_1449);
and U2608 (N_2608,N_1165,N_1065);
and U2609 (N_2609,N_1359,N_1780);
and U2610 (N_2610,N_1648,N_1124);
nor U2611 (N_2611,N_1627,N_1988);
or U2612 (N_2612,N_1033,N_1073);
and U2613 (N_2613,N_1057,N_1645);
nor U2614 (N_2614,N_1261,N_1900);
nor U2615 (N_2615,N_1099,N_1536);
or U2616 (N_2616,N_1503,N_1928);
nand U2617 (N_2617,N_1055,N_1799);
or U2618 (N_2618,N_1061,N_1559);
nand U2619 (N_2619,N_1203,N_1529);
xnor U2620 (N_2620,N_1155,N_1999);
nor U2621 (N_2621,N_1721,N_1824);
or U2622 (N_2622,N_1520,N_1937);
nand U2623 (N_2623,N_1490,N_1165);
nand U2624 (N_2624,N_1750,N_1464);
and U2625 (N_2625,N_1345,N_1992);
or U2626 (N_2626,N_1197,N_1983);
xor U2627 (N_2627,N_1602,N_1117);
nor U2628 (N_2628,N_1100,N_1431);
and U2629 (N_2629,N_1565,N_1062);
nand U2630 (N_2630,N_1565,N_1600);
and U2631 (N_2631,N_1243,N_1658);
nand U2632 (N_2632,N_1911,N_1104);
or U2633 (N_2633,N_1776,N_1827);
nor U2634 (N_2634,N_1782,N_1748);
and U2635 (N_2635,N_1562,N_1539);
and U2636 (N_2636,N_1780,N_1711);
nand U2637 (N_2637,N_1409,N_1911);
or U2638 (N_2638,N_1598,N_1809);
or U2639 (N_2639,N_1683,N_1960);
and U2640 (N_2640,N_1859,N_1762);
nor U2641 (N_2641,N_1926,N_1309);
nor U2642 (N_2642,N_1028,N_1229);
or U2643 (N_2643,N_1579,N_1060);
or U2644 (N_2644,N_1678,N_1459);
nor U2645 (N_2645,N_1696,N_1018);
xor U2646 (N_2646,N_1740,N_1773);
and U2647 (N_2647,N_1232,N_1651);
nand U2648 (N_2648,N_1545,N_1314);
and U2649 (N_2649,N_1826,N_1571);
and U2650 (N_2650,N_1850,N_1223);
and U2651 (N_2651,N_1060,N_1805);
nand U2652 (N_2652,N_1909,N_1104);
nor U2653 (N_2653,N_1648,N_1820);
and U2654 (N_2654,N_1872,N_1857);
or U2655 (N_2655,N_1871,N_1216);
nand U2656 (N_2656,N_1432,N_1853);
xnor U2657 (N_2657,N_1058,N_1079);
xnor U2658 (N_2658,N_1176,N_1272);
or U2659 (N_2659,N_1542,N_1328);
or U2660 (N_2660,N_1465,N_1527);
or U2661 (N_2661,N_1455,N_1053);
nand U2662 (N_2662,N_1510,N_1058);
nor U2663 (N_2663,N_1542,N_1580);
and U2664 (N_2664,N_1426,N_1946);
nor U2665 (N_2665,N_1131,N_1097);
and U2666 (N_2666,N_1039,N_1431);
or U2667 (N_2667,N_1317,N_1439);
nand U2668 (N_2668,N_1296,N_1701);
and U2669 (N_2669,N_1446,N_1580);
nor U2670 (N_2670,N_1247,N_1285);
nand U2671 (N_2671,N_1774,N_1559);
and U2672 (N_2672,N_1264,N_1706);
nand U2673 (N_2673,N_1958,N_1817);
nand U2674 (N_2674,N_1588,N_1638);
or U2675 (N_2675,N_1758,N_1225);
and U2676 (N_2676,N_1654,N_1297);
xnor U2677 (N_2677,N_1581,N_1660);
or U2678 (N_2678,N_1703,N_1706);
or U2679 (N_2679,N_1418,N_1497);
and U2680 (N_2680,N_1680,N_1005);
nand U2681 (N_2681,N_1695,N_1920);
nand U2682 (N_2682,N_1585,N_1052);
nor U2683 (N_2683,N_1396,N_1978);
nand U2684 (N_2684,N_1713,N_1608);
or U2685 (N_2685,N_1228,N_1257);
or U2686 (N_2686,N_1511,N_1034);
xnor U2687 (N_2687,N_1786,N_1937);
nand U2688 (N_2688,N_1275,N_1216);
nand U2689 (N_2689,N_1753,N_1495);
xor U2690 (N_2690,N_1110,N_1727);
nor U2691 (N_2691,N_1254,N_1697);
nand U2692 (N_2692,N_1043,N_1639);
nand U2693 (N_2693,N_1480,N_1417);
or U2694 (N_2694,N_1811,N_1410);
xor U2695 (N_2695,N_1000,N_1238);
and U2696 (N_2696,N_1591,N_1398);
and U2697 (N_2697,N_1340,N_1850);
or U2698 (N_2698,N_1907,N_1738);
nand U2699 (N_2699,N_1278,N_1452);
nand U2700 (N_2700,N_1290,N_1433);
nor U2701 (N_2701,N_1893,N_1637);
and U2702 (N_2702,N_1766,N_1409);
nor U2703 (N_2703,N_1012,N_1264);
or U2704 (N_2704,N_1619,N_1466);
xor U2705 (N_2705,N_1483,N_1967);
xor U2706 (N_2706,N_1306,N_1923);
xor U2707 (N_2707,N_1492,N_1777);
nor U2708 (N_2708,N_1739,N_1160);
xor U2709 (N_2709,N_1577,N_1739);
nor U2710 (N_2710,N_1371,N_1585);
nor U2711 (N_2711,N_1580,N_1135);
nand U2712 (N_2712,N_1313,N_1242);
and U2713 (N_2713,N_1155,N_1641);
nand U2714 (N_2714,N_1980,N_1473);
xor U2715 (N_2715,N_1679,N_1150);
nor U2716 (N_2716,N_1522,N_1675);
and U2717 (N_2717,N_1509,N_1264);
xor U2718 (N_2718,N_1216,N_1075);
or U2719 (N_2719,N_1841,N_1023);
or U2720 (N_2720,N_1662,N_1794);
xnor U2721 (N_2721,N_1538,N_1046);
or U2722 (N_2722,N_1036,N_1399);
xnor U2723 (N_2723,N_1481,N_1497);
nor U2724 (N_2724,N_1502,N_1934);
nand U2725 (N_2725,N_1655,N_1893);
nor U2726 (N_2726,N_1240,N_1249);
nand U2727 (N_2727,N_1876,N_1143);
xor U2728 (N_2728,N_1545,N_1972);
nor U2729 (N_2729,N_1270,N_1849);
xnor U2730 (N_2730,N_1828,N_1096);
nor U2731 (N_2731,N_1810,N_1293);
nor U2732 (N_2732,N_1451,N_1984);
nor U2733 (N_2733,N_1415,N_1168);
nand U2734 (N_2734,N_1353,N_1244);
or U2735 (N_2735,N_1914,N_1905);
nand U2736 (N_2736,N_1849,N_1480);
xnor U2737 (N_2737,N_1225,N_1390);
and U2738 (N_2738,N_1676,N_1630);
and U2739 (N_2739,N_1017,N_1454);
and U2740 (N_2740,N_1798,N_1828);
or U2741 (N_2741,N_1860,N_1654);
nor U2742 (N_2742,N_1586,N_1646);
nand U2743 (N_2743,N_1967,N_1598);
and U2744 (N_2744,N_1135,N_1529);
nor U2745 (N_2745,N_1811,N_1698);
or U2746 (N_2746,N_1475,N_1882);
or U2747 (N_2747,N_1275,N_1149);
nand U2748 (N_2748,N_1374,N_1615);
or U2749 (N_2749,N_1518,N_1695);
nor U2750 (N_2750,N_1128,N_1511);
nor U2751 (N_2751,N_1697,N_1099);
and U2752 (N_2752,N_1456,N_1253);
xnor U2753 (N_2753,N_1725,N_1713);
xnor U2754 (N_2754,N_1779,N_1787);
nand U2755 (N_2755,N_1142,N_1954);
or U2756 (N_2756,N_1335,N_1470);
or U2757 (N_2757,N_1290,N_1649);
xnor U2758 (N_2758,N_1052,N_1809);
xor U2759 (N_2759,N_1753,N_1571);
nand U2760 (N_2760,N_1055,N_1328);
nor U2761 (N_2761,N_1941,N_1532);
and U2762 (N_2762,N_1238,N_1408);
or U2763 (N_2763,N_1355,N_1176);
nor U2764 (N_2764,N_1917,N_1009);
xor U2765 (N_2765,N_1360,N_1506);
nor U2766 (N_2766,N_1407,N_1933);
xnor U2767 (N_2767,N_1708,N_1860);
and U2768 (N_2768,N_1844,N_1455);
nor U2769 (N_2769,N_1770,N_1593);
nor U2770 (N_2770,N_1779,N_1889);
xnor U2771 (N_2771,N_1062,N_1925);
xnor U2772 (N_2772,N_1081,N_1528);
nor U2773 (N_2773,N_1982,N_1214);
nor U2774 (N_2774,N_1429,N_1084);
xnor U2775 (N_2775,N_1274,N_1252);
and U2776 (N_2776,N_1922,N_1196);
nor U2777 (N_2777,N_1556,N_1006);
or U2778 (N_2778,N_1813,N_1793);
and U2779 (N_2779,N_1332,N_1625);
nand U2780 (N_2780,N_1421,N_1616);
nand U2781 (N_2781,N_1335,N_1025);
nand U2782 (N_2782,N_1526,N_1251);
nor U2783 (N_2783,N_1281,N_1374);
xnor U2784 (N_2784,N_1731,N_1301);
or U2785 (N_2785,N_1990,N_1910);
or U2786 (N_2786,N_1812,N_1608);
nor U2787 (N_2787,N_1177,N_1493);
and U2788 (N_2788,N_1708,N_1058);
and U2789 (N_2789,N_1027,N_1279);
and U2790 (N_2790,N_1116,N_1932);
xnor U2791 (N_2791,N_1503,N_1554);
nor U2792 (N_2792,N_1245,N_1869);
and U2793 (N_2793,N_1742,N_1430);
xnor U2794 (N_2794,N_1050,N_1159);
nor U2795 (N_2795,N_1736,N_1567);
nor U2796 (N_2796,N_1549,N_1939);
nor U2797 (N_2797,N_1870,N_1003);
and U2798 (N_2798,N_1906,N_1394);
nor U2799 (N_2799,N_1604,N_1865);
or U2800 (N_2800,N_1266,N_1766);
xnor U2801 (N_2801,N_1179,N_1186);
nand U2802 (N_2802,N_1175,N_1243);
xor U2803 (N_2803,N_1868,N_1802);
or U2804 (N_2804,N_1074,N_1860);
or U2805 (N_2805,N_1254,N_1282);
nor U2806 (N_2806,N_1885,N_1048);
and U2807 (N_2807,N_1355,N_1527);
and U2808 (N_2808,N_1734,N_1066);
nor U2809 (N_2809,N_1571,N_1403);
and U2810 (N_2810,N_1808,N_1309);
nand U2811 (N_2811,N_1125,N_1702);
and U2812 (N_2812,N_1404,N_1992);
nor U2813 (N_2813,N_1425,N_1785);
xor U2814 (N_2814,N_1135,N_1525);
nor U2815 (N_2815,N_1686,N_1400);
xor U2816 (N_2816,N_1495,N_1229);
or U2817 (N_2817,N_1530,N_1923);
nor U2818 (N_2818,N_1122,N_1404);
xnor U2819 (N_2819,N_1943,N_1850);
nand U2820 (N_2820,N_1962,N_1308);
xor U2821 (N_2821,N_1108,N_1048);
nor U2822 (N_2822,N_1454,N_1874);
nor U2823 (N_2823,N_1577,N_1565);
and U2824 (N_2824,N_1507,N_1487);
nor U2825 (N_2825,N_1968,N_1379);
xor U2826 (N_2826,N_1962,N_1842);
or U2827 (N_2827,N_1585,N_1909);
and U2828 (N_2828,N_1791,N_1552);
or U2829 (N_2829,N_1775,N_1053);
nand U2830 (N_2830,N_1529,N_1091);
xor U2831 (N_2831,N_1897,N_1269);
xnor U2832 (N_2832,N_1171,N_1633);
nand U2833 (N_2833,N_1567,N_1116);
nand U2834 (N_2834,N_1771,N_1612);
or U2835 (N_2835,N_1268,N_1760);
xnor U2836 (N_2836,N_1371,N_1807);
or U2837 (N_2837,N_1282,N_1134);
and U2838 (N_2838,N_1396,N_1529);
nand U2839 (N_2839,N_1972,N_1722);
and U2840 (N_2840,N_1441,N_1636);
or U2841 (N_2841,N_1126,N_1640);
xnor U2842 (N_2842,N_1181,N_1333);
nand U2843 (N_2843,N_1810,N_1722);
nor U2844 (N_2844,N_1933,N_1174);
and U2845 (N_2845,N_1852,N_1537);
or U2846 (N_2846,N_1009,N_1352);
xor U2847 (N_2847,N_1175,N_1860);
or U2848 (N_2848,N_1833,N_1562);
and U2849 (N_2849,N_1037,N_1268);
xnor U2850 (N_2850,N_1834,N_1971);
nand U2851 (N_2851,N_1300,N_1325);
and U2852 (N_2852,N_1213,N_1523);
xnor U2853 (N_2853,N_1410,N_1632);
nand U2854 (N_2854,N_1968,N_1427);
nand U2855 (N_2855,N_1433,N_1449);
and U2856 (N_2856,N_1768,N_1598);
xor U2857 (N_2857,N_1315,N_1936);
and U2858 (N_2858,N_1215,N_1019);
nand U2859 (N_2859,N_1065,N_1488);
nor U2860 (N_2860,N_1099,N_1416);
xnor U2861 (N_2861,N_1135,N_1402);
and U2862 (N_2862,N_1504,N_1898);
xor U2863 (N_2863,N_1742,N_1311);
and U2864 (N_2864,N_1362,N_1799);
nand U2865 (N_2865,N_1613,N_1393);
nor U2866 (N_2866,N_1549,N_1902);
or U2867 (N_2867,N_1005,N_1491);
or U2868 (N_2868,N_1049,N_1753);
and U2869 (N_2869,N_1884,N_1678);
xor U2870 (N_2870,N_1778,N_1305);
and U2871 (N_2871,N_1140,N_1700);
nand U2872 (N_2872,N_1551,N_1468);
and U2873 (N_2873,N_1987,N_1490);
nand U2874 (N_2874,N_1725,N_1002);
xor U2875 (N_2875,N_1345,N_1685);
xor U2876 (N_2876,N_1104,N_1253);
and U2877 (N_2877,N_1422,N_1521);
nand U2878 (N_2878,N_1246,N_1670);
xor U2879 (N_2879,N_1674,N_1166);
or U2880 (N_2880,N_1201,N_1262);
and U2881 (N_2881,N_1673,N_1863);
or U2882 (N_2882,N_1417,N_1308);
and U2883 (N_2883,N_1355,N_1434);
xnor U2884 (N_2884,N_1641,N_1436);
nor U2885 (N_2885,N_1940,N_1687);
nor U2886 (N_2886,N_1734,N_1730);
nor U2887 (N_2887,N_1964,N_1135);
xnor U2888 (N_2888,N_1569,N_1374);
or U2889 (N_2889,N_1984,N_1734);
nor U2890 (N_2890,N_1901,N_1893);
nor U2891 (N_2891,N_1695,N_1373);
or U2892 (N_2892,N_1775,N_1103);
nand U2893 (N_2893,N_1909,N_1869);
and U2894 (N_2894,N_1371,N_1206);
nand U2895 (N_2895,N_1999,N_1791);
and U2896 (N_2896,N_1697,N_1354);
nand U2897 (N_2897,N_1297,N_1827);
or U2898 (N_2898,N_1191,N_1023);
nand U2899 (N_2899,N_1396,N_1658);
nor U2900 (N_2900,N_1741,N_1416);
nand U2901 (N_2901,N_1790,N_1991);
xnor U2902 (N_2902,N_1145,N_1384);
and U2903 (N_2903,N_1411,N_1333);
nand U2904 (N_2904,N_1435,N_1823);
xor U2905 (N_2905,N_1364,N_1313);
nand U2906 (N_2906,N_1221,N_1565);
xor U2907 (N_2907,N_1084,N_1372);
xnor U2908 (N_2908,N_1870,N_1367);
or U2909 (N_2909,N_1370,N_1329);
nand U2910 (N_2910,N_1907,N_1748);
nand U2911 (N_2911,N_1225,N_1675);
nand U2912 (N_2912,N_1480,N_1199);
nand U2913 (N_2913,N_1111,N_1335);
nand U2914 (N_2914,N_1914,N_1040);
xor U2915 (N_2915,N_1222,N_1810);
xnor U2916 (N_2916,N_1888,N_1289);
and U2917 (N_2917,N_1832,N_1062);
xnor U2918 (N_2918,N_1261,N_1313);
nor U2919 (N_2919,N_1074,N_1762);
nor U2920 (N_2920,N_1232,N_1202);
nand U2921 (N_2921,N_1629,N_1497);
nor U2922 (N_2922,N_1274,N_1625);
and U2923 (N_2923,N_1209,N_1514);
nand U2924 (N_2924,N_1110,N_1076);
nand U2925 (N_2925,N_1325,N_1748);
nand U2926 (N_2926,N_1448,N_1962);
nor U2927 (N_2927,N_1470,N_1611);
nand U2928 (N_2928,N_1648,N_1762);
or U2929 (N_2929,N_1065,N_1158);
nor U2930 (N_2930,N_1361,N_1272);
nand U2931 (N_2931,N_1262,N_1250);
and U2932 (N_2932,N_1066,N_1978);
xor U2933 (N_2933,N_1313,N_1349);
or U2934 (N_2934,N_1161,N_1279);
or U2935 (N_2935,N_1919,N_1126);
nor U2936 (N_2936,N_1838,N_1737);
nand U2937 (N_2937,N_1964,N_1794);
nand U2938 (N_2938,N_1598,N_1363);
nor U2939 (N_2939,N_1641,N_1710);
xor U2940 (N_2940,N_1633,N_1340);
and U2941 (N_2941,N_1291,N_1693);
nor U2942 (N_2942,N_1956,N_1655);
xor U2943 (N_2943,N_1999,N_1651);
xor U2944 (N_2944,N_1681,N_1866);
xor U2945 (N_2945,N_1988,N_1087);
or U2946 (N_2946,N_1290,N_1898);
or U2947 (N_2947,N_1887,N_1468);
and U2948 (N_2948,N_1921,N_1161);
xor U2949 (N_2949,N_1791,N_1345);
xnor U2950 (N_2950,N_1484,N_1116);
or U2951 (N_2951,N_1539,N_1649);
xor U2952 (N_2952,N_1594,N_1451);
or U2953 (N_2953,N_1626,N_1800);
and U2954 (N_2954,N_1642,N_1530);
nor U2955 (N_2955,N_1869,N_1521);
nand U2956 (N_2956,N_1120,N_1888);
and U2957 (N_2957,N_1174,N_1131);
nand U2958 (N_2958,N_1073,N_1025);
and U2959 (N_2959,N_1943,N_1186);
xor U2960 (N_2960,N_1584,N_1666);
and U2961 (N_2961,N_1607,N_1848);
nor U2962 (N_2962,N_1171,N_1809);
xnor U2963 (N_2963,N_1509,N_1446);
xnor U2964 (N_2964,N_1279,N_1699);
nor U2965 (N_2965,N_1241,N_1460);
or U2966 (N_2966,N_1779,N_1864);
nand U2967 (N_2967,N_1836,N_1703);
nor U2968 (N_2968,N_1659,N_1621);
and U2969 (N_2969,N_1306,N_1370);
or U2970 (N_2970,N_1724,N_1118);
or U2971 (N_2971,N_1298,N_1619);
nand U2972 (N_2972,N_1248,N_1974);
xnor U2973 (N_2973,N_1798,N_1229);
nor U2974 (N_2974,N_1321,N_1822);
nand U2975 (N_2975,N_1931,N_1280);
and U2976 (N_2976,N_1796,N_1646);
or U2977 (N_2977,N_1422,N_1315);
and U2978 (N_2978,N_1693,N_1749);
nand U2979 (N_2979,N_1602,N_1298);
nand U2980 (N_2980,N_1912,N_1964);
xnor U2981 (N_2981,N_1706,N_1743);
or U2982 (N_2982,N_1422,N_1468);
and U2983 (N_2983,N_1152,N_1301);
or U2984 (N_2984,N_1384,N_1634);
xnor U2985 (N_2985,N_1010,N_1347);
or U2986 (N_2986,N_1253,N_1243);
nor U2987 (N_2987,N_1874,N_1580);
xor U2988 (N_2988,N_1582,N_1262);
and U2989 (N_2989,N_1722,N_1279);
and U2990 (N_2990,N_1013,N_1358);
or U2991 (N_2991,N_1280,N_1877);
xnor U2992 (N_2992,N_1407,N_1441);
xnor U2993 (N_2993,N_1849,N_1185);
or U2994 (N_2994,N_1651,N_1941);
and U2995 (N_2995,N_1789,N_1607);
xor U2996 (N_2996,N_1385,N_1668);
and U2997 (N_2997,N_1435,N_1314);
and U2998 (N_2998,N_1130,N_1922);
nor U2999 (N_2999,N_1051,N_1299);
xnor UO_0 (O_0,N_2292,N_2039);
or UO_1 (O_1,N_2330,N_2360);
nand UO_2 (O_2,N_2644,N_2365);
nor UO_3 (O_3,N_2731,N_2976);
nand UO_4 (O_4,N_2498,N_2073);
nand UO_5 (O_5,N_2478,N_2736);
or UO_6 (O_6,N_2439,N_2595);
nand UO_7 (O_7,N_2719,N_2729);
and UO_8 (O_8,N_2616,N_2371);
nor UO_9 (O_9,N_2100,N_2465);
nor UO_10 (O_10,N_2176,N_2187);
xnor UO_11 (O_11,N_2219,N_2528);
or UO_12 (O_12,N_2566,N_2254);
or UO_13 (O_13,N_2312,N_2996);
or UO_14 (O_14,N_2916,N_2377);
xor UO_15 (O_15,N_2770,N_2687);
nor UO_16 (O_16,N_2127,N_2799);
nor UO_17 (O_17,N_2400,N_2994);
nand UO_18 (O_18,N_2024,N_2751);
xor UO_19 (O_19,N_2581,N_2180);
nand UO_20 (O_20,N_2295,N_2072);
xor UO_21 (O_21,N_2332,N_2970);
xnor UO_22 (O_22,N_2317,N_2630);
and UO_23 (O_23,N_2211,N_2392);
and UO_24 (O_24,N_2434,N_2138);
and UO_25 (O_25,N_2645,N_2756);
or UO_26 (O_26,N_2730,N_2798);
nand UO_27 (O_27,N_2413,N_2261);
and UO_28 (O_28,N_2135,N_2833);
or UO_29 (O_29,N_2071,N_2085);
nor UO_30 (O_30,N_2386,N_2558);
or UO_31 (O_31,N_2381,N_2605);
xor UO_32 (O_32,N_2245,N_2412);
nand UO_33 (O_33,N_2411,N_2054);
or UO_34 (O_34,N_2390,N_2097);
nor UO_35 (O_35,N_2568,N_2503);
and UO_36 (O_36,N_2524,N_2713);
xnor UO_37 (O_37,N_2949,N_2957);
nor UO_38 (O_38,N_2603,N_2422);
nor UO_39 (O_39,N_2734,N_2712);
nand UO_40 (O_40,N_2746,N_2325);
nor UO_41 (O_41,N_2574,N_2410);
or UO_42 (O_42,N_2011,N_2841);
xor UO_43 (O_43,N_2843,N_2140);
nand UO_44 (O_44,N_2518,N_2896);
and UO_45 (O_45,N_2920,N_2940);
or UO_46 (O_46,N_2326,N_2336);
or UO_47 (O_47,N_2702,N_2075);
nand UO_48 (O_48,N_2469,N_2271);
and UO_49 (O_49,N_2293,N_2108);
or UO_50 (O_50,N_2851,N_2419);
nor UO_51 (O_51,N_2895,N_2682);
and UO_52 (O_52,N_2701,N_2221);
xnor UO_53 (O_53,N_2043,N_2821);
xnor UO_54 (O_54,N_2253,N_2119);
nor UO_55 (O_55,N_2366,N_2619);
xnor UO_56 (O_56,N_2372,N_2923);
or UO_57 (O_57,N_2264,N_2796);
xnor UO_58 (O_58,N_2456,N_2881);
and UO_59 (O_59,N_2868,N_2786);
xor UO_60 (O_60,N_2234,N_2888);
xor UO_61 (O_61,N_2549,N_2569);
nor UO_62 (O_62,N_2250,N_2463);
and UO_63 (O_63,N_2811,N_2276);
or UO_64 (O_64,N_2307,N_2107);
and UO_65 (O_65,N_2753,N_2808);
nand UO_66 (O_66,N_2583,N_2178);
xor UO_67 (O_67,N_2198,N_2132);
nor UO_68 (O_68,N_2783,N_2305);
and UO_69 (O_69,N_2597,N_2398);
and UO_70 (O_70,N_2093,N_2184);
xor UO_71 (O_71,N_2692,N_2338);
xor UO_72 (O_72,N_2709,N_2785);
nor UO_73 (O_73,N_2829,N_2532);
and UO_74 (O_74,N_2046,N_2792);
xnor UO_75 (O_75,N_2448,N_2860);
or UO_76 (O_76,N_2420,N_2815);
nand UO_77 (O_77,N_2711,N_2450);
nor UO_78 (O_78,N_2113,N_2077);
and UO_79 (O_79,N_2871,N_2846);
xor UO_80 (O_80,N_2329,N_2502);
and UO_81 (O_81,N_2737,N_2334);
xor UO_82 (O_82,N_2002,N_2214);
and UO_83 (O_83,N_2742,N_2070);
nand UO_84 (O_84,N_2267,N_2089);
nand UO_85 (O_85,N_2678,N_2651);
and UO_86 (O_86,N_2006,N_2385);
and UO_87 (O_87,N_2580,N_2637);
or UO_88 (O_88,N_2534,N_2354);
and UO_89 (O_89,N_2015,N_2417);
nand UO_90 (O_90,N_2589,N_2794);
nor UO_91 (O_91,N_2356,N_2927);
or UO_92 (O_92,N_2509,N_2231);
and UO_93 (O_93,N_2810,N_2800);
or UO_94 (O_94,N_2766,N_2299);
nor UO_95 (O_95,N_2368,N_2752);
nor UO_96 (O_96,N_2975,N_2690);
or UO_97 (O_97,N_2035,N_2009);
and UO_98 (O_98,N_2714,N_2150);
and UO_99 (O_99,N_2435,N_2579);
nand UO_100 (O_100,N_2879,N_2215);
and UO_101 (O_101,N_2470,N_2216);
nor UO_102 (O_102,N_2206,N_2159);
xor UO_103 (O_103,N_2521,N_2062);
or UO_104 (O_104,N_2930,N_2672);
xnor UO_105 (O_105,N_2546,N_2931);
and UO_106 (O_106,N_2019,N_2902);
and UO_107 (O_107,N_2486,N_2715);
nand UO_108 (O_108,N_2225,N_2196);
nand UO_109 (O_109,N_2956,N_2983);
xor UO_110 (O_110,N_2080,N_2220);
nor UO_111 (O_111,N_2488,N_2194);
nor UO_112 (O_112,N_2535,N_2727);
nand UO_113 (O_113,N_2660,N_2563);
and UO_114 (O_114,N_2144,N_2166);
or UO_115 (O_115,N_2269,N_2228);
nor UO_116 (O_116,N_2707,N_2958);
nand UO_117 (O_117,N_2614,N_2606);
nor UO_118 (O_118,N_2747,N_2001);
nor UO_119 (O_119,N_2161,N_2852);
nand UO_120 (O_120,N_2748,N_2476);
nor UO_121 (O_121,N_2491,N_2874);
and UO_122 (O_122,N_2865,N_2936);
nand UO_123 (O_123,N_2255,N_2241);
or UO_124 (O_124,N_2716,N_2732);
and UO_125 (O_125,N_2133,N_2530);
and UO_126 (O_126,N_2803,N_2617);
and UO_127 (O_127,N_2912,N_2723);
nor UO_128 (O_128,N_2205,N_2838);
and UO_129 (O_129,N_2437,N_2671);
nor UO_130 (O_130,N_2939,N_2472);
or UO_131 (O_131,N_2370,N_2082);
xnor UO_132 (O_132,N_2531,N_2102);
xnor UO_133 (O_133,N_2683,N_2240);
xor UO_134 (O_134,N_2397,N_2827);
or UO_135 (O_135,N_2944,N_2513);
nor UO_136 (O_136,N_2979,N_2117);
xor UO_137 (O_137,N_2899,N_2275);
nand UO_138 (O_138,N_2512,N_2555);
nand UO_139 (O_139,N_2157,N_2327);
nand UO_140 (O_140,N_2084,N_2428);
xnor UO_141 (O_141,N_2608,N_2935);
nor UO_142 (O_142,N_2167,N_2806);
nor UO_143 (O_143,N_2493,N_2812);
nand UO_144 (O_144,N_2506,N_2725);
or UO_145 (O_145,N_2848,N_2952);
nand UO_146 (O_146,N_2677,N_2265);
and UO_147 (O_147,N_2367,N_2318);
or UO_148 (O_148,N_2646,N_2622);
and UO_149 (O_149,N_2067,N_2757);
xor UO_150 (O_150,N_2954,N_2867);
or UO_151 (O_151,N_2131,N_2499);
xor UO_152 (O_152,N_2027,N_2304);
nor UO_153 (O_153,N_2567,N_2768);
nor UO_154 (O_154,N_2056,N_2373);
or UO_155 (O_155,N_2125,N_2331);
nor UO_156 (O_156,N_2691,N_2320);
nand UO_157 (O_157,N_2416,N_2995);
nand UO_158 (O_158,N_2090,N_2349);
and UO_159 (O_159,N_2919,N_2076);
nand UO_160 (O_160,N_2459,N_2230);
nand UO_161 (O_161,N_2012,N_2765);
nor UO_162 (O_162,N_2190,N_2802);
nand UO_163 (O_163,N_2328,N_2489);
nor UO_164 (O_164,N_2175,N_2044);
nand UO_165 (O_165,N_2351,N_2246);
nor UO_166 (O_166,N_2591,N_2309);
and UO_167 (O_167,N_2733,N_2183);
nor UO_168 (O_168,N_2624,N_2778);
or UO_169 (O_169,N_2032,N_2648);
and UO_170 (O_170,N_2817,N_2037);
xnor UO_171 (O_171,N_2130,N_2383);
xor UO_172 (O_172,N_2620,N_2844);
and UO_173 (O_173,N_2586,N_2659);
nand UO_174 (O_174,N_2041,N_2876);
xor UO_175 (O_175,N_2281,N_2855);
or UO_176 (O_176,N_2301,N_2950);
nand UO_177 (O_177,N_2629,N_2985);
xor UO_178 (O_178,N_2654,N_2163);
nand UO_179 (O_179,N_2441,N_2197);
nand UO_180 (O_180,N_2744,N_2200);
nand UO_181 (O_181,N_2721,N_2378);
and UO_182 (O_182,N_2953,N_2929);
or UO_183 (O_183,N_2455,N_2164);
nor UO_184 (O_184,N_2092,N_2143);
nor UO_185 (O_185,N_2227,N_2947);
or UO_186 (O_186,N_2505,N_2182);
or UO_187 (O_187,N_2830,N_2280);
or UO_188 (O_188,N_2273,N_2462);
xor UO_189 (O_189,N_2050,N_2741);
nor UO_190 (O_190,N_2551,N_2086);
and UO_191 (O_191,N_2514,N_2475);
or UO_192 (O_192,N_2051,N_2653);
xnor UO_193 (O_193,N_2965,N_2487);
nand UO_194 (O_194,N_2823,N_2618);
nor UO_195 (O_195,N_2461,N_2835);
or UO_196 (O_196,N_2507,N_2961);
or UO_197 (O_197,N_2064,N_2836);
xnor UO_198 (O_198,N_2394,N_2519);
nand UO_199 (O_199,N_2495,N_2527);
and UO_200 (O_200,N_2421,N_2887);
and UO_201 (O_201,N_2118,N_2155);
and UO_202 (O_202,N_2625,N_2872);
xor UO_203 (O_203,N_2376,N_2943);
or UO_204 (O_204,N_2447,N_2602);
and UO_205 (O_205,N_2763,N_2652);
or UO_206 (O_206,N_2847,N_2233);
xor UO_207 (O_207,N_2700,N_2477);
or UO_208 (O_208,N_2485,N_2708);
and UO_209 (O_209,N_2705,N_2226);
nor UO_210 (O_210,N_2500,N_2818);
or UO_211 (O_211,N_2516,N_2316);
and UO_212 (O_212,N_2526,N_2703);
or UO_213 (O_213,N_2596,N_2666);
and UO_214 (O_214,N_2793,N_2758);
xor UO_215 (O_215,N_2669,N_2286);
nor UO_216 (O_216,N_2880,N_2402);
xor UO_217 (O_217,N_2856,N_2193);
nand UO_218 (O_218,N_2169,N_2081);
nand UO_219 (O_219,N_2340,N_2826);
or UO_220 (O_220,N_2529,N_2662);
nor UO_221 (O_221,N_2875,N_2955);
nand UO_222 (O_222,N_2387,N_2128);
nor UO_223 (O_223,N_2680,N_2932);
or UO_224 (O_224,N_2698,N_2988);
nor UO_225 (O_225,N_2021,N_2302);
and UO_226 (O_226,N_2631,N_2091);
and UO_227 (O_227,N_2882,N_2460);
nand UO_228 (O_228,N_2972,N_2425);
and UO_229 (O_229,N_2112,N_2480);
xor UO_230 (O_230,N_2772,N_2423);
nor UO_231 (O_231,N_2650,N_2904);
nor UO_232 (O_232,N_2969,N_2415);
nor UO_233 (O_233,N_2426,N_2688);
xor UO_234 (O_234,N_2160,N_2542);
nand UO_235 (O_235,N_2098,N_2718);
or UO_236 (O_236,N_2490,N_2473);
nand UO_237 (O_237,N_2152,N_2199);
nor UO_238 (O_238,N_2883,N_2642);
nand UO_239 (O_239,N_2989,N_2224);
nand UO_240 (O_240,N_2186,N_2681);
or UO_241 (O_241,N_2822,N_2928);
xnor UO_242 (O_242,N_2481,N_2268);
and UO_243 (O_243,N_2791,N_2539);
or UO_244 (O_244,N_2023,N_2834);
nor UO_245 (O_245,N_2839,N_2594);
or UO_246 (O_246,N_2104,N_2446);
xnor UO_247 (O_247,N_2548,N_2162);
nor UO_248 (O_248,N_2258,N_2750);
nand UO_249 (O_249,N_2743,N_2000);
xnor UO_250 (O_250,N_2877,N_2977);
and UO_251 (O_251,N_2592,N_2869);
and UO_252 (O_252,N_2863,N_2572);
nor UO_253 (O_253,N_2915,N_2571);
nor UO_254 (O_254,N_2418,N_2389);
or UO_255 (O_255,N_2556,N_2828);
or UO_256 (O_256,N_2430,N_2083);
nor UO_257 (O_257,N_2760,N_2171);
nand UO_258 (O_258,N_2065,N_2116);
or UO_259 (O_259,N_2388,N_2686);
or UO_260 (O_260,N_2892,N_2464);
nand UO_261 (O_261,N_2345,N_2355);
nand UO_262 (O_262,N_2893,N_2278);
and UO_263 (O_263,N_2195,N_2306);
nor UO_264 (O_264,N_2382,N_2926);
and UO_265 (O_265,N_2636,N_2026);
xnor UO_266 (O_266,N_2344,N_2759);
nor UO_267 (O_267,N_2008,N_2873);
nand UO_268 (O_268,N_2795,N_2343);
nor UO_269 (O_269,N_2003,N_2192);
xnor UO_270 (O_270,N_2361,N_2966);
nand UO_271 (O_271,N_2561,N_2754);
nand UO_272 (O_272,N_2545,N_2445);
and UO_273 (O_273,N_2639,N_2626);
nor UO_274 (O_274,N_2628,N_2523);
or UO_275 (O_275,N_2153,N_2609);
and UO_276 (O_276,N_2761,N_2287);
xnor UO_277 (O_277,N_2238,N_2212);
xnor UO_278 (O_278,N_2266,N_2739);
or UO_279 (O_279,N_2993,N_2474);
xnor UO_280 (O_280,N_2951,N_2886);
or UO_281 (O_281,N_2964,N_2982);
or UO_282 (O_282,N_2864,N_2122);
or UO_283 (O_283,N_2096,N_2170);
nor UO_284 (O_284,N_2058,N_2909);
nand UO_285 (O_285,N_2068,N_2668);
and UO_286 (O_286,N_2676,N_2501);
nand UO_287 (O_287,N_2962,N_2693);
or UO_288 (O_288,N_2780,N_2429);
or UO_289 (O_289,N_2570,N_2109);
nor UO_290 (O_290,N_2126,N_2517);
nand UO_291 (O_291,N_2764,N_2154);
xor UO_292 (O_292,N_2028,N_2087);
nand UO_293 (O_293,N_2726,N_2053);
nand UO_294 (O_294,N_2177,N_2057);
xor UO_295 (O_295,N_2897,N_2059);
or UO_296 (O_296,N_2640,N_2560);
and UO_297 (O_297,N_2249,N_2277);
nor UO_298 (O_298,N_2735,N_2358);
nand UO_299 (O_299,N_2638,N_2635);
nor UO_300 (O_300,N_2740,N_2079);
nand UO_301 (O_301,N_2576,N_2244);
nand UO_302 (O_302,N_2937,N_2997);
nor UO_303 (O_303,N_2536,N_2562);
xor UO_304 (O_304,N_2854,N_2862);
xor UO_305 (O_305,N_2906,N_2728);
or UO_306 (O_306,N_2088,N_2657);
nor UO_307 (O_307,N_2438,N_2840);
or UO_308 (O_308,N_2934,N_2820);
nor UO_309 (O_309,N_2363,N_2968);
or UO_310 (O_310,N_2272,N_2380);
and UO_311 (O_311,N_2203,N_2313);
and UO_312 (O_312,N_2384,N_2337);
and UO_313 (O_313,N_2031,N_2859);
nand UO_314 (O_314,N_2910,N_2452);
and UO_315 (O_315,N_2717,N_2663);
or UO_316 (O_316,N_2350,N_2296);
and UO_317 (O_317,N_2670,N_2788);
xnor UO_318 (O_318,N_2223,N_2471);
and UO_319 (O_319,N_2781,N_2120);
or UO_320 (O_320,N_2809,N_2504);
and UO_321 (O_321,N_2992,N_2005);
or UO_322 (O_322,N_2999,N_2252);
nand UO_323 (O_323,N_2905,N_2814);
nor UO_324 (O_324,N_2158,N_2137);
or UO_325 (O_325,N_2172,N_2577);
or UO_326 (O_326,N_2837,N_2925);
and UO_327 (O_327,N_2453,N_2364);
or UO_328 (O_328,N_2938,N_2235);
or UO_329 (O_329,N_2458,N_2149);
nand UO_330 (O_330,N_2339,N_2615);
nor UO_331 (O_331,N_2511,N_2298);
or UO_332 (O_332,N_2342,N_2825);
and UO_333 (O_333,N_2346,N_2424);
and UO_334 (O_334,N_2482,N_2396);
nor UO_335 (O_335,N_2229,N_2291);
nand UO_336 (O_336,N_2946,N_2971);
nor UO_337 (O_337,N_2103,N_2559);
nand UO_338 (O_338,N_2007,N_2391);
xor UO_339 (O_339,N_2393,N_2805);
and UO_340 (O_340,N_2239,N_2496);
and UO_341 (O_341,N_2553,N_2061);
nor UO_342 (O_342,N_2789,N_2494);
xor UO_343 (O_343,N_2399,N_2724);
xor UO_344 (O_344,N_2352,N_2941);
or UO_345 (O_345,N_2134,N_2807);
nand UO_346 (O_346,N_2599,N_2924);
or UO_347 (O_347,N_2774,N_2901);
or UO_348 (O_348,N_2018,N_2404);
nand UO_349 (O_349,N_2684,N_2816);
nor UO_350 (O_350,N_2259,N_2767);
xnor UO_351 (O_351,N_2270,N_2801);
nor UO_352 (O_352,N_2210,N_2319);
and UO_353 (O_353,N_2374,N_2933);
nor UO_354 (O_354,N_2236,N_2921);
nand UO_355 (O_355,N_2903,N_2036);
or UO_356 (O_356,N_2124,N_2066);
xnor UO_357 (O_357,N_2607,N_2362);
xor UO_358 (O_358,N_2121,N_2649);
xor UO_359 (O_359,N_2322,N_2738);
and UO_360 (O_360,N_2565,N_2123);
nand UO_361 (O_361,N_2858,N_2308);
xor UO_362 (O_362,N_2771,N_2247);
nor UO_363 (O_363,N_2468,N_2537);
and UO_364 (O_364,N_2348,N_2525);
nor UO_365 (O_365,N_2853,N_2538);
or UO_366 (O_366,N_2694,N_2889);
or UO_367 (O_367,N_2288,N_2341);
and UO_368 (O_368,N_2866,N_2611);
nor UO_369 (O_369,N_2911,N_2168);
or UO_370 (O_370,N_2279,N_2689);
or UO_371 (O_371,N_2401,N_2959);
or UO_372 (O_372,N_2101,N_2706);
or UO_373 (O_373,N_2824,N_2990);
or UO_374 (O_374,N_2664,N_2633);
xnor UO_375 (O_375,N_2942,N_2790);
xnor UO_376 (O_376,N_2948,N_2894);
xor UO_377 (O_377,N_2074,N_2251);
nor UO_378 (O_378,N_2395,N_2333);
xor UO_379 (O_379,N_2454,N_2623);
nand UO_380 (O_380,N_2675,N_2359);
or UO_381 (O_381,N_2034,N_2641);
and UO_382 (O_382,N_2347,N_2467);
or UO_383 (O_383,N_2573,N_2773);
nor UO_384 (O_384,N_2020,N_2787);
or UO_385 (O_385,N_2141,N_2353);
nand UO_386 (O_386,N_2845,N_2991);
nor UO_387 (O_387,N_2048,N_2217);
nor UO_388 (O_388,N_2522,N_2405);
xor UO_389 (O_389,N_2627,N_2777);
or UO_390 (O_390,N_2408,N_2369);
nand UO_391 (O_391,N_2403,N_2179);
and UO_392 (O_392,N_2543,N_2049);
and UO_393 (O_393,N_2045,N_2656);
or UO_394 (O_394,N_2819,N_2311);
and UO_395 (O_395,N_2016,N_2173);
nor UO_396 (O_396,N_2960,N_2310);
or UO_397 (O_397,N_2181,N_2237);
or UO_398 (O_398,N_2095,N_2443);
or UO_399 (O_399,N_2878,N_2584);
or UO_400 (O_400,N_2967,N_2202);
nor UO_401 (O_401,N_2025,N_2661);
and UO_402 (O_402,N_2604,N_2047);
xor UO_403 (O_403,N_2797,N_2375);
xor UO_404 (O_404,N_2078,N_2665);
and UO_405 (O_405,N_2831,N_2520);
xnor UO_406 (O_406,N_2842,N_2963);
nand UO_407 (O_407,N_2945,N_2588);
xor UO_408 (O_408,N_2598,N_2643);
nand UO_409 (O_409,N_2634,N_2578);
or UO_410 (O_410,N_2442,N_2263);
nor UO_411 (O_411,N_2357,N_2321);
nand UO_412 (O_412,N_2762,N_2069);
nand UO_413 (O_413,N_2655,N_2479);
nand UO_414 (O_414,N_2297,N_2891);
nor UO_415 (O_415,N_2554,N_2204);
nor UO_416 (O_416,N_2055,N_2457);
or UO_417 (O_417,N_2300,N_2188);
nand UO_418 (O_418,N_2174,N_2587);
xor UO_419 (O_419,N_2704,N_2185);
nor UO_420 (O_420,N_2804,N_2449);
and UO_421 (O_421,N_2564,N_2890);
nor UO_422 (O_422,N_2914,N_2213);
xnor UO_423 (O_423,N_2984,N_2497);
nor UO_424 (O_424,N_2784,N_2974);
and UO_425 (O_425,N_2593,N_2207);
xor UO_426 (O_426,N_2303,N_2191);
xor UO_427 (O_427,N_2014,N_2466);
xnor UO_428 (O_428,N_2612,N_2907);
or UO_429 (O_429,N_2980,N_2755);
or UO_430 (O_430,N_2674,N_2285);
xnor UO_431 (O_431,N_2775,N_2232);
and UO_432 (O_432,N_2115,N_2508);
and UO_433 (O_433,N_2699,N_2335);
and UO_434 (O_434,N_2040,N_2610);
nor UO_435 (O_435,N_2433,N_2030);
and UO_436 (O_436,N_2813,N_2600);
nand UO_437 (O_437,N_2379,N_2575);
xor UO_438 (O_438,N_2492,N_2552);
and UO_439 (O_439,N_2544,N_2290);
or UO_440 (O_440,N_2981,N_2679);
nor UO_441 (O_441,N_2621,N_2658);
nor UO_442 (O_442,N_2111,N_2973);
or UO_443 (O_443,N_2861,N_2029);
nor UO_444 (O_444,N_2632,N_2148);
and UO_445 (O_445,N_2289,N_2129);
nand UO_446 (O_446,N_2274,N_2436);
xnor UO_447 (O_447,N_2284,N_2720);
and UO_448 (O_448,N_2033,N_2218);
xnor UO_449 (O_449,N_2248,N_2114);
and UO_450 (O_450,N_2998,N_2209);
or UO_451 (O_451,N_2099,N_2885);
xnor UO_452 (O_452,N_2884,N_2849);
and UO_453 (O_453,N_2776,N_2922);
xor UO_454 (O_454,N_2483,N_2256);
xnor UO_455 (O_455,N_2582,N_2324);
and UO_456 (O_456,N_2647,N_2156);
xnor UO_457 (O_457,N_2136,N_2004);
and UO_458 (O_458,N_2145,N_2913);
nor UO_459 (O_459,N_2696,N_2315);
or UO_460 (O_460,N_2105,N_2697);
nand UO_461 (O_461,N_2431,N_2407);
nand UO_462 (O_462,N_2722,N_2440);
nor UO_463 (O_463,N_2745,N_2022);
xnor UO_464 (O_464,N_2533,N_2667);
xor UO_465 (O_465,N_2540,N_2779);
and UO_466 (O_466,N_2294,N_2262);
or UO_467 (O_467,N_2900,N_2613);
and UO_468 (O_468,N_2484,N_2257);
and UO_469 (O_469,N_2782,N_2052);
nor UO_470 (O_470,N_2432,N_2409);
nand UO_471 (O_471,N_2094,N_2282);
nand UO_472 (O_472,N_2601,N_2060);
xnor UO_473 (O_473,N_2986,N_2917);
nor UO_474 (O_474,N_2710,N_2013);
xor UO_475 (O_475,N_2243,N_2146);
or UO_476 (O_476,N_2323,N_2139);
or UO_477 (O_477,N_2260,N_2406);
nand UO_478 (O_478,N_2414,N_2189);
xor UO_479 (O_479,N_2870,N_2451);
and UO_480 (O_480,N_2063,N_2515);
and UO_481 (O_481,N_2987,N_2673);
and UO_482 (O_482,N_2832,N_2242);
or UO_483 (O_483,N_2222,N_2898);
or UO_484 (O_484,N_2769,N_2547);
xor UO_485 (O_485,N_2427,N_2017);
nor UO_486 (O_486,N_2106,N_2444);
and UO_487 (O_487,N_2918,N_2541);
nand UO_488 (O_488,N_2042,N_2147);
nor UO_489 (O_489,N_2585,N_2283);
xnor UO_490 (O_490,N_2557,N_2201);
or UO_491 (O_491,N_2208,N_2850);
nand UO_492 (O_492,N_2685,N_2314);
xnor UO_493 (O_493,N_2749,N_2550);
nor UO_494 (O_494,N_2695,N_2590);
nand UO_495 (O_495,N_2110,N_2151);
and UO_496 (O_496,N_2038,N_2165);
and UO_497 (O_497,N_2978,N_2010);
nor UO_498 (O_498,N_2857,N_2142);
xor UO_499 (O_499,N_2908,N_2510);
endmodule