module basic_1500_15000_2000_10_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_595,In_1130);
nor U1 (N_1,In_1182,In_1085);
or U2 (N_2,In_1140,In_1297);
and U3 (N_3,In_1367,In_22);
nand U4 (N_4,In_1124,In_1242);
nand U5 (N_5,In_173,In_227);
nor U6 (N_6,In_344,In_96);
xnor U7 (N_7,In_457,In_1436);
xor U8 (N_8,In_1307,In_838);
nand U9 (N_9,In_514,In_521);
or U10 (N_10,In_804,In_743);
nand U11 (N_11,In_63,In_978);
nor U12 (N_12,In_477,In_836);
or U13 (N_13,In_2,In_724);
and U14 (N_14,In_175,In_382);
nand U15 (N_15,In_1319,In_852);
xor U16 (N_16,In_1430,In_1334);
and U17 (N_17,In_1168,In_646);
nand U18 (N_18,In_1463,In_592);
nor U19 (N_19,In_15,In_988);
nor U20 (N_20,In_36,In_651);
nand U21 (N_21,In_919,In_768);
nor U22 (N_22,In_594,In_167);
xnor U23 (N_23,In_402,In_327);
or U24 (N_24,In_1,In_814);
nand U25 (N_25,In_587,In_678);
xor U26 (N_26,In_195,In_1070);
or U27 (N_27,In_26,In_1427);
nor U28 (N_28,In_1026,In_278);
nor U29 (N_29,In_722,In_1399);
and U30 (N_30,In_1008,In_1094);
xor U31 (N_31,In_631,In_77);
or U32 (N_32,In_830,In_7);
or U33 (N_33,In_1120,In_259);
and U34 (N_34,In_627,In_757);
or U35 (N_35,In_150,In_95);
and U36 (N_36,In_100,In_276);
nand U37 (N_37,In_650,In_418);
xnor U38 (N_38,In_212,In_356);
xnor U39 (N_39,In_737,In_1386);
and U40 (N_40,In_954,In_1377);
and U41 (N_41,In_380,In_384);
nand U42 (N_42,In_1284,In_1477);
nor U43 (N_43,In_704,In_489);
nor U44 (N_44,In_1429,In_670);
nor U45 (N_45,In_376,In_1300);
nand U46 (N_46,In_1243,In_185);
nand U47 (N_47,In_1178,In_1180);
xnor U48 (N_48,In_80,In_285);
xnor U49 (N_49,In_531,In_107);
nor U50 (N_50,In_471,In_644);
nor U51 (N_51,In_1145,In_741);
nand U52 (N_52,In_624,In_681);
nor U53 (N_53,In_779,In_200);
nand U54 (N_54,In_1425,In_470);
nor U55 (N_55,In_1308,In_186);
nand U56 (N_56,In_949,In_321);
nand U57 (N_57,In_235,In_1495);
or U58 (N_58,In_997,In_536);
or U59 (N_59,In_1002,In_328);
and U60 (N_60,In_4,In_1160);
nor U61 (N_61,In_809,In_1121);
nand U62 (N_62,In_430,In_1318);
nand U63 (N_63,In_220,In_1332);
nand U64 (N_64,In_714,In_1322);
nand U65 (N_65,In_238,In_1460);
or U66 (N_66,In_1195,In_940);
nor U67 (N_67,In_1155,In_144);
and U68 (N_68,In_1150,In_811);
and U69 (N_69,In_142,In_657);
nor U70 (N_70,In_574,In_65);
and U71 (N_71,In_194,In_1447);
and U72 (N_72,In_106,In_796);
nand U73 (N_73,In_744,In_1360);
or U74 (N_74,In_635,In_1281);
or U75 (N_75,In_1207,In_821);
and U76 (N_76,In_441,In_476);
nor U77 (N_77,In_597,In_968);
nand U78 (N_78,In_226,In_46);
and U79 (N_79,In_1456,In_297);
nand U80 (N_80,In_525,In_1376);
or U81 (N_81,In_899,In_456);
or U82 (N_82,In_160,In_1191);
nor U83 (N_83,In_605,In_1273);
and U84 (N_84,In_1470,In_691);
nor U85 (N_85,In_905,In_1383);
and U86 (N_86,In_9,In_1406);
xor U87 (N_87,In_1446,In_1362);
or U88 (N_88,In_926,In_562);
nor U89 (N_89,In_67,In_388);
xor U90 (N_90,In_1415,In_257);
nor U91 (N_91,In_1075,In_1315);
and U92 (N_92,In_892,In_797);
and U93 (N_93,In_964,In_921);
or U94 (N_94,In_172,In_329);
or U95 (N_95,In_295,In_867);
and U96 (N_96,In_1064,In_1489);
nor U97 (N_97,In_783,In_287);
and U98 (N_98,In_707,In_122);
xor U99 (N_99,In_480,In_1363);
or U100 (N_100,In_566,In_519);
nor U101 (N_101,In_951,In_551);
nor U102 (N_102,In_878,In_1053);
nor U103 (N_103,In_1198,In_1230);
nor U104 (N_104,In_213,In_1012);
xnor U105 (N_105,In_1067,In_529);
or U106 (N_106,In_364,In_945);
and U107 (N_107,In_1078,In_452);
nand U108 (N_108,In_1357,In_720);
nor U109 (N_109,In_91,In_740);
or U110 (N_110,In_409,In_166);
or U111 (N_111,In_601,In_1465);
and U112 (N_112,In_1340,In_711);
or U113 (N_113,In_400,In_1074);
nand U114 (N_114,In_101,In_849);
xor U115 (N_115,In_647,In_831);
or U116 (N_116,In_228,In_1439);
nor U117 (N_117,In_206,In_1263);
or U118 (N_118,In_333,In_214);
and U119 (N_119,In_511,In_458);
nand U120 (N_120,In_1077,In_1022);
nand U121 (N_121,In_423,In_1203);
xnor U122 (N_122,In_1431,In_1401);
nand U123 (N_123,In_718,In_170);
nor U124 (N_124,In_338,In_883);
or U125 (N_125,In_346,In_1112);
nor U126 (N_126,In_1143,In_1205);
nand U127 (N_127,In_298,In_1418);
and U128 (N_128,In_370,In_1210);
nand U129 (N_129,In_1073,In_429);
or U130 (N_130,In_1005,In_368);
nor U131 (N_131,In_199,In_1158);
and U132 (N_132,In_974,In_880);
xnor U133 (N_133,In_1040,In_1494);
and U134 (N_134,In_1286,In_1006);
and U135 (N_135,In_1214,In_303);
xnor U136 (N_136,In_588,In_121);
xnor U137 (N_137,In_856,In_19);
and U138 (N_138,In_977,In_469);
or U139 (N_139,In_1048,In_1424);
and U140 (N_140,In_515,In_440);
nand U141 (N_141,In_1434,In_119);
nand U142 (N_142,In_1017,In_62);
and U143 (N_143,In_275,In_729);
or U144 (N_144,In_1096,In_727);
and U145 (N_145,In_1051,In_403);
nand U146 (N_146,In_1353,In_1254);
or U147 (N_147,In_98,In_1468);
xnor U148 (N_148,In_443,In_596);
nor U149 (N_149,In_1234,In_1212);
nand U150 (N_150,In_555,In_911);
nor U151 (N_151,In_1268,In_171);
and U152 (N_152,In_1396,In_1391);
or U153 (N_153,In_25,In_358);
or U154 (N_154,In_1476,In_1084);
or U155 (N_155,In_148,In_985);
or U156 (N_156,In_539,In_1330);
xor U157 (N_157,In_255,In_516);
xnor U158 (N_158,In_349,In_599);
nand U159 (N_159,In_381,In_794);
nand U160 (N_160,In_1335,In_1302);
or U161 (N_161,In_1416,In_967);
nand U162 (N_162,In_1350,In_363);
nand U163 (N_163,In_1147,In_1449);
nor U164 (N_164,In_258,In_558);
nor U165 (N_165,In_820,In_585);
or U166 (N_166,In_1274,In_1080);
nand U167 (N_167,In_1486,In_215);
or U168 (N_168,In_313,In_526);
or U169 (N_169,In_712,In_571);
and U170 (N_170,In_1245,In_270);
and U171 (N_171,In_773,In_475);
or U172 (N_172,In_196,In_941);
or U173 (N_173,In_563,In_850);
nand U174 (N_174,In_94,In_1272);
and U175 (N_175,In_1370,In_732);
and U176 (N_176,In_1271,In_667);
nor U177 (N_177,In_990,In_986);
and U178 (N_178,In_1375,In_554);
or U179 (N_179,In_1090,In_1141);
nand U180 (N_180,In_581,In_372);
and U181 (N_181,In_672,In_948);
nand U182 (N_182,In_1255,In_247);
nor U183 (N_183,In_1410,In_1157);
nor U184 (N_184,In_689,In_626);
nand U185 (N_185,In_580,In_1204);
or U186 (N_186,In_898,In_746);
nand U187 (N_187,In_508,In_696);
nor U188 (N_188,In_1438,In_854);
nand U189 (N_189,In_767,In_318);
nand U190 (N_190,In_1146,In_924);
and U191 (N_191,In_1134,In_896);
and U192 (N_192,In_216,In_161);
nor U193 (N_193,In_556,In_130);
and U194 (N_194,In_1451,In_771);
or U195 (N_195,In_633,In_66);
nand U196 (N_196,In_97,In_618);
or U197 (N_197,In_436,In_791);
nor U198 (N_198,In_404,In_90);
and U199 (N_199,In_345,In_1173);
and U200 (N_200,In_994,In_164);
and U201 (N_201,In_1065,In_1188);
nand U202 (N_202,In_759,In_777);
nor U203 (N_203,In_64,In_1009);
nand U204 (N_204,In_739,In_512);
nand U205 (N_205,In_57,In_132);
and U206 (N_206,In_742,In_1235);
nand U207 (N_207,In_503,In_1052);
or U208 (N_208,In_316,In_1341);
nor U209 (N_209,In_455,In_1221);
nand U210 (N_210,In_1231,In_1260);
or U211 (N_211,In_544,In_638);
or U212 (N_212,In_1079,In_653);
or U213 (N_213,In_352,In_1414);
nor U214 (N_214,In_60,In_156);
and U215 (N_215,In_145,In_396);
nor U216 (N_216,In_1497,In_813);
xnor U217 (N_217,In_801,In_362);
xnor U218 (N_218,In_61,In_643);
and U219 (N_219,In_1232,In_1156);
nor U220 (N_220,In_1384,In_426);
or U221 (N_221,In_1482,In_233);
nand U222 (N_222,In_1473,In_864);
xnor U223 (N_223,In_210,In_1021);
xnor U224 (N_224,In_537,In_890);
xnor U225 (N_225,In_41,In_885);
nor U226 (N_226,In_1305,In_825);
and U227 (N_227,In_1217,In_386);
nand U228 (N_228,In_12,In_187);
nor U229 (N_229,In_1224,In_523);
and U230 (N_230,In_1385,In_420);
or U231 (N_231,In_939,In_583);
nand U232 (N_232,In_760,In_593);
and U233 (N_233,In_659,In_1374);
and U234 (N_234,In_296,In_900);
xor U235 (N_235,In_1445,In_464);
nor U236 (N_236,In_241,In_871);
nor U237 (N_237,In_873,In_1458);
nand U238 (N_238,In_1264,In_1102);
xor U239 (N_239,In_33,In_548);
xor U240 (N_240,In_221,In_1366);
nand U241 (N_241,In_586,In_851);
xor U242 (N_242,In_857,In_1033);
and U243 (N_243,In_218,In_932);
and U244 (N_244,In_942,In_11);
and U245 (N_245,In_394,In_1488);
nand U246 (N_246,In_666,In_474);
xnor U247 (N_247,In_1209,In_1310);
nand U248 (N_248,In_568,In_385);
and U249 (N_249,In_654,In_962);
and U250 (N_250,In_1487,In_855);
nand U251 (N_251,In_365,In_1252);
and U252 (N_252,In_674,In_1337);
nand U253 (N_253,In_800,In_1197);
and U254 (N_254,In_845,In_550);
and U255 (N_255,In_863,In_600);
and U256 (N_256,In_341,In_559);
nor U257 (N_257,In_565,In_472);
nand U258 (N_258,In_553,In_431);
or U259 (N_259,In_1151,In_1136);
nand U260 (N_260,In_1041,In_808);
and U261 (N_261,In_1110,In_0);
xnor U262 (N_262,In_13,In_243);
nor U263 (N_263,In_683,In_294);
and U264 (N_264,In_1276,In_840);
or U265 (N_265,In_1038,In_570);
nor U266 (N_266,In_937,In_591);
or U267 (N_267,In_865,In_1119);
nor U268 (N_268,In_963,In_522);
nor U269 (N_269,In_546,In_427);
and U270 (N_270,In_1139,In_828);
nor U271 (N_271,In_1324,In_279);
nor U272 (N_272,In_127,In_909);
nand U273 (N_273,In_782,In_961);
or U274 (N_274,In_648,In_695);
and U275 (N_275,In_438,In_1405);
or U276 (N_276,In_1059,In_24);
and U277 (N_277,In_753,In_378);
or U278 (N_278,In_1251,In_1450);
nor U279 (N_279,In_182,In_658);
xnor U280 (N_280,In_1138,In_1037);
nor U281 (N_281,In_151,In_1089);
or U282 (N_282,In_645,In_1137);
nor U283 (N_283,In_1201,In_157);
and U284 (N_284,In_1149,In_752);
nand U285 (N_285,In_280,In_1492);
xnor U286 (N_286,In_834,In_1423);
and U287 (N_287,In_611,In_1083);
nor U288 (N_288,In_697,In_882);
nor U289 (N_289,In_787,In_334);
and U290 (N_290,In_518,In_35);
or U291 (N_291,In_675,In_1480);
and U292 (N_292,In_224,In_128);
nand U293 (N_293,In_219,In_1013);
nand U294 (N_294,In_1219,In_884);
or U295 (N_295,In_922,In_314);
and U296 (N_296,In_1199,In_823);
and U297 (N_297,In_223,In_1154);
nand U298 (N_298,In_904,In_1298);
nand U299 (N_299,In_506,In_609);
nand U300 (N_300,In_290,In_561);
and U301 (N_301,In_110,In_21);
or U302 (N_302,In_293,In_1250);
or U303 (N_303,In_299,In_108);
and U304 (N_304,In_973,In_676);
and U305 (N_305,In_1400,In_958);
and U306 (N_306,In_894,In_459);
nand U307 (N_307,In_143,In_1356);
nand U308 (N_308,In_1166,In_463);
nand U309 (N_309,In_615,In_640);
and U310 (N_310,In_578,In_10);
and U311 (N_311,In_414,In_1211);
nor U312 (N_312,In_50,In_1227);
nor U313 (N_313,In_237,In_982);
or U314 (N_314,In_168,In_1082);
or U315 (N_315,In_509,In_861);
or U316 (N_316,In_844,In_114);
and U317 (N_317,In_750,In_495);
and U318 (N_318,In_342,In_39);
nor U319 (N_319,In_661,In_54);
and U320 (N_320,In_1411,In_590);
nand U321 (N_321,In_309,In_513);
and U322 (N_322,In_542,In_826);
nor U323 (N_323,In_1010,In_913);
and U324 (N_324,In_1389,In_662);
nand U325 (N_325,In_1185,In_1057);
nor U326 (N_326,In_282,In_795);
or U327 (N_327,In_879,In_1311);
nor U328 (N_328,In_895,In_184);
or U329 (N_329,In_231,In_68);
or U330 (N_330,In_728,In_573);
xor U331 (N_331,In_1184,In_792);
and U332 (N_332,In_1233,In_1056);
or U333 (N_333,In_319,In_250);
xnor U334 (N_334,In_1175,In_209);
nor U335 (N_335,In_154,In_1493);
xnor U336 (N_336,In_1003,In_1426);
xor U337 (N_337,In_1379,In_876);
nand U338 (N_338,In_639,In_1348);
or U339 (N_339,In_162,In_869);
xor U340 (N_340,In_1131,In_907);
and U341 (N_341,In_1034,In_118);
or U342 (N_342,In_802,In_607);
or U343 (N_343,In_1000,In_1265);
nor U344 (N_344,In_1179,In_306);
nand U345 (N_345,In_85,In_222);
nor U346 (N_346,In_421,In_240);
xnor U347 (N_347,In_625,In_1444);
nand U348 (N_348,In_283,In_1291);
xnor U349 (N_349,In_1479,In_1317);
nor U350 (N_350,In_541,In_1023);
and U351 (N_351,In_762,In_159);
or U352 (N_352,In_415,In_311);
and U353 (N_353,In_776,In_1100);
and U354 (N_354,In_693,In_189);
nor U355 (N_355,In_908,In_1187);
xnor U356 (N_356,In_103,In_938);
nor U357 (N_357,In_1485,In_1448);
nor U358 (N_358,In_266,In_82);
and U359 (N_359,In_286,In_636);
nand U360 (N_360,In_972,In_1129);
nor U361 (N_361,In_367,In_1111);
xnor U362 (N_362,In_824,In_1229);
xnor U363 (N_363,In_843,In_608);
nand U364 (N_364,In_1464,In_866);
and U365 (N_365,In_304,In_1466);
nor U366 (N_366,In_976,In_960);
nor U367 (N_367,In_1279,In_500);
xnor U368 (N_368,In_793,In_970);
and U369 (N_369,In_910,In_398);
or U370 (N_370,In_956,In_407);
nor U371 (N_371,In_999,In_383);
nor U372 (N_372,In_897,In_1413);
nor U373 (N_373,In_72,In_181);
nor U374 (N_374,In_950,In_1177);
nand U375 (N_375,In_450,In_133);
or U376 (N_376,In_1469,In_1314);
nor U377 (N_377,In_1270,In_390);
nor U378 (N_378,In_1398,In_1359);
nor U379 (N_379,In_564,In_1164);
and U380 (N_380,In_1001,In_798);
or U381 (N_381,In_1301,In_139);
xnor U382 (N_382,In_1196,In_620);
nand U383 (N_383,In_351,In_113);
nor U384 (N_384,In_579,In_1194);
nor U385 (N_385,In_770,In_1043);
or U386 (N_386,In_694,In_389);
xor U387 (N_387,In_1382,In_702);
nand U388 (N_388,In_485,In_373);
or U389 (N_389,In_1381,In_59);
nand U390 (N_390,In_253,In_1088);
and U391 (N_391,In_229,In_1031);
and U392 (N_392,In_131,In_393);
or U393 (N_393,In_1351,In_1186);
nand U394 (N_394,In_460,In_395);
nand U395 (N_395,In_1290,In_315);
or U396 (N_396,In_174,In_687);
or U397 (N_397,In_629,In_1069);
nand U398 (N_398,In_769,In_262);
nor U399 (N_399,In_134,In_481);
nand U400 (N_400,In_1393,In_507);
nor U401 (N_401,In_641,In_1039);
or U402 (N_402,In_682,In_354);
or U403 (N_403,In_1020,In_102);
nor U404 (N_404,In_1115,In_1066);
or U405 (N_405,In_140,In_1228);
or U406 (N_406,In_547,In_1461);
and U407 (N_407,In_1299,In_630);
nand U408 (N_408,In_211,In_355);
and U409 (N_409,In_731,In_1365);
nand U410 (N_410,In_991,In_252);
nand U411 (N_411,In_291,In_392);
nand U412 (N_412,In_331,In_466);
and U413 (N_413,In_1371,In_527);
xnor U414 (N_414,In_273,In_1086);
nand U415 (N_415,In_83,In_339);
nand U416 (N_416,In_621,In_1108);
or U417 (N_417,In_1262,In_1135);
nand U418 (N_418,In_14,In_842);
and U419 (N_419,In_628,In_330);
or U420 (N_420,In_1126,In_1035);
nor U421 (N_421,In_1117,In_86);
or U422 (N_422,In_264,In_1433);
nand U423 (N_423,In_1257,In_1174);
xnor U424 (N_424,In_971,In_141);
nand U425 (N_425,In_419,In_366);
nor U426 (N_426,In_1481,In_505);
and U427 (N_427,In_572,In_188);
nand U428 (N_428,In_923,In_1285);
and U429 (N_429,In_1170,In_806);
xor U430 (N_430,In_1435,In_428);
and U431 (N_431,In_1123,In_69);
nand U432 (N_432,In_934,In_302);
nand U433 (N_433,In_1459,In_781);
nor U434 (N_434,In_1215,In_493);
xor U435 (N_435,In_176,In_20);
or U436 (N_436,In_263,In_1068);
nor U437 (N_437,In_1030,In_1019);
and U438 (N_438,In_129,In_391);
or U439 (N_439,In_1183,In_818);
nand U440 (N_440,In_1213,In_78);
and U441 (N_441,In_766,In_685);
nor U442 (N_442,In_1133,In_747);
nand U443 (N_443,In_1327,In_205);
and U444 (N_444,In_325,In_55);
and U445 (N_445,In_1058,In_1256);
nand U446 (N_446,In_178,In_467);
or U447 (N_447,In_320,In_946);
nor U448 (N_448,In_668,In_1428);
nand U449 (N_449,In_112,In_163);
xor U450 (N_450,In_730,In_853);
or U451 (N_451,In_1397,In_260);
nor U452 (N_452,In_1113,In_1192);
and U453 (N_453,In_1333,In_560);
and U454 (N_454,In_1062,In_528);
nor U455 (N_455,In_817,In_1127);
nor U456 (N_456,In_989,In_56);
nor U457 (N_457,In_272,In_534);
or U458 (N_458,In_785,In_1453);
and U459 (N_459,In_716,In_520);
nand U460 (N_460,In_758,In_765);
nor U461 (N_461,In_288,In_1025);
nor U462 (N_462,In_761,In_1246);
nand U463 (N_463,In_952,In_1422);
and U464 (N_464,In_755,In_1189);
nand U465 (N_465,In_16,In_1338);
nand U466 (N_466,In_417,In_1325);
nand U467 (N_467,In_1220,In_17);
nand U468 (N_468,In_1364,In_1159);
and U469 (N_469,In_708,In_987);
nor U470 (N_470,In_28,In_1015);
nand U471 (N_471,In_269,In_837);
nor U472 (N_472,In_772,In_52);
nor U473 (N_473,In_204,In_1114);
or U474 (N_474,In_268,In_444);
nand U475 (N_475,In_679,In_669);
and U476 (N_476,In_317,In_87);
nand U477 (N_477,In_925,In_1046);
xor U478 (N_478,In_931,In_1283);
nand U479 (N_479,In_1063,In_6);
xor U480 (N_480,In_723,In_1498);
or U481 (N_481,In_575,In_775);
nand U482 (N_482,In_891,In_1467);
and U483 (N_483,In_197,In_1420);
or U484 (N_484,In_74,In_893);
nor U485 (N_485,In_790,In_401);
nand U486 (N_486,In_1152,In_610);
or U487 (N_487,In_535,In_589);
nor U488 (N_488,In_335,In_1060);
or U489 (N_489,In_735,In_1355);
and U490 (N_490,In_498,In_1372);
or U491 (N_491,In_1225,In_684);
nand U492 (N_492,In_677,In_1095);
or U493 (N_493,In_18,In_369);
nand U494 (N_494,In_120,In_998);
xor U495 (N_495,In_1253,In_1047);
or U496 (N_496,In_1472,In_225);
nand U497 (N_497,In_815,In_1239);
and U498 (N_498,In_917,In_501);
xor U499 (N_499,In_1167,In_1216);
and U500 (N_500,In_680,In_1144);
nor U501 (N_501,In_265,In_715);
or U502 (N_502,In_245,In_721);
and U503 (N_503,In_552,In_875);
xor U504 (N_504,In_31,In_1161);
and U505 (N_505,In_1107,In_1148);
nor U506 (N_506,In_73,In_690);
nand U507 (N_507,In_1091,In_1104);
or U508 (N_508,In_1105,In_1101);
xor U509 (N_509,In_51,In_374);
nand U510 (N_510,In_1087,In_8);
and U511 (N_511,In_499,In_149);
nor U512 (N_512,In_347,In_1471);
nor U513 (N_513,In_123,In_1172);
nor U514 (N_514,In_1269,In_1326);
and U515 (N_515,In_359,In_432);
or U516 (N_516,In_1238,In_482);
nor U517 (N_517,In_435,In_1499);
nand U518 (N_518,In_256,In_111);
nor U519 (N_519,In_191,In_710);
or U520 (N_520,In_343,In_1044);
nor U521 (N_521,In_701,In_1442);
nand U522 (N_522,In_902,In_1496);
nor U523 (N_523,In_1118,In_816);
or U524 (N_524,In_1347,In_84);
nor U525 (N_525,In_397,In_1014);
xnor U526 (N_526,In_1241,In_439);
nand U527 (N_527,In_1304,In_230);
or U528 (N_528,In_545,In_289);
nor U529 (N_529,In_901,In_1027);
nand U530 (N_530,In_1387,In_447);
xor U531 (N_531,In_993,In_789);
nor U532 (N_532,In_966,In_350);
nor U533 (N_533,In_38,In_1153);
or U534 (N_534,In_524,In_835);
nor U535 (N_535,In_706,In_207);
and U536 (N_536,In_981,In_1412);
nor U537 (N_537,In_115,In_357);
or U538 (N_538,In_1097,In_424);
or U539 (N_539,In_445,In_203);
xor U540 (N_540,In_336,In_468);
nor U541 (N_541,In_1004,In_1050);
nand U542 (N_542,In_872,In_652);
and U543 (N_543,In_619,In_1054);
nor U544 (N_544,In_557,In_75);
or U545 (N_545,In_705,In_881);
nand U546 (N_546,In_935,In_569);
nor U547 (N_547,In_969,In_1061);
and U548 (N_548,In_37,In_292);
and U549 (N_549,In_664,In_125);
and U550 (N_550,In_1344,In_584);
xor U551 (N_551,In_1349,In_1282);
or U552 (N_552,In_1457,In_1042);
nor U553 (N_553,In_1259,In_606);
xnor U554 (N_554,In_217,In_944);
nor U555 (N_555,In_312,In_1028);
nor U556 (N_556,In_877,In_1474);
nand U557 (N_557,In_1202,In_846);
nor U558 (N_558,In_124,In_190);
or U559 (N_559,In_153,In_726);
nand U560 (N_560,In_1128,In_784);
or U561 (N_561,In_612,In_324);
and U562 (N_562,In_478,In_44);
and U563 (N_563,In_1358,In_1103);
nor U564 (N_564,In_1122,In_248);
or U565 (N_565,In_617,In_76);
or U566 (N_566,In_1029,In_254);
or U567 (N_567,In_451,In_99);
nand U568 (N_568,In_1267,In_660);
or U569 (N_569,In_42,In_1024);
nor U570 (N_570,In_576,In_30);
nand U571 (N_571,In_604,In_1277);
or U572 (N_572,In_138,In_437);
nand U573 (N_573,In_688,In_58);
nor U574 (N_574,In_408,In_1419);
nand U575 (N_575,In_713,In_700);
nand U576 (N_576,In_92,In_959);
nand U577 (N_577,In_927,In_249);
nor U578 (N_578,In_267,In_332);
nand U579 (N_579,In_1490,In_137);
nor U580 (N_580,In_996,In_1484);
and U581 (N_581,In_1380,In_1171);
or U582 (N_582,In_1045,In_399);
and U583 (N_583,In_48,In_751);
or U584 (N_584,In_847,In_947);
and U585 (N_585,In_1395,In_1222);
or U586 (N_586,In_860,In_839);
nand U587 (N_587,In_780,In_1373);
nand U588 (N_588,In_870,In_433);
and U589 (N_589,In_868,In_81);
xor U590 (N_590,In_1011,In_1441);
nor U591 (N_591,In_1266,In_1226);
or U592 (N_592,In_1336,In_1176);
and U593 (N_593,In_208,In_244);
or U594 (N_594,In_1258,In_819);
or U595 (N_595,In_656,In_1249);
or U596 (N_596,In_1352,In_23);
xnor U597 (N_597,In_271,In_116);
and U598 (N_598,In_337,In_105);
or U599 (N_599,In_920,In_916);
or U600 (N_600,In_32,In_1165);
or U601 (N_601,In_655,In_5);
or U602 (N_602,In_165,In_1236);
or U603 (N_603,In_1193,In_242);
nand U604 (N_604,In_918,In_749);
or U605 (N_605,In_692,In_799);
xnor U606 (N_606,In_461,In_858);
and U607 (N_607,In_45,In_530);
nand U608 (N_608,In_305,In_1392);
xnor U609 (N_609,In_1218,In_487);
and U610 (N_610,In_169,In_301);
and U611 (N_611,In_27,In_1142);
nand U612 (N_612,In_549,In_377);
and U613 (N_613,In_915,In_1443);
and U614 (N_614,In_89,In_486);
nor U615 (N_615,In_1163,In_488);
xor U616 (N_616,In_1071,In_1288);
and U617 (N_617,In_832,In_1346);
xnor U618 (N_618,In_1125,In_109);
or U619 (N_619,In_179,In_1407);
or U620 (N_620,In_53,In_1437);
or U621 (N_621,In_40,In_928);
nand U622 (N_622,In_413,In_841);
or U623 (N_623,In_1394,In_829);
nand U624 (N_624,In_719,In_284);
and U625 (N_625,In_155,In_454);
or U626 (N_626,In_1289,In_239);
nor U627 (N_627,In_1478,In_502);
nor U628 (N_628,In_126,In_1109);
nor U629 (N_629,In_1321,In_1390);
or U630 (N_630,In_1016,In_953);
or U631 (N_631,In_361,In_492);
nand U632 (N_632,In_326,In_494);
xnor U633 (N_633,In_807,In_533);
or U634 (N_634,In_634,In_745);
and U635 (N_635,In_43,In_71);
nand U636 (N_636,In_567,In_980);
or U637 (N_637,In_490,In_1007);
nand U638 (N_638,In_387,In_642);
xnor U639 (N_639,In_1275,In_774);
nor U640 (N_640,In_1296,In_1036);
nand U641 (N_641,In_425,In_277);
and U642 (N_642,In_379,In_274);
or U643 (N_643,In_827,In_754);
nor U644 (N_644,In_202,In_34);
nor U645 (N_645,In_1329,In_406);
or U646 (N_646,In_79,In_1404);
and U647 (N_647,In_1206,In_1181);
and U648 (N_648,In_183,In_308);
nand U649 (N_649,In_1368,In_1018);
or U650 (N_650,In_717,In_889);
and U651 (N_651,In_348,In_1316);
and U652 (N_652,In_803,In_422);
or U653 (N_653,In_975,In_698);
nand U654 (N_654,In_543,In_788);
nand U655 (N_655,In_323,In_446);
or U656 (N_656,In_632,In_1452);
nor U657 (N_657,In_538,In_3);
nand U658 (N_658,In_180,In_906);
xor U659 (N_659,In_251,In_1076);
or U660 (N_660,In_434,In_859);
or U661 (N_661,In_483,In_577);
nand U662 (N_662,In_903,In_1278);
nand U663 (N_663,In_1099,In_1200);
and U664 (N_664,In_193,In_1081);
nand U665 (N_665,In_497,In_614);
or U666 (N_666,In_637,In_1354);
nand U667 (N_667,In_371,In_147);
nand U668 (N_668,In_1293,In_1032);
and U669 (N_669,In_353,In_410);
nand U670 (N_670,In_613,In_1421);
or U671 (N_671,In_862,In_957);
nor U672 (N_672,In_686,In_93);
xnor U673 (N_673,In_1055,In_1312);
nand U674 (N_674,In_484,In_411);
or U675 (N_675,In_47,In_232);
or U676 (N_676,In_360,In_699);
or U677 (N_677,In_146,In_1106);
or U678 (N_678,In_491,In_887);
or U679 (N_679,In_1361,In_602);
nand U680 (N_680,In_1223,In_1132);
nand U681 (N_681,In_763,In_1049);
or U682 (N_682,In_1303,In_416);
xor U683 (N_683,In_822,In_152);
and U684 (N_684,In_504,In_812);
or U685 (N_685,In_1462,In_340);
and U686 (N_686,In_738,In_1208);
nand U687 (N_687,In_736,In_810);
xor U688 (N_688,In_1093,In_1320);
or U689 (N_689,In_510,In_1295);
or U690 (N_690,In_448,In_1247);
nor U691 (N_691,In_70,In_733);
nor U692 (N_692,In_805,In_1440);
and U693 (N_693,In_1432,In_1323);
xnor U694 (N_694,In_848,In_449);
nor U695 (N_695,In_1190,In_1280);
or U696 (N_696,In_914,In_673);
nand U697 (N_697,In_1328,In_1331);
nor U698 (N_698,In_929,In_192);
and U699 (N_699,In_1483,In_1343);
nor U700 (N_700,In_236,In_496);
or U701 (N_701,In_1116,In_1408);
and U702 (N_702,In_1342,In_1072);
nor U703 (N_703,In_1455,In_1339);
xor U704 (N_704,In_104,In_933);
xor U705 (N_705,In_1287,In_158);
nor U706 (N_706,In_912,In_540);
or U707 (N_707,In_983,In_665);
nor U708 (N_708,In_300,In_649);
nor U709 (N_709,In_1403,In_833);
or U710 (N_710,In_1369,In_1491);
or U711 (N_711,In_1261,In_1475);
nand U712 (N_712,In_49,In_453);
nand U713 (N_713,In_874,In_622);
nand U714 (N_714,In_778,In_995);
nand U715 (N_715,In_936,In_1345);
and U716 (N_716,In_703,In_756);
and U717 (N_717,In_135,In_748);
xor U718 (N_718,In_955,In_517);
or U719 (N_719,In_281,In_582);
or U720 (N_720,In_405,In_1309);
and U721 (N_721,In_1237,In_992);
nor U722 (N_722,In_623,In_462);
nor U723 (N_723,In_375,In_1402);
and U724 (N_724,In_532,In_1388);
nand U725 (N_725,In_234,In_1092);
and U726 (N_726,In_1292,In_663);
nand U727 (N_727,In_465,In_88);
or U728 (N_728,In_888,In_764);
nor U729 (N_729,In_198,In_1248);
or U730 (N_730,In_943,In_136);
nor U731 (N_731,In_1294,In_246);
nand U732 (N_732,In_930,In_1378);
xnor U733 (N_733,In_1098,In_1409);
nand U734 (N_734,In_117,In_598);
or U735 (N_735,In_886,In_473);
or U736 (N_736,In_965,In_734);
nand U737 (N_737,In_1169,In_1306);
and U738 (N_738,In_1162,In_786);
nand U739 (N_739,In_322,In_442);
nor U740 (N_740,In_979,In_479);
or U741 (N_741,In_177,In_603);
and U742 (N_742,In_725,In_201);
nor U743 (N_743,In_1417,In_310);
nand U744 (N_744,In_412,In_1313);
nand U745 (N_745,In_984,In_709);
nand U746 (N_746,In_29,In_1244);
and U747 (N_747,In_1454,In_1240);
or U748 (N_748,In_261,In_307);
and U749 (N_749,In_616,In_671);
and U750 (N_750,In_1269,In_1104);
and U751 (N_751,In_1167,In_285);
nand U752 (N_752,In_616,In_905);
and U753 (N_753,In_1402,In_1294);
and U754 (N_754,In_1202,In_179);
nor U755 (N_755,In_689,In_106);
nor U756 (N_756,In_206,In_1099);
nor U757 (N_757,In_673,In_251);
or U758 (N_758,In_432,In_709);
and U759 (N_759,In_379,In_701);
nor U760 (N_760,In_669,In_831);
nor U761 (N_761,In_353,In_1364);
or U762 (N_762,In_1268,In_215);
or U763 (N_763,In_755,In_1324);
and U764 (N_764,In_343,In_815);
nor U765 (N_765,In_1439,In_705);
xnor U766 (N_766,In_1444,In_1391);
and U767 (N_767,In_1297,In_666);
nor U768 (N_768,In_503,In_1459);
and U769 (N_769,In_686,In_478);
nor U770 (N_770,In_148,In_730);
nor U771 (N_771,In_507,In_538);
nand U772 (N_772,In_585,In_571);
xnor U773 (N_773,In_862,In_705);
nor U774 (N_774,In_86,In_1200);
nand U775 (N_775,In_629,In_197);
and U776 (N_776,In_95,In_1163);
or U777 (N_777,In_1160,In_99);
or U778 (N_778,In_692,In_581);
xnor U779 (N_779,In_877,In_1456);
or U780 (N_780,In_1296,In_1265);
nand U781 (N_781,In_1416,In_258);
nand U782 (N_782,In_1229,In_257);
nand U783 (N_783,In_1266,In_319);
nand U784 (N_784,In_491,In_135);
and U785 (N_785,In_483,In_1138);
nor U786 (N_786,In_389,In_495);
and U787 (N_787,In_930,In_945);
and U788 (N_788,In_314,In_375);
nand U789 (N_789,In_1369,In_904);
nand U790 (N_790,In_367,In_656);
nor U791 (N_791,In_80,In_425);
nand U792 (N_792,In_114,In_339);
and U793 (N_793,In_85,In_1364);
and U794 (N_794,In_1299,In_936);
or U795 (N_795,In_463,In_1173);
nand U796 (N_796,In_72,In_213);
or U797 (N_797,In_93,In_561);
nor U798 (N_798,In_1498,In_462);
nor U799 (N_799,In_171,In_342);
nand U800 (N_800,In_229,In_692);
nand U801 (N_801,In_1398,In_794);
and U802 (N_802,In_486,In_248);
nor U803 (N_803,In_633,In_176);
or U804 (N_804,In_330,In_1052);
nand U805 (N_805,In_606,In_1064);
and U806 (N_806,In_1313,In_117);
and U807 (N_807,In_1299,In_834);
and U808 (N_808,In_993,In_1462);
or U809 (N_809,In_602,In_655);
nor U810 (N_810,In_599,In_430);
or U811 (N_811,In_151,In_361);
xor U812 (N_812,In_1372,In_1284);
nand U813 (N_813,In_451,In_1237);
or U814 (N_814,In_352,In_328);
nor U815 (N_815,In_691,In_351);
nand U816 (N_816,In_116,In_672);
or U817 (N_817,In_1209,In_556);
and U818 (N_818,In_1233,In_1405);
or U819 (N_819,In_1175,In_979);
nor U820 (N_820,In_689,In_1433);
or U821 (N_821,In_1334,In_445);
or U822 (N_822,In_1106,In_644);
or U823 (N_823,In_1165,In_914);
nor U824 (N_824,In_556,In_191);
and U825 (N_825,In_115,In_1330);
nand U826 (N_826,In_682,In_1236);
or U827 (N_827,In_476,In_757);
or U828 (N_828,In_700,In_45);
nand U829 (N_829,In_297,In_404);
and U830 (N_830,In_723,In_27);
xor U831 (N_831,In_761,In_1336);
nor U832 (N_832,In_410,In_1472);
nand U833 (N_833,In_926,In_623);
and U834 (N_834,In_698,In_1342);
nand U835 (N_835,In_715,In_1145);
or U836 (N_836,In_508,In_1237);
or U837 (N_837,In_922,In_512);
nand U838 (N_838,In_713,In_601);
nand U839 (N_839,In_732,In_1451);
and U840 (N_840,In_288,In_249);
nand U841 (N_841,In_358,In_835);
nand U842 (N_842,In_616,In_923);
nand U843 (N_843,In_1388,In_892);
nor U844 (N_844,In_314,In_1228);
or U845 (N_845,In_761,In_821);
nand U846 (N_846,In_936,In_644);
nand U847 (N_847,In_747,In_462);
and U848 (N_848,In_1247,In_654);
nor U849 (N_849,In_423,In_204);
nand U850 (N_850,In_632,In_726);
nand U851 (N_851,In_1312,In_280);
nand U852 (N_852,In_142,In_56);
and U853 (N_853,In_383,In_159);
nor U854 (N_854,In_717,In_799);
xnor U855 (N_855,In_618,In_232);
or U856 (N_856,In_478,In_1102);
nor U857 (N_857,In_51,In_1184);
nor U858 (N_858,In_396,In_972);
nor U859 (N_859,In_1280,In_522);
and U860 (N_860,In_237,In_875);
and U861 (N_861,In_644,In_173);
xor U862 (N_862,In_505,In_778);
or U863 (N_863,In_1434,In_956);
nor U864 (N_864,In_872,In_1110);
and U865 (N_865,In_294,In_641);
or U866 (N_866,In_214,In_122);
nand U867 (N_867,In_87,In_1308);
nor U868 (N_868,In_1389,In_238);
nor U869 (N_869,In_404,In_474);
nand U870 (N_870,In_206,In_988);
or U871 (N_871,In_163,In_545);
or U872 (N_872,In_18,In_255);
nand U873 (N_873,In_802,In_579);
and U874 (N_874,In_84,In_770);
and U875 (N_875,In_278,In_1012);
nand U876 (N_876,In_791,In_535);
nand U877 (N_877,In_1360,In_1106);
xor U878 (N_878,In_545,In_5);
xor U879 (N_879,In_566,In_1084);
and U880 (N_880,In_297,In_335);
nor U881 (N_881,In_1259,In_1397);
and U882 (N_882,In_538,In_1105);
nand U883 (N_883,In_321,In_735);
and U884 (N_884,In_917,In_146);
or U885 (N_885,In_825,In_934);
nor U886 (N_886,In_951,In_1369);
nor U887 (N_887,In_462,In_988);
or U888 (N_888,In_288,In_475);
or U889 (N_889,In_372,In_830);
xnor U890 (N_890,In_935,In_1260);
nor U891 (N_891,In_1091,In_879);
nand U892 (N_892,In_395,In_524);
nor U893 (N_893,In_517,In_930);
and U894 (N_894,In_830,In_709);
or U895 (N_895,In_212,In_721);
and U896 (N_896,In_78,In_79);
or U897 (N_897,In_1244,In_585);
nand U898 (N_898,In_440,In_816);
or U899 (N_899,In_60,In_204);
xnor U900 (N_900,In_1328,In_135);
or U901 (N_901,In_78,In_400);
or U902 (N_902,In_1094,In_1207);
or U903 (N_903,In_9,In_71);
nor U904 (N_904,In_579,In_950);
nand U905 (N_905,In_1383,In_240);
and U906 (N_906,In_420,In_1086);
or U907 (N_907,In_1130,In_1168);
or U908 (N_908,In_495,In_552);
nor U909 (N_909,In_914,In_1171);
and U910 (N_910,In_893,In_718);
nor U911 (N_911,In_828,In_803);
nor U912 (N_912,In_587,In_400);
nand U913 (N_913,In_432,In_1020);
and U914 (N_914,In_1107,In_1096);
and U915 (N_915,In_93,In_203);
xor U916 (N_916,In_598,In_1107);
or U917 (N_917,In_900,In_1225);
nand U918 (N_918,In_488,In_1329);
and U919 (N_919,In_1154,In_495);
and U920 (N_920,In_1206,In_1458);
and U921 (N_921,In_272,In_318);
and U922 (N_922,In_1218,In_966);
nor U923 (N_923,In_1109,In_180);
and U924 (N_924,In_358,In_1489);
or U925 (N_925,In_1433,In_630);
or U926 (N_926,In_6,In_34);
nor U927 (N_927,In_407,In_694);
and U928 (N_928,In_691,In_1072);
nand U929 (N_929,In_159,In_843);
nand U930 (N_930,In_248,In_150);
xor U931 (N_931,In_553,In_1010);
and U932 (N_932,In_1137,In_994);
xor U933 (N_933,In_1431,In_504);
xor U934 (N_934,In_901,In_697);
and U935 (N_935,In_214,In_686);
nor U936 (N_936,In_999,In_16);
and U937 (N_937,In_214,In_1242);
and U938 (N_938,In_541,In_843);
and U939 (N_939,In_1409,In_726);
nand U940 (N_940,In_535,In_1354);
and U941 (N_941,In_776,In_1035);
and U942 (N_942,In_473,In_76);
or U943 (N_943,In_141,In_378);
and U944 (N_944,In_441,In_1233);
nand U945 (N_945,In_1424,In_1434);
and U946 (N_946,In_43,In_411);
and U947 (N_947,In_86,In_185);
nand U948 (N_948,In_864,In_352);
nand U949 (N_949,In_554,In_1064);
nor U950 (N_950,In_419,In_823);
and U951 (N_951,In_1486,In_293);
and U952 (N_952,In_218,In_1278);
nand U953 (N_953,In_269,In_927);
nor U954 (N_954,In_1466,In_126);
nand U955 (N_955,In_310,In_652);
nand U956 (N_956,In_1248,In_1229);
or U957 (N_957,In_1121,In_901);
nor U958 (N_958,In_914,In_257);
nand U959 (N_959,In_861,In_483);
nand U960 (N_960,In_44,In_672);
nor U961 (N_961,In_544,In_334);
nand U962 (N_962,In_202,In_559);
xor U963 (N_963,In_1455,In_194);
or U964 (N_964,In_302,In_1466);
nor U965 (N_965,In_785,In_381);
and U966 (N_966,In_2,In_1258);
and U967 (N_967,In_255,In_1047);
and U968 (N_968,In_264,In_59);
or U969 (N_969,In_691,In_1001);
nor U970 (N_970,In_851,In_1449);
or U971 (N_971,In_479,In_1106);
xor U972 (N_972,In_1,In_769);
or U973 (N_973,In_1071,In_1304);
or U974 (N_974,In_120,In_1349);
or U975 (N_975,In_771,In_44);
or U976 (N_976,In_34,In_965);
xor U977 (N_977,In_1410,In_982);
nor U978 (N_978,In_1061,In_648);
xnor U979 (N_979,In_196,In_347);
nor U980 (N_980,In_304,In_80);
and U981 (N_981,In_248,In_1178);
xnor U982 (N_982,In_819,In_441);
or U983 (N_983,In_285,In_1108);
nor U984 (N_984,In_405,In_869);
nand U985 (N_985,In_318,In_79);
xor U986 (N_986,In_815,In_573);
nand U987 (N_987,In_895,In_1430);
and U988 (N_988,In_340,In_582);
and U989 (N_989,In_288,In_627);
or U990 (N_990,In_1107,In_1349);
nor U991 (N_991,In_1483,In_711);
and U992 (N_992,In_1396,In_162);
nor U993 (N_993,In_155,In_901);
nor U994 (N_994,In_1094,In_281);
and U995 (N_995,In_819,In_98);
or U996 (N_996,In_365,In_589);
nor U997 (N_997,In_1288,In_1471);
or U998 (N_998,In_926,In_608);
nor U999 (N_999,In_684,In_42);
nor U1000 (N_1000,In_184,In_1109);
or U1001 (N_1001,In_982,In_867);
or U1002 (N_1002,In_811,In_362);
and U1003 (N_1003,In_594,In_801);
nor U1004 (N_1004,In_1178,In_62);
nor U1005 (N_1005,In_1070,In_320);
nand U1006 (N_1006,In_1049,In_249);
or U1007 (N_1007,In_1239,In_348);
nand U1008 (N_1008,In_270,In_350);
and U1009 (N_1009,In_1398,In_655);
nor U1010 (N_1010,In_757,In_799);
nand U1011 (N_1011,In_1223,In_1224);
or U1012 (N_1012,In_163,In_990);
or U1013 (N_1013,In_944,In_402);
and U1014 (N_1014,In_257,In_763);
and U1015 (N_1015,In_681,In_1223);
nand U1016 (N_1016,In_832,In_344);
xor U1017 (N_1017,In_1317,In_1092);
nand U1018 (N_1018,In_401,In_783);
nand U1019 (N_1019,In_1227,In_651);
and U1020 (N_1020,In_990,In_152);
or U1021 (N_1021,In_225,In_60);
or U1022 (N_1022,In_353,In_998);
nand U1023 (N_1023,In_455,In_152);
nand U1024 (N_1024,In_1465,In_1295);
xnor U1025 (N_1025,In_425,In_802);
nor U1026 (N_1026,In_1204,In_30);
and U1027 (N_1027,In_5,In_1272);
or U1028 (N_1028,In_638,In_1074);
or U1029 (N_1029,In_185,In_934);
nor U1030 (N_1030,In_790,In_37);
nor U1031 (N_1031,In_499,In_857);
nand U1032 (N_1032,In_1106,In_1009);
and U1033 (N_1033,In_1252,In_878);
or U1034 (N_1034,In_1265,In_1157);
and U1035 (N_1035,In_713,In_826);
or U1036 (N_1036,In_1130,In_472);
or U1037 (N_1037,In_348,In_206);
or U1038 (N_1038,In_609,In_38);
or U1039 (N_1039,In_303,In_1163);
nor U1040 (N_1040,In_1371,In_1350);
nand U1041 (N_1041,In_833,In_897);
xnor U1042 (N_1042,In_832,In_725);
or U1043 (N_1043,In_1393,In_1207);
and U1044 (N_1044,In_680,In_976);
xnor U1045 (N_1045,In_1155,In_810);
or U1046 (N_1046,In_1056,In_1295);
nor U1047 (N_1047,In_503,In_572);
and U1048 (N_1048,In_733,In_998);
xnor U1049 (N_1049,In_807,In_1281);
nor U1050 (N_1050,In_1290,In_1485);
nand U1051 (N_1051,In_621,In_653);
and U1052 (N_1052,In_247,In_1236);
and U1053 (N_1053,In_1032,In_873);
xor U1054 (N_1054,In_136,In_859);
and U1055 (N_1055,In_379,In_303);
nand U1056 (N_1056,In_1001,In_141);
and U1057 (N_1057,In_375,In_1371);
nor U1058 (N_1058,In_1207,In_349);
and U1059 (N_1059,In_1084,In_788);
and U1060 (N_1060,In_707,In_548);
or U1061 (N_1061,In_478,In_1199);
nor U1062 (N_1062,In_457,In_1148);
or U1063 (N_1063,In_745,In_900);
xor U1064 (N_1064,In_1293,In_505);
or U1065 (N_1065,In_1207,In_1189);
or U1066 (N_1066,In_584,In_880);
xor U1067 (N_1067,In_167,In_642);
and U1068 (N_1068,In_1179,In_960);
nor U1069 (N_1069,In_233,In_118);
nor U1070 (N_1070,In_215,In_1119);
nor U1071 (N_1071,In_916,In_871);
nand U1072 (N_1072,In_1477,In_1332);
or U1073 (N_1073,In_408,In_352);
or U1074 (N_1074,In_933,In_282);
or U1075 (N_1075,In_1067,In_1064);
or U1076 (N_1076,In_15,In_80);
xor U1077 (N_1077,In_1122,In_22);
nor U1078 (N_1078,In_613,In_56);
nor U1079 (N_1079,In_523,In_50);
or U1080 (N_1080,In_723,In_1147);
or U1081 (N_1081,In_105,In_1351);
nand U1082 (N_1082,In_49,In_396);
nor U1083 (N_1083,In_576,In_568);
nor U1084 (N_1084,In_400,In_818);
or U1085 (N_1085,In_1369,In_1052);
or U1086 (N_1086,In_250,In_88);
nor U1087 (N_1087,In_211,In_1138);
nand U1088 (N_1088,In_425,In_1251);
nand U1089 (N_1089,In_580,In_538);
xnor U1090 (N_1090,In_90,In_696);
nand U1091 (N_1091,In_672,In_1474);
or U1092 (N_1092,In_407,In_1356);
nor U1093 (N_1093,In_673,In_1012);
nand U1094 (N_1094,In_339,In_31);
nand U1095 (N_1095,In_337,In_1258);
and U1096 (N_1096,In_865,In_671);
nor U1097 (N_1097,In_504,In_217);
xor U1098 (N_1098,In_143,In_649);
and U1099 (N_1099,In_496,In_1108);
nand U1100 (N_1100,In_227,In_577);
or U1101 (N_1101,In_609,In_593);
or U1102 (N_1102,In_832,In_931);
or U1103 (N_1103,In_1157,In_334);
and U1104 (N_1104,In_183,In_465);
nand U1105 (N_1105,In_1049,In_55);
nor U1106 (N_1106,In_178,In_787);
nor U1107 (N_1107,In_659,In_32);
nand U1108 (N_1108,In_287,In_700);
nand U1109 (N_1109,In_981,In_112);
or U1110 (N_1110,In_1451,In_1250);
nand U1111 (N_1111,In_1383,In_594);
nand U1112 (N_1112,In_976,In_999);
and U1113 (N_1113,In_954,In_308);
nor U1114 (N_1114,In_336,In_315);
xor U1115 (N_1115,In_718,In_458);
and U1116 (N_1116,In_369,In_1005);
and U1117 (N_1117,In_460,In_1288);
xor U1118 (N_1118,In_1012,In_404);
nand U1119 (N_1119,In_988,In_884);
nand U1120 (N_1120,In_684,In_1142);
or U1121 (N_1121,In_894,In_1061);
and U1122 (N_1122,In_1096,In_272);
nand U1123 (N_1123,In_1271,In_1364);
nand U1124 (N_1124,In_367,In_1443);
nand U1125 (N_1125,In_844,In_390);
nand U1126 (N_1126,In_428,In_587);
nand U1127 (N_1127,In_580,In_21);
and U1128 (N_1128,In_538,In_396);
nor U1129 (N_1129,In_187,In_1254);
or U1130 (N_1130,In_605,In_795);
nor U1131 (N_1131,In_1275,In_1072);
or U1132 (N_1132,In_830,In_586);
and U1133 (N_1133,In_1241,In_902);
or U1134 (N_1134,In_1065,In_562);
and U1135 (N_1135,In_582,In_1209);
nand U1136 (N_1136,In_431,In_903);
nand U1137 (N_1137,In_1464,In_119);
or U1138 (N_1138,In_100,In_1014);
nand U1139 (N_1139,In_1434,In_311);
nand U1140 (N_1140,In_893,In_606);
nor U1141 (N_1141,In_345,In_113);
or U1142 (N_1142,In_1496,In_281);
or U1143 (N_1143,In_977,In_245);
nand U1144 (N_1144,In_405,In_810);
nand U1145 (N_1145,In_483,In_931);
or U1146 (N_1146,In_427,In_906);
and U1147 (N_1147,In_434,In_317);
and U1148 (N_1148,In_660,In_783);
or U1149 (N_1149,In_18,In_828);
nor U1150 (N_1150,In_578,In_1137);
and U1151 (N_1151,In_1021,In_1403);
nand U1152 (N_1152,In_700,In_516);
nand U1153 (N_1153,In_839,In_971);
or U1154 (N_1154,In_1019,In_1300);
and U1155 (N_1155,In_778,In_279);
nor U1156 (N_1156,In_133,In_426);
nand U1157 (N_1157,In_656,In_118);
xnor U1158 (N_1158,In_203,In_798);
nor U1159 (N_1159,In_1496,In_214);
nand U1160 (N_1160,In_785,In_644);
nor U1161 (N_1161,In_785,In_620);
nand U1162 (N_1162,In_1026,In_717);
and U1163 (N_1163,In_18,In_636);
nor U1164 (N_1164,In_1065,In_450);
nor U1165 (N_1165,In_502,In_1380);
and U1166 (N_1166,In_895,In_891);
nand U1167 (N_1167,In_1279,In_666);
nor U1168 (N_1168,In_811,In_1330);
or U1169 (N_1169,In_323,In_1426);
and U1170 (N_1170,In_107,In_777);
or U1171 (N_1171,In_1078,In_33);
nand U1172 (N_1172,In_1125,In_1480);
nand U1173 (N_1173,In_326,In_115);
or U1174 (N_1174,In_300,In_495);
or U1175 (N_1175,In_800,In_1077);
xor U1176 (N_1176,In_1227,In_556);
nand U1177 (N_1177,In_928,In_803);
and U1178 (N_1178,In_182,In_834);
nor U1179 (N_1179,In_1450,In_117);
or U1180 (N_1180,In_773,In_620);
or U1181 (N_1181,In_638,In_18);
nand U1182 (N_1182,In_1069,In_313);
nand U1183 (N_1183,In_41,In_721);
xor U1184 (N_1184,In_52,In_287);
nor U1185 (N_1185,In_871,In_1264);
and U1186 (N_1186,In_1149,In_712);
nor U1187 (N_1187,In_137,In_256);
or U1188 (N_1188,In_1393,In_219);
or U1189 (N_1189,In_1430,In_1108);
nor U1190 (N_1190,In_1382,In_684);
or U1191 (N_1191,In_1162,In_1103);
xnor U1192 (N_1192,In_523,In_1035);
xor U1193 (N_1193,In_719,In_886);
and U1194 (N_1194,In_412,In_481);
or U1195 (N_1195,In_848,In_668);
or U1196 (N_1196,In_996,In_405);
and U1197 (N_1197,In_484,In_102);
and U1198 (N_1198,In_1283,In_1115);
and U1199 (N_1199,In_242,In_702);
or U1200 (N_1200,In_1304,In_1164);
and U1201 (N_1201,In_705,In_1107);
nor U1202 (N_1202,In_1235,In_123);
nor U1203 (N_1203,In_757,In_264);
nand U1204 (N_1204,In_855,In_919);
and U1205 (N_1205,In_1190,In_116);
and U1206 (N_1206,In_1134,In_869);
or U1207 (N_1207,In_545,In_145);
xor U1208 (N_1208,In_397,In_115);
nor U1209 (N_1209,In_398,In_462);
nand U1210 (N_1210,In_1498,In_872);
and U1211 (N_1211,In_1073,In_1359);
and U1212 (N_1212,In_144,In_714);
or U1213 (N_1213,In_726,In_1471);
nand U1214 (N_1214,In_68,In_611);
nor U1215 (N_1215,In_1153,In_895);
or U1216 (N_1216,In_541,In_1036);
xnor U1217 (N_1217,In_1315,In_1495);
nor U1218 (N_1218,In_1337,In_1140);
nand U1219 (N_1219,In_107,In_1351);
and U1220 (N_1220,In_566,In_1079);
or U1221 (N_1221,In_345,In_682);
nor U1222 (N_1222,In_386,In_586);
or U1223 (N_1223,In_738,In_642);
nand U1224 (N_1224,In_1427,In_1434);
or U1225 (N_1225,In_1139,In_664);
and U1226 (N_1226,In_256,In_807);
or U1227 (N_1227,In_602,In_693);
xor U1228 (N_1228,In_192,In_359);
and U1229 (N_1229,In_12,In_855);
or U1230 (N_1230,In_585,In_333);
xor U1231 (N_1231,In_1348,In_1140);
nor U1232 (N_1232,In_887,In_1172);
and U1233 (N_1233,In_472,In_1365);
or U1234 (N_1234,In_1076,In_1328);
nand U1235 (N_1235,In_790,In_816);
or U1236 (N_1236,In_333,In_1201);
nand U1237 (N_1237,In_470,In_289);
or U1238 (N_1238,In_1115,In_602);
nand U1239 (N_1239,In_545,In_1058);
and U1240 (N_1240,In_35,In_1337);
and U1241 (N_1241,In_723,In_1176);
xnor U1242 (N_1242,In_641,In_406);
nand U1243 (N_1243,In_1486,In_329);
and U1244 (N_1244,In_96,In_556);
xor U1245 (N_1245,In_1294,In_1220);
nor U1246 (N_1246,In_114,In_1264);
nand U1247 (N_1247,In_126,In_1055);
nor U1248 (N_1248,In_375,In_279);
or U1249 (N_1249,In_166,In_1368);
nor U1250 (N_1250,In_202,In_661);
nand U1251 (N_1251,In_195,In_855);
nand U1252 (N_1252,In_746,In_979);
and U1253 (N_1253,In_365,In_1407);
xnor U1254 (N_1254,In_1484,In_1047);
nor U1255 (N_1255,In_1325,In_688);
nor U1256 (N_1256,In_1135,In_1260);
nor U1257 (N_1257,In_136,In_653);
nand U1258 (N_1258,In_1261,In_237);
and U1259 (N_1259,In_1102,In_1093);
nand U1260 (N_1260,In_12,In_664);
or U1261 (N_1261,In_223,In_856);
nor U1262 (N_1262,In_238,In_1216);
nand U1263 (N_1263,In_923,In_1341);
or U1264 (N_1264,In_832,In_122);
or U1265 (N_1265,In_1088,In_793);
nand U1266 (N_1266,In_764,In_474);
nand U1267 (N_1267,In_862,In_880);
nand U1268 (N_1268,In_685,In_274);
nor U1269 (N_1269,In_1249,In_105);
and U1270 (N_1270,In_988,In_1394);
nand U1271 (N_1271,In_207,In_276);
and U1272 (N_1272,In_391,In_35);
nor U1273 (N_1273,In_1154,In_1116);
or U1274 (N_1274,In_657,In_415);
or U1275 (N_1275,In_1229,In_75);
or U1276 (N_1276,In_737,In_491);
or U1277 (N_1277,In_876,In_384);
nand U1278 (N_1278,In_976,In_996);
nand U1279 (N_1279,In_958,In_252);
nand U1280 (N_1280,In_115,In_1380);
or U1281 (N_1281,In_631,In_884);
nor U1282 (N_1282,In_1191,In_446);
nor U1283 (N_1283,In_808,In_333);
xnor U1284 (N_1284,In_970,In_665);
nand U1285 (N_1285,In_1191,In_1447);
nand U1286 (N_1286,In_353,In_387);
nor U1287 (N_1287,In_1064,In_1303);
and U1288 (N_1288,In_1022,In_126);
nor U1289 (N_1289,In_1379,In_955);
nand U1290 (N_1290,In_858,In_1396);
nor U1291 (N_1291,In_1356,In_1105);
nand U1292 (N_1292,In_1370,In_481);
and U1293 (N_1293,In_8,In_1474);
nor U1294 (N_1294,In_1274,In_335);
and U1295 (N_1295,In_97,In_716);
and U1296 (N_1296,In_421,In_222);
xor U1297 (N_1297,In_820,In_910);
or U1298 (N_1298,In_1477,In_1098);
and U1299 (N_1299,In_1051,In_719);
or U1300 (N_1300,In_59,In_66);
or U1301 (N_1301,In_266,In_375);
nand U1302 (N_1302,In_189,In_601);
nor U1303 (N_1303,In_133,In_284);
nor U1304 (N_1304,In_666,In_1258);
nand U1305 (N_1305,In_334,In_1055);
nand U1306 (N_1306,In_133,In_564);
nor U1307 (N_1307,In_1228,In_1303);
nand U1308 (N_1308,In_1005,In_1418);
nand U1309 (N_1309,In_387,In_1408);
nor U1310 (N_1310,In_837,In_497);
nor U1311 (N_1311,In_1128,In_900);
and U1312 (N_1312,In_1402,In_1267);
nand U1313 (N_1313,In_1318,In_865);
and U1314 (N_1314,In_779,In_7);
nand U1315 (N_1315,In_612,In_1301);
and U1316 (N_1316,In_499,In_746);
nor U1317 (N_1317,In_4,In_1365);
nor U1318 (N_1318,In_721,In_746);
nor U1319 (N_1319,In_597,In_32);
or U1320 (N_1320,In_1214,In_803);
xnor U1321 (N_1321,In_1304,In_291);
or U1322 (N_1322,In_1013,In_1272);
xor U1323 (N_1323,In_52,In_1296);
and U1324 (N_1324,In_813,In_545);
or U1325 (N_1325,In_323,In_173);
and U1326 (N_1326,In_635,In_350);
nor U1327 (N_1327,In_647,In_714);
or U1328 (N_1328,In_1108,In_485);
and U1329 (N_1329,In_255,In_176);
and U1330 (N_1330,In_1430,In_1309);
or U1331 (N_1331,In_813,In_1461);
nor U1332 (N_1332,In_1350,In_644);
or U1333 (N_1333,In_787,In_407);
or U1334 (N_1334,In_221,In_1272);
or U1335 (N_1335,In_1427,In_1248);
xor U1336 (N_1336,In_104,In_1447);
nand U1337 (N_1337,In_642,In_778);
and U1338 (N_1338,In_733,In_505);
or U1339 (N_1339,In_880,In_824);
and U1340 (N_1340,In_886,In_1294);
and U1341 (N_1341,In_48,In_1070);
nor U1342 (N_1342,In_848,In_1271);
nor U1343 (N_1343,In_1343,In_1291);
or U1344 (N_1344,In_244,In_1396);
nor U1345 (N_1345,In_21,In_1168);
nor U1346 (N_1346,In_340,In_417);
or U1347 (N_1347,In_1470,In_153);
nor U1348 (N_1348,In_1252,In_1231);
nor U1349 (N_1349,In_453,In_1178);
nor U1350 (N_1350,In_315,In_1307);
and U1351 (N_1351,In_229,In_1204);
xor U1352 (N_1352,In_1362,In_499);
or U1353 (N_1353,In_290,In_1389);
nor U1354 (N_1354,In_936,In_796);
nand U1355 (N_1355,In_359,In_900);
xor U1356 (N_1356,In_159,In_1196);
nor U1357 (N_1357,In_949,In_1386);
nand U1358 (N_1358,In_6,In_1347);
and U1359 (N_1359,In_200,In_281);
and U1360 (N_1360,In_280,In_383);
and U1361 (N_1361,In_828,In_1425);
or U1362 (N_1362,In_163,In_124);
and U1363 (N_1363,In_145,In_469);
and U1364 (N_1364,In_633,In_709);
or U1365 (N_1365,In_1142,In_429);
and U1366 (N_1366,In_224,In_91);
nor U1367 (N_1367,In_586,In_437);
nand U1368 (N_1368,In_765,In_680);
nand U1369 (N_1369,In_1473,In_1480);
nor U1370 (N_1370,In_347,In_1359);
nand U1371 (N_1371,In_895,In_415);
or U1372 (N_1372,In_1255,In_66);
nor U1373 (N_1373,In_869,In_966);
nor U1374 (N_1374,In_834,In_201);
and U1375 (N_1375,In_257,In_447);
xor U1376 (N_1376,In_975,In_302);
nor U1377 (N_1377,In_634,In_616);
or U1378 (N_1378,In_859,In_1277);
and U1379 (N_1379,In_140,In_114);
and U1380 (N_1380,In_980,In_199);
and U1381 (N_1381,In_362,In_1017);
nor U1382 (N_1382,In_252,In_477);
and U1383 (N_1383,In_899,In_1305);
nor U1384 (N_1384,In_762,In_125);
and U1385 (N_1385,In_611,In_140);
or U1386 (N_1386,In_154,In_262);
nand U1387 (N_1387,In_131,In_555);
nor U1388 (N_1388,In_1184,In_1438);
or U1389 (N_1389,In_1384,In_701);
nor U1390 (N_1390,In_940,In_1062);
or U1391 (N_1391,In_1249,In_97);
nand U1392 (N_1392,In_1160,In_883);
and U1393 (N_1393,In_162,In_235);
and U1394 (N_1394,In_718,In_1466);
nand U1395 (N_1395,In_145,In_439);
nor U1396 (N_1396,In_664,In_557);
or U1397 (N_1397,In_664,In_967);
and U1398 (N_1398,In_765,In_1425);
nand U1399 (N_1399,In_1102,In_298);
or U1400 (N_1400,In_1401,In_872);
nand U1401 (N_1401,In_213,In_115);
or U1402 (N_1402,In_1097,In_585);
xnor U1403 (N_1403,In_84,In_478);
nor U1404 (N_1404,In_80,In_1118);
xnor U1405 (N_1405,In_574,In_1018);
or U1406 (N_1406,In_208,In_152);
nor U1407 (N_1407,In_276,In_509);
and U1408 (N_1408,In_402,In_1103);
nor U1409 (N_1409,In_142,In_1122);
nor U1410 (N_1410,In_1475,In_572);
xnor U1411 (N_1411,In_1074,In_691);
or U1412 (N_1412,In_1077,In_264);
nor U1413 (N_1413,In_937,In_691);
nand U1414 (N_1414,In_1123,In_95);
and U1415 (N_1415,In_438,In_1259);
and U1416 (N_1416,In_671,In_1387);
or U1417 (N_1417,In_275,In_1141);
and U1418 (N_1418,In_814,In_797);
nor U1419 (N_1419,In_615,In_1150);
nand U1420 (N_1420,In_1057,In_1110);
nor U1421 (N_1421,In_1171,In_167);
nor U1422 (N_1422,In_1292,In_1418);
nor U1423 (N_1423,In_819,In_207);
nand U1424 (N_1424,In_93,In_952);
nor U1425 (N_1425,In_537,In_1013);
and U1426 (N_1426,In_284,In_514);
nor U1427 (N_1427,In_744,In_918);
or U1428 (N_1428,In_993,In_1429);
and U1429 (N_1429,In_1189,In_477);
nor U1430 (N_1430,In_429,In_683);
or U1431 (N_1431,In_1079,In_633);
and U1432 (N_1432,In_313,In_696);
nor U1433 (N_1433,In_1257,In_752);
or U1434 (N_1434,In_1231,In_932);
nand U1435 (N_1435,In_359,In_588);
nor U1436 (N_1436,In_881,In_694);
and U1437 (N_1437,In_1385,In_110);
nand U1438 (N_1438,In_471,In_3);
nand U1439 (N_1439,In_486,In_1065);
and U1440 (N_1440,In_1382,In_208);
nor U1441 (N_1441,In_436,In_727);
nand U1442 (N_1442,In_686,In_1182);
xor U1443 (N_1443,In_1002,In_1271);
and U1444 (N_1444,In_441,In_751);
nor U1445 (N_1445,In_1346,In_207);
and U1446 (N_1446,In_582,In_826);
and U1447 (N_1447,In_474,In_303);
nand U1448 (N_1448,In_966,In_1329);
nand U1449 (N_1449,In_1398,In_959);
nor U1450 (N_1450,In_521,In_674);
and U1451 (N_1451,In_401,In_1056);
nand U1452 (N_1452,In_461,In_601);
nor U1453 (N_1453,In_223,In_467);
nand U1454 (N_1454,In_684,In_655);
nor U1455 (N_1455,In_77,In_1261);
or U1456 (N_1456,In_1214,In_509);
nand U1457 (N_1457,In_1181,In_15);
or U1458 (N_1458,In_1063,In_973);
nor U1459 (N_1459,In_221,In_189);
nor U1460 (N_1460,In_358,In_1323);
nand U1461 (N_1461,In_758,In_32);
nand U1462 (N_1462,In_1109,In_378);
or U1463 (N_1463,In_403,In_1258);
nand U1464 (N_1464,In_1280,In_288);
nor U1465 (N_1465,In_934,In_512);
nor U1466 (N_1466,In_628,In_1374);
and U1467 (N_1467,In_1192,In_100);
or U1468 (N_1468,In_461,In_136);
and U1469 (N_1469,In_1241,In_1094);
or U1470 (N_1470,In_133,In_1368);
nand U1471 (N_1471,In_903,In_194);
and U1472 (N_1472,In_1128,In_1021);
nand U1473 (N_1473,In_89,In_118);
and U1474 (N_1474,In_1000,In_719);
nand U1475 (N_1475,In_180,In_1444);
or U1476 (N_1476,In_1097,In_50);
nor U1477 (N_1477,In_1228,In_52);
or U1478 (N_1478,In_3,In_653);
and U1479 (N_1479,In_721,In_1231);
nand U1480 (N_1480,In_663,In_755);
nor U1481 (N_1481,In_714,In_495);
nor U1482 (N_1482,In_1213,In_1046);
xor U1483 (N_1483,In_883,In_678);
xor U1484 (N_1484,In_561,In_967);
nor U1485 (N_1485,In_1157,In_490);
or U1486 (N_1486,In_517,In_585);
or U1487 (N_1487,In_1397,In_293);
and U1488 (N_1488,In_651,In_816);
nor U1489 (N_1489,In_1136,In_673);
and U1490 (N_1490,In_976,In_797);
or U1491 (N_1491,In_1255,In_957);
and U1492 (N_1492,In_650,In_474);
nand U1493 (N_1493,In_1369,In_843);
xnor U1494 (N_1494,In_1183,In_1051);
nand U1495 (N_1495,In_350,In_750);
nor U1496 (N_1496,In_399,In_855);
xnor U1497 (N_1497,In_587,In_696);
nand U1498 (N_1498,In_631,In_1241);
nor U1499 (N_1499,In_17,In_559);
nand U1500 (N_1500,N_853,N_652);
nand U1501 (N_1501,N_910,N_383);
xnor U1502 (N_1502,N_366,N_1494);
nand U1503 (N_1503,N_179,N_1408);
and U1504 (N_1504,N_1386,N_1156);
nor U1505 (N_1505,N_350,N_997);
nand U1506 (N_1506,N_1285,N_646);
nor U1507 (N_1507,N_712,N_1341);
and U1508 (N_1508,N_500,N_268);
or U1509 (N_1509,N_390,N_1005);
and U1510 (N_1510,N_17,N_126);
or U1511 (N_1511,N_94,N_358);
and U1512 (N_1512,N_679,N_284);
nor U1513 (N_1513,N_1446,N_983);
xor U1514 (N_1514,N_989,N_305);
nand U1515 (N_1515,N_36,N_1233);
nor U1516 (N_1516,N_556,N_831);
nand U1517 (N_1517,N_525,N_589);
or U1518 (N_1518,N_1464,N_1270);
nor U1519 (N_1519,N_52,N_637);
nand U1520 (N_1520,N_357,N_484);
and U1521 (N_1521,N_76,N_406);
nand U1522 (N_1522,N_335,N_1470);
and U1523 (N_1523,N_842,N_422);
and U1524 (N_1524,N_1375,N_794);
nand U1525 (N_1525,N_253,N_63);
nand U1526 (N_1526,N_766,N_1373);
nor U1527 (N_1527,N_982,N_1283);
nand U1528 (N_1528,N_323,N_1287);
or U1529 (N_1529,N_854,N_631);
nor U1530 (N_1530,N_746,N_1184);
and U1531 (N_1531,N_685,N_310);
or U1532 (N_1532,N_1453,N_561);
and U1533 (N_1533,N_1317,N_784);
nor U1534 (N_1534,N_1152,N_18);
or U1535 (N_1535,N_1170,N_509);
nand U1536 (N_1536,N_1249,N_998);
nor U1537 (N_1537,N_662,N_1312);
nand U1538 (N_1538,N_674,N_707);
or U1539 (N_1539,N_1062,N_1151);
nand U1540 (N_1540,N_461,N_936);
or U1541 (N_1541,N_93,N_1467);
and U1542 (N_1542,N_583,N_340);
nand U1543 (N_1543,N_687,N_45);
or U1544 (N_1544,N_1463,N_499);
xnor U1545 (N_1545,N_751,N_105);
and U1546 (N_1546,N_302,N_324);
and U1547 (N_1547,N_981,N_57);
nand U1548 (N_1548,N_557,N_1058);
nand U1549 (N_1549,N_949,N_1024);
nand U1550 (N_1550,N_153,N_1242);
or U1551 (N_1551,N_404,N_287);
nand U1552 (N_1552,N_378,N_41);
or U1553 (N_1553,N_480,N_1206);
nand U1554 (N_1554,N_1426,N_1038);
nor U1555 (N_1555,N_431,N_527);
nand U1556 (N_1556,N_196,N_1411);
or U1557 (N_1557,N_344,N_1085);
or U1558 (N_1558,N_772,N_992);
nand U1559 (N_1559,N_584,N_329);
nand U1560 (N_1560,N_919,N_1288);
or U1561 (N_1561,N_782,N_1339);
or U1562 (N_1562,N_1313,N_1271);
and U1563 (N_1563,N_501,N_1168);
and U1564 (N_1564,N_701,N_569);
and U1565 (N_1565,N_192,N_942);
nor U1566 (N_1566,N_748,N_13);
nand U1567 (N_1567,N_606,N_1350);
nor U1568 (N_1568,N_724,N_675);
nand U1569 (N_1569,N_803,N_1396);
nand U1570 (N_1570,N_16,N_623);
nand U1571 (N_1571,N_6,N_25);
nor U1572 (N_1572,N_504,N_1105);
nor U1573 (N_1573,N_700,N_219);
nor U1574 (N_1574,N_514,N_103);
nor U1575 (N_1575,N_551,N_211);
nand U1576 (N_1576,N_950,N_974);
or U1577 (N_1577,N_1070,N_777);
nor U1578 (N_1578,N_75,N_475);
or U1579 (N_1579,N_190,N_1109);
and U1580 (N_1580,N_279,N_1003);
nor U1581 (N_1581,N_764,N_1043);
nor U1582 (N_1582,N_1089,N_448);
xnor U1583 (N_1583,N_194,N_574);
nor U1584 (N_1584,N_1268,N_1051);
xor U1585 (N_1585,N_1099,N_1000);
and U1586 (N_1586,N_800,N_108);
and U1587 (N_1587,N_388,N_1358);
nand U1588 (N_1588,N_188,N_1418);
nor U1589 (N_1589,N_1338,N_1110);
nor U1590 (N_1590,N_879,N_1247);
and U1591 (N_1591,N_314,N_1141);
and U1592 (N_1592,N_166,N_1262);
nor U1593 (N_1593,N_161,N_1333);
xor U1594 (N_1594,N_655,N_1314);
nand U1595 (N_1595,N_601,N_1286);
nand U1596 (N_1596,N_596,N_487);
and U1597 (N_1597,N_498,N_222);
nand U1598 (N_1598,N_787,N_537);
or U1599 (N_1599,N_934,N_49);
nor U1600 (N_1600,N_79,N_859);
nor U1601 (N_1601,N_672,N_418);
nor U1602 (N_1602,N_621,N_814);
nand U1603 (N_1603,N_1423,N_670);
nor U1604 (N_1604,N_1441,N_410);
xnor U1605 (N_1605,N_1295,N_1325);
or U1606 (N_1606,N_1497,N_58);
nand U1607 (N_1607,N_96,N_432);
nand U1608 (N_1608,N_2,N_1328);
or U1609 (N_1609,N_916,N_603);
or U1610 (N_1610,N_1033,N_534);
xnor U1611 (N_1611,N_463,N_334);
or U1612 (N_1612,N_636,N_812);
or U1613 (N_1613,N_191,N_201);
nand U1614 (N_1614,N_1366,N_1476);
or U1615 (N_1615,N_1133,N_586);
nor U1616 (N_1616,N_1034,N_1297);
and U1617 (N_1617,N_688,N_411);
nand U1618 (N_1618,N_35,N_817);
and U1619 (N_1619,N_1017,N_593);
or U1620 (N_1620,N_907,N_1150);
nand U1621 (N_1621,N_1444,N_107);
nor U1622 (N_1622,N_237,N_479);
and U1623 (N_1623,N_138,N_1129);
and U1624 (N_1624,N_1007,N_200);
or U1625 (N_1625,N_1395,N_884);
or U1626 (N_1626,N_808,N_1304);
or U1627 (N_1627,N_1445,N_752);
nand U1628 (N_1628,N_78,N_1102);
and U1629 (N_1629,N_506,N_767);
nand U1630 (N_1630,N_795,N_619);
and U1631 (N_1631,N_239,N_540);
and U1632 (N_1632,N_1347,N_451);
nor U1633 (N_1633,N_924,N_649);
nor U1634 (N_1634,N_644,N_186);
nand U1635 (N_1635,N_1210,N_1404);
nand U1636 (N_1636,N_294,N_880);
and U1637 (N_1637,N_1094,N_640);
nor U1638 (N_1638,N_909,N_715);
nand U1639 (N_1639,N_882,N_154);
or U1640 (N_1640,N_897,N_810);
and U1641 (N_1641,N_783,N_469);
nand U1642 (N_1642,N_277,N_667);
nand U1643 (N_1643,N_1468,N_532);
nand U1644 (N_1644,N_172,N_1037);
and U1645 (N_1645,N_682,N_592);
nor U1646 (N_1646,N_1278,N_825);
nand U1647 (N_1647,N_1485,N_734);
nand U1648 (N_1648,N_677,N_454);
nand U1649 (N_1649,N_155,N_316);
or U1650 (N_1650,N_804,N_1010);
xor U1651 (N_1651,N_261,N_1267);
nor U1652 (N_1652,N_81,N_1498);
nand U1653 (N_1653,N_394,N_131);
or U1654 (N_1654,N_470,N_1213);
and U1655 (N_1655,N_1360,N_89);
and U1656 (N_1656,N_1078,N_1425);
nand U1657 (N_1657,N_124,N_379);
nor U1658 (N_1658,N_526,N_1415);
or U1659 (N_1659,N_477,N_260);
xor U1660 (N_1660,N_262,N_1290);
or U1661 (N_1661,N_208,N_564);
nand U1662 (N_1662,N_732,N_903);
nor U1663 (N_1663,N_252,N_474);
or U1664 (N_1664,N_1348,N_71);
nand U1665 (N_1665,N_729,N_642);
and U1666 (N_1666,N_587,N_369);
nand U1667 (N_1667,N_1088,N_1071);
xnor U1668 (N_1668,N_40,N_1186);
nand U1669 (N_1669,N_42,N_12);
xnor U1670 (N_1670,N_877,N_915);
or U1671 (N_1671,N_923,N_64);
or U1672 (N_1672,N_645,N_1394);
and U1673 (N_1673,N_607,N_444);
or U1674 (N_1674,N_1238,N_1457);
and U1675 (N_1675,N_616,N_553);
nand U1676 (N_1676,N_790,N_1119);
nand U1677 (N_1677,N_1368,N_355);
nand U1678 (N_1678,N_1044,N_1443);
nand U1679 (N_1679,N_1157,N_960);
or U1680 (N_1680,N_1009,N_288);
nor U1681 (N_1681,N_549,N_872);
nor U1682 (N_1682,N_22,N_1334);
nor U1683 (N_1683,N_1020,N_398);
nand U1684 (N_1684,N_176,N_898);
nor U1685 (N_1685,N_478,N_168);
nand U1686 (N_1686,N_46,N_317);
and U1687 (N_1687,N_11,N_1202);
and U1688 (N_1688,N_72,N_414);
nand U1689 (N_1689,N_683,N_691);
or U1690 (N_1690,N_1039,N_273);
nand U1691 (N_1691,N_1371,N_405);
nand U1692 (N_1692,N_1264,N_867);
or U1693 (N_1693,N_32,N_1201);
and U1694 (N_1694,N_906,N_1194);
nand U1695 (N_1695,N_212,N_571);
or U1696 (N_1696,N_612,N_720);
or U1697 (N_1697,N_7,N_993);
nor U1698 (N_1698,N_833,N_956);
nand U1699 (N_1699,N_87,N_1257);
nor U1700 (N_1700,N_890,N_1482);
nor U1701 (N_1701,N_259,N_468);
nor U1702 (N_1702,N_146,N_1231);
nand U1703 (N_1703,N_535,N_1065);
or U1704 (N_1704,N_615,N_427);
or U1705 (N_1705,N_604,N_581);
nand U1706 (N_1706,N_522,N_1075);
or U1707 (N_1707,N_929,N_727);
nand U1708 (N_1708,N_778,N_733);
nor U1709 (N_1709,N_100,N_696);
nand U1710 (N_1710,N_330,N_488);
nor U1711 (N_1711,N_312,N_97);
nor U1712 (N_1712,N_135,N_351);
and U1713 (N_1713,N_1123,N_1298);
nor U1714 (N_1714,N_95,N_241);
nor U1715 (N_1715,N_1057,N_958);
nand U1716 (N_1716,N_940,N_1319);
xor U1717 (N_1717,N_231,N_823);
and U1718 (N_1718,N_1148,N_1310);
xor U1719 (N_1719,N_1438,N_546);
nor U1720 (N_1720,N_1493,N_676);
nand U1721 (N_1721,N_141,N_954);
xnor U1722 (N_1722,N_321,N_492);
nor U1723 (N_1723,N_336,N_1437);
nor U1724 (N_1724,N_913,N_1336);
and U1725 (N_1725,N_1180,N_348);
and U1726 (N_1726,N_1155,N_1200);
xor U1727 (N_1727,N_523,N_1289);
nand U1728 (N_1728,N_695,N_1128);
nand U1729 (N_1729,N_507,N_442);
or U1730 (N_1730,N_705,N_1045);
and U1731 (N_1731,N_888,N_1211);
nand U1732 (N_1732,N_918,N_1393);
nor U1733 (N_1733,N_1047,N_311);
or U1734 (N_1734,N_1196,N_1234);
or U1735 (N_1735,N_1054,N_1093);
or U1736 (N_1736,N_403,N_1377);
or U1737 (N_1737,N_1309,N_223);
xnor U1738 (N_1738,N_570,N_1203);
and U1739 (N_1739,N_548,N_1473);
or U1740 (N_1740,N_495,N_893);
and U1741 (N_1741,N_743,N_757);
nor U1742 (N_1742,N_159,N_216);
or U1743 (N_1743,N_1436,N_1417);
nor U1744 (N_1744,N_1145,N_1299);
and U1745 (N_1745,N_56,N_684);
or U1746 (N_1746,N_1307,N_263);
or U1747 (N_1747,N_1232,N_663);
or U1748 (N_1748,N_973,N_598);
nor U1749 (N_1749,N_568,N_741);
and U1750 (N_1750,N_1471,N_524);
nor U1751 (N_1751,N_1452,N_789);
or U1752 (N_1752,N_567,N_1204);
nor U1753 (N_1753,N_892,N_445);
nand U1754 (N_1754,N_515,N_953);
xnor U1755 (N_1755,N_293,N_31);
nor U1756 (N_1756,N_1191,N_1013);
nor U1757 (N_1757,N_19,N_425);
nor U1758 (N_1758,N_372,N_401);
xor U1759 (N_1759,N_512,N_681);
nor U1760 (N_1760,N_1219,N_744);
or U1761 (N_1761,N_1107,N_780);
or U1762 (N_1762,N_271,N_1385);
xor U1763 (N_1763,N_98,N_1014);
nor U1764 (N_1764,N_133,N_1069);
or U1765 (N_1765,N_1035,N_1272);
nand U1766 (N_1766,N_354,N_1134);
and U1767 (N_1767,N_1274,N_38);
or U1768 (N_1768,N_559,N_985);
and U1769 (N_1769,N_362,N_453);
nand U1770 (N_1770,N_249,N_1087);
nor U1771 (N_1771,N_1082,N_69);
or U1772 (N_1772,N_728,N_65);
xnor U1773 (N_1773,N_112,N_1161);
and U1774 (N_1774,N_1029,N_420);
nor U1775 (N_1775,N_761,N_1303);
and U1776 (N_1776,N_828,N_709);
xor U1777 (N_1777,N_24,N_862);
nor U1778 (N_1778,N_242,N_1064);
nand U1779 (N_1779,N_286,N_742);
or U1780 (N_1780,N_333,N_827);
or U1781 (N_1781,N_143,N_1177);
nand U1782 (N_1782,N_338,N_1120);
and U1783 (N_1783,N_434,N_55);
nor U1784 (N_1784,N_303,N_1337);
nand U1785 (N_1785,N_449,N_554);
nor U1786 (N_1786,N_489,N_628);
nand U1787 (N_1787,N_821,N_1430);
or U1788 (N_1788,N_197,N_1451);
nor U1789 (N_1789,N_624,N_1046);
nand U1790 (N_1790,N_326,N_666);
nor U1791 (N_1791,N_1012,N_1023);
and U1792 (N_1792,N_210,N_1390);
nand U1793 (N_1793,N_835,N_1052);
nand U1794 (N_1794,N_1098,N_137);
nor U1795 (N_1795,N_174,N_182);
nor U1796 (N_1796,N_60,N_891);
xnor U1797 (N_1797,N_639,N_1146);
nor U1798 (N_1798,N_1127,N_660);
and U1799 (N_1799,N_868,N_673);
nand U1800 (N_1800,N_1015,N_1032);
or U1801 (N_1801,N_1248,N_796);
or U1802 (N_1802,N_1488,N_984);
or U1803 (N_1803,N_387,N_632);
nand U1804 (N_1804,N_1136,N_295);
or U1805 (N_1805,N_1228,N_1217);
or U1806 (N_1806,N_1412,N_1409);
nor U1807 (N_1807,N_585,N_446);
and U1808 (N_1808,N_23,N_84);
or U1809 (N_1809,N_1113,N_125);
nand U1810 (N_1810,N_622,N_80);
or U1811 (N_1811,N_1369,N_306);
xnor U1812 (N_1812,N_1022,N_162);
and U1813 (N_1813,N_1226,N_145);
nand U1814 (N_1814,N_37,N_1469);
or U1815 (N_1815,N_441,N_502);
xnor U1816 (N_1816,N_1080,N_101);
nand U1817 (N_1817,N_352,N_713);
xnor U1818 (N_1818,N_832,N_1086);
xnor U1819 (N_1819,N_1439,N_920);
nor U1820 (N_1820,N_735,N_873);
nor U1821 (N_1821,N_205,N_493);
nand U1822 (N_1822,N_1096,N_356);
and U1823 (N_1823,N_409,N_952);
nor U1824 (N_1824,N_830,N_1164);
or U1825 (N_1825,N_206,N_834);
or U1826 (N_1826,N_904,N_1079);
nor U1827 (N_1827,N_121,N_1066);
xnor U1828 (N_1828,N_102,N_738);
and U1829 (N_1829,N_988,N_417);
or U1830 (N_1830,N_1137,N_170);
and U1831 (N_1831,N_160,N_457);
or U1832 (N_1832,N_1308,N_214);
nand U1833 (N_1833,N_1112,N_359);
nor U1834 (N_1834,N_364,N_1101);
nor U1835 (N_1835,N_963,N_1084);
nor U1836 (N_1836,N_1067,N_819);
and U1837 (N_1837,N_327,N_1261);
xnor U1838 (N_1838,N_965,N_521);
xor U1839 (N_1839,N_801,N_1315);
or U1840 (N_1840,N_30,N_481);
or U1841 (N_1841,N_473,N_1380);
and U1842 (N_1842,N_129,N_408);
and U1843 (N_1843,N_508,N_247);
or U1844 (N_1844,N_43,N_465);
nand U1845 (N_1845,N_456,N_901);
and U1846 (N_1846,N_932,N_987);
nor U1847 (N_1847,N_1365,N_1049);
xor U1848 (N_1848,N_1300,N_243);
nand U1849 (N_1849,N_320,N_1001);
xor U1850 (N_1850,N_313,N_1421);
nor U1851 (N_1851,N_1461,N_1025);
nand U1852 (N_1852,N_389,N_1171);
nand U1853 (N_1853,N_199,N_1154);
and U1854 (N_1854,N_1382,N_964);
and U1855 (N_1855,N_232,N_962);
or U1856 (N_1856,N_722,N_1108);
or U1857 (N_1857,N_285,N_1215);
or U1858 (N_1858,N_1207,N_943);
and U1859 (N_1859,N_1306,N_718);
and U1860 (N_1860,N_440,N_594);
and U1861 (N_1861,N_1092,N_1379);
nand U1862 (N_1862,N_51,N_861);
xor U1863 (N_1863,N_977,N_1173);
or U1864 (N_1864,N_999,N_959);
or U1865 (N_1865,N_386,N_692);
or U1866 (N_1866,N_541,N_439);
nand U1867 (N_1867,N_693,N_1008);
or U1868 (N_1868,N_694,N_149);
and U1869 (N_1869,N_533,N_1160);
nand U1870 (N_1870,N_171,N_653);
or U1871 (N_1871,N_204,N_610);
or U1872 (N_1872,N_120,N_1002);
nor U1873 (N_1873,N_462,N_1162);
and U1874 (N_1874,N_215,N_1374);
xor U1875 (N_1875,N_980,N_221);
and U1876 (N_1876,N_826,N_908);
nor U1877 (N_1877,N_1031,N_605);
nor U1878 (N_1878,N_245,N_1172);
nor U1879 (N_1879,N_597,N_1489);
xnor U1880 (N_1880,N_829,N_224);
nand U1881 (N_1881,N_704,N_577);
or U1882 (N_1882,N_1240,N_491);
nand U1883 (N_1883,N_368,N_1130);
nor U1884 (N_1884,N_874,N_807);
and U1885 (N_1885,N_1074,N_374);
or U1886 (N_1886,N_678,N_88);
or U1887 (N_1887,N_809,N_1332);
or U1888 (N_1888,N_319,N_476);
nor U1889 (N_1889,N_979,N_276);
nand U1890 (N_1890,N_922,N_633);
nor U1891 (N_1891,N_250,N_545);
or U1892 (N_1892,N_180,N_968);
nor U1893 (N_1893,N_301,N_818);
nor U1894 (N_1894,N_278,N_1149);
nand U1895 (N_1895,N_300,N_1147);
nor U1896 (N_1896,N_698,N_1125);
xor U1897 (N_1897,N_1209,N_459);
nor U1898 (N_1898,N_1305,N_773);
and U1899 (N_1899,N_134,N_856);
or U1900 (N_1900,N_505,N_308);
nand U1901 (N_1901,N_881,N_1381);
nand U1902 (N_1902,N_382,N_367);
nor U1903 (N_1903,N_402,N_325);
nand U1904 (N_1904,N_1006,N_122);
nand U1905 (N_1905,N_142,N_1163);
and U1906 (N_1906,N_1167,N_342);
and U1907 (N_1907,N_1188,N_307);
nor U1908 (N_1908,N_702,N_28);
and U1909 (N_1909,N_50,N_951);
nand U1910 (N_1910,N_151,N_739);
or U1911 (N_1911,N_885,N_130);
and U1912 (N_1912,N_73,N_15);
nand U1913 (N_1913,N_8,N_421);
or U1914 (N_1914,N_443,N_1175);
nand U1915 (N_1915,N_948,N_227);
or U1916 (N_1916,N_1355,N_990);
or U1917 (N_1917,N_233,N_792);
nor U1918 (N_1918,N_157,N_471);
nand U1919 (N_1919,N_1392,N_274);
nand U1920 (N_1920,N_883,N_747);
nand U1921 (N_1921,N_207,N_905);
nand U1922 (N_1922,N_1454,N_376);
nand U1923 (N_1923,N_1401,N_238);
or U1924 (N_1924,N_1474,N_719);
nor U1925 (N_1925,N_590,N_460);
nor U1926 (N_1926,N_246,N_1398);
or U1927 (N_1927,N_1356,N_1197);
xnor U1928 (N_1928,N_635,N_711);
and U1929 (N_1929,N_1433,N_1083);
and U1930 (N_1930,N_716,N_297);
nor U1931 (N_1931,N_1260,N_1391);
nor U1932 (N_1932,N_163,N_1499);
nand U1933 (N_1933,N_519,N_1330);
xnor U1934 (N_1934,N_1258,N_218);
nand U1935 (N_1935,N_339,N_343);
nor U1936 (N_1936,N_740,N_14);
nand U1937 (N_1937,N_1118,N_1449);
nand U1938 (N_1938,N_798,N_578);
nand U1939 (N_1939,N_455,N_1205);
and U1940 (N_1940,N_697,N_1486);
nand U1941 (N_1941,N_656,N_429);
nor U1942 (N_1942,N_996,N_654);
and U1943 (N_1943,N_244,N_627);
nand U1944 (N_1944,N_931,N_485);
nand U1945 (N_1945,N_562,N_935);
or U1946 (N_1946,N_1361,N_822);
xor U1947 (N_1947,N_1345,N_529);
and U1948 (N_1948,N_797,N_1259);
nor U1949 (N_1949,N_1077,N_435);
nor U1950 (N_1950,N_657,N_391);
nand U1951 (N_1951,N_689,N_1318);
nand U1952 (N_1952,N_753,N_428);
or U1953 (N_1953,N_1400,N_1114);
nand U1954 (N_1954,N_813,N_802);
or U1955 (N_1955,N_1220,N_1121);
nor U1956 (N_1956,N_44,N_1224);
nand U1957 (N_1957,N_599,N_68);
or U1958 (N_1958,N_33,N_365);
nand U1959 (N_1959,N_926,N_1349);
and U1960 (N_1960,N_195,N_322);
and U1961 (N_1961,N_1,N_1021);
xor U1962 (N_1962,N_1060,N_1329);
and U1963 (N_1963,N_618,N_127);
nand U1964 (N_1964,N_1427,N_114);
and U1965 (N_1965,N_1424,N_516);
nand U1966 (N_1966,N_270,N_779);
or U1967 (N_1967,N_213,N_1208);
or U1968 (N_1968,N_1252,N_5);
and U1969 (N_1969,N_1399,N_781);
nor U1970 (N_1970,N_272,N_900);
nand U1971 (N_1971,N_1181,N_1346);
nand U1972 (N_1972,N_855,N_1402);
nor U1973 (N_1973,N_1144,N_1491);
nand U1974 (N_1974,N_1056,N_1422);
and U1975 (N_1975,N_824,N_415);
and U1976 (N_1976,N_1323,N_641);
or U1977 (N_1977,N_961,N_878);
xnor U1978 (N_1978,N_256,N_1169);
nor U1979 (N_1979,N_1097,N_9);
nand U1980 (N_1980,N_538,N_725);
nand U1981 (N_1981,N_217,N_1273);
nor U1982 (N_1982,N_1028,N_1076);
nand U1983 (N_1983,N_774,N_175);
nand U1984 (N_1984,N_638,N_430);
and U1985 (N_1985,N_370,N_1414);
nand U1986 (N_1986,N_1284,N_167);
nand U1987 (N_1987,N_144,N_202);
xnor U1988 (N_1988,N_1363,N_1063);
or U1989 (N_1989,N_543,N_703);
xnor U1990 (N_1990,N_332,N_1458);
or U1991 (N_1991,N_966,N_419);
and U1992 (N_1992,N_1255,N_511);
nand U1993 (N_1993,N_412,N_1225);
and U1994 (N_1994,N_331,N_1004);
xnor U1995 (N_1995,N_1405,N_225);
or U1996 (N_1996,N_914,N_1103);
and U1997 (N_1997,N_1327,N_184);
nand U1998 (N_1998,N_264,N_1340);
and U1999 (N_1999,N_928,N_309);
and U2000 (N_2000,N_1265,N_496);
and U2001 (N_2001,N_54,N_1359);
and U2002 (N_2002,N_1251,N_1447);
or U2003 (N_2003,N_1322,N_234);
and U2004 (N_2004,N_1331,N_1440);
nor U2005 (N_2005,N_770,N_1245);
or U2006 (N_2006,N_1176,N_1413);
nor U2007 (N_2007,N_1104,N_299);
or U2008 (N_2008,N_289,N_510);
nor U2009 (N_2009,N_793,N_1055);
xor U2010 (N_2010,N_664,N_851);
and U2011 (N_2011,N_450,N_816);
nand U2012 (N_2012,N_630,N_1227);
nor U2013 (N_2013,N_230,N_927);
nor U2014 (N_2014,N_92,N_1253);
nand U2015 (N_2015,N_710,N_400);
nor U2016 (N_2016,N_189,N_1480);
nor U2017 (N_2017,N_91,N_48);
nand U2018 (N_2018,N_257,N_799);
or U2019 (N_2019,N_128,N_173);
nand U2020 (N_2020,N_721,N_542);
xor U2021 (N_2021,N_116,N_1042);
nor U2022 (N_2022,N_290,N_531);
nor U2023 (N_2023,N_1455,N_839);
nor U2024 (N_2024,N_836,N_1434);
xor U2025 (N_2025,N_1388,N_433);
and U2026 (N_2026,N_1292,N_1481);
xor U2027 (N_2027,N_1256,N_513);
nor U2028 (N_2028,N_967,N_1229);
nor U2029 (N_2029,N_850,N_731);
and U2030 (N_2030,N_609,N_47);
or U2031 (N_2031,N_458,N_1218);
nand U2032 (N_2032,N_1320,N_1354);
nand U2033 (N_2033,N_395,N_1142);
or U2034 (N_2034,N_1143,N_737);
nor U2035 (N_2035,N_20,N_363);
nor U2036 (N_2036,N_1432,N_690);
nand U2037 (N_2037,N_106,N_659);
nand U2038 (N_2038,N_820,N_925);
xor U2039 (N_2039,N_1484,N_346);
nor U2040 (N_2040,N_1428,N_1465);
nor U2041 (N_2041,N_811,N_1479);
and U2042 (N_2042,N_617,N_1053);
xnor U2043 (N_2043,N_841,N_1236);
and U2044 (N_2044,N_1041,N_1282);
and U2045 (N_2045,N_281,N_494);
or U2046 (N_2046,N_930,N_292);
or U2047 (N_2047,N_228,N_860);
nor U2048 (N_2048,N_360,N_582);
and U2049 (N_2049,N_377,N_1230);
nand U2050 (N_2050,N_66,N_558);
or U2051 (N_2051,N_53,N_341);
and U2052 (N_2052,N_1073,N_304);
nor U2053 (N_2053,N_1448,N_1195);
xor U2054 (N_2054,N_423,N_1036);
and U2055 (N_2055,N_490,N_1179);
or U2056 (N_2056,N_1344,N_668);
or U2057 (N_2057,N_132,N_140);
xor U2058 (N_2058,N_876,N_1193);
or U2059 (N_2059,N_1132,N_318);
nor U2060 (N_2060,N_1296,N_648);
or U2061 (N_2061,N_902,N_118);
nand U2062 (N_2062,N_756,N_1124);
and U2063 (N_2063,N_1367,N_113);
nor U2064 (N_2064,N_59,N_328);
and U2065 (N_2065,N_866,N_139);
or U2066 (N_2066,N_745,N_1116);
and U2067 (N_2067,N_869,N_1372);
or U2068 (N_2068,N_939,N_1407);
nand U2069 (N_2069,N_437,N_1091);
and U2070 (N_2070,N_275,N_438);
nor U2071 (N_2071,N_969,N_957);
nand U2072 (N_2072,N_1362,N_466);
nor U2073 (N_2073,N_651,N_39);
and U2074 (N_2074,N_1174,N_1478);
and U2075 (N_2075,N_1192,N_847);
and U2076 (N_2076,N_576,N_588);
nand U2077 (N_2077,N_258,N_283);
and U2078 (N_2078,N_248,N_104);
nor U2079 (N_2079,N_109,N_267);
or U2080 (N_2080,N_911,N_1254);
or U2081 (N_2081,N_547,N_373);
nor U2082 (N_2082,N_536,N_1135);
and U2083 (N_2083,N_865,N_1450);
or U2084 (N_2084,N_846,N_572);
or U2085 (N_2085,N_1378,N_528);
nand U2086 (N_2086,N_1275,N_544);
and U2087 (N_2087,N_385,N_483);
nor U2088 (N_2088,N_115,N_613);
xor U2089 (N_2089,N_845,N_1187);
nor U2090 (N_2090,N_658,N_413);
and U2091 (N_2091,N_62,N_291);
xor U2092 (N_2092,N_1212,N_843);
and U2093 (N_2093,N_436,N_183);
xor U2094 (N_2094,N_472,N_560);
nor U2095 (N_2095,N_875,N_1081);
nor U2096 (N_2096,N_933,N_1495);
or U2097 (N_2097,N_647,N_1068);
or U2098 (N_2098,N_187,N_769);
or U2099 (N_2099,N_226,N_1357);
and U2100 (N_2100,N_838,N_643);
nor U2101 (N_2101,N_1026,N_384);
and U2102 (N_2102,N_1239,N_1243);
nor U2103 (N_2103,N_1431,N_380);
nor U2104 (N_2104,N_1159,N_887);
nor U2105 (N_2105,N_1462,N_119);
or U2106 (N_2106,N_699,N_392);
nor U2107 (N_2107,N_986,N_1280);
and U2108 (N_2108,N_625,N_1335);
and U2109 (N_2109,N_520,N_265);
nor U2110 (N_2110,N_70,N_759);
nand U2111 (N_2111,N_1250,N_844);
nor U2112 (N_2112,N_1235,N_169);
or U2113 (N_2113,N_849,N_152);
or U2114 (N_2114,N_995,N_1221);
nor U2115 (N_2115,N_1324,N_1095);
nor U2116 (N_2116,N_198,N_424);
and U2117 (N_2117,N_917,N_650);
nand U2118 (N_2118,N_858,N_1126);
or U2119 (N_2119,N_1420,N_1019);
or U2120 (N_2120,N_347,N_754);
nor U2121 (N_2121,N_1050,N_1276);
nand U2122 (N_2122,N_1472,N_1246);
nor U2123 (N_2123,N_467,N_1466);
or U2124 (N_2124,N_1279,N_77);
and U2125 (N_2125,N_315,N_1198);
nand U2126 (N_2126,N_136,N_482);
nand U2127 (N_2127,N_156,N_1460);
and U2128 (N_2128,N_111,N_220);
and U2129 (N_2129,N_947,N_337);
and U2130 (N_2130,N_1241,N_1406);
or U2131 (N_2131,N_486,N_1311);
or U2132 (N_2132,N_10,N_530);
nor U2133 (N_2133,N_1294,N_591);
and U2134 (N_2134,N_407,N_1410);
or U2135 (N_2135,N_1376,N_1199);
nand U2136 (N_2136,N_29,N_148);
and U2137 (N_2137,N_1138,N_349);
xor U2138 (N_2138,N_251,N_1277);
or U2139 (N_2139,N_452,N_1351);
nand U2140 (N_2140,N_837,N_381);
nand U2141 (N_2141,N_1429,N_1166);
xnor U2142 (N_2142,N_726,N_600);
nand U2143 (N_2143,N_353,N_941);
and U2144 (N_2144,N_563,N_375);
nor U2145 (N_2145,N_629,N_1165);
or U2146 (N_2146,N_686,N_1061);
nor U2147 (N_2147,N_805,N_665);
nor U2148 (N_2148,N_345,N_0);
nand U2149 (N_2149,N_978,N_776);
and U2150 (N_2150,N_975,N_1016);
and U2151 (N_2151,N_765,N_921);
nand U2152 (N_2152,N_3,N_994);
and U2153 (N_2153,N_27,N_706);
xnor U2154 (N_2154,N_1185,N_1222);
nor U2155 (N_2155,N_1342,N_912);
or U2156 (N_2156,N_397,N_626);
nor U2157 (N_2157,N_815,N_755);
nor U2158 (N_2158,N_566,N_1353);
and U2159 (N_2159,N_1139,N_1140);
nand U2160 (N_2160,N_1456,N_416);
xnor U2161 (N_2161,N_730,N_67);
and U2162 (N_2162,N_871,N_178);
nand U2163 (N_2163,N_282,N_447);
and U2164 (N_2164,N_886,N_4);
or U2165 (N_2165,N_972,N_864);
and U2166 (N_2166,N_158,N_1492);
and U2167 (N_2167,N_1387,N_1316);
and U2168 (N_2168,N_857,N_848);
nor U2169 (N_2169,N_1459,N_1483);
xor U2170 (N_2170,N_1100,N_99);
nor U2171 (N_2171,N_895,N_762);
and U2172 (N_2172,N_614,N_1442);
xor U2173 (N_2173,N_946,N_1370);
or U2174 (N_2174,N_634,N_164);
and U2175 (N_2175,N_209,N_361);
nand U2176 (N_2176,N_938,N_266);
or U2177 (N_2177,N_1496,N_396);
xor U2178 (N_2178,N_1384,N_944);
and U2179 (N_2179,N_937,N_1178);
and U2180 (N_2180,N_61,N_889);
nand U2181 (N_2181,N_894,N_1291);
nor U2182 (N_2182,N_680,N_760);
nor U2183 (N_2183,N_785,N_1090);
xnor U2184 (N_2184,N_863,N_235);
nand U2185 (N_2185,N_1403,N_852);
or U2186 (N_2186,N_976,N_608);
nand U2187 (N_2187,N_749,N_775);
and U2188 (N_2188,N_1321,N_840);
nor U2189 (N_2189,N_1416,N_896);
and U2190 (N_2190,N_254,N_565);
xnor U2191 (N_2191,N_970,N_1383);
and U2192 (N_2192,N_758,N_503);
or U2193 (N_2193,N_1153,N_1475);
nor U2194 (N_2194,N_255,N_1237);
nand U2195 (N_2195,N_518,N_714);
nand U2196 (N_2196,N_661,N_1214);
and U2197 (N_2197,N_611,N_177);
nand U2198 (N_2198,N_899,N_1111);
nand U2199 (N_2199,N_771,N_1011);
and U2200 (N_2200,N_791,N_82);
or U2201 (N_2201,N_150,N_185);
nand U2202 (N_2202,N_1182,N_620);
nor U2203 (N_2203,N_269,N_1352);
nor U2204 (N_2204,N_575,N_1117);
nor U2205 (N_2205,N_371,N_1216);
nor U2206 (N_2206,N_117,N_555);
nor U2207 (N_2207,N_165,N_1030);
or U2208 (N_2208,N_1027,N_426);
nor U2209 (N_2209,N_229,N_86);
and U2210 (N_2210,N_1190,N_74);
or U2211 (N_2211,N_26,N_203);
or U2212 (N_2212,N_573,N_181);
and U2213 (N_2213,N_1477,N_193);
or U2214 (N_2214,N_602,N_1435);
nor U2215 (N_2215,N_579,N_1106);
xor U2216 (N_2216,N_1326,N_1263);
nand U2217 (N_2217,N_552,N_90);
or U2218 (N_2218,N_1293,N_595);
nor U2219 (N_2219,N_147,N_1302);
and U2220 (N_2220,N_280,N_750);
nor U2221 (N_2221,N_517,N_1223);
xnor U2222 (N_2222,N_1389,N_1040);
or U2223 (N_2223,N_1183,N_736);
nor U2224 (N_2224,N_786,N_85);
and U2225 (N_2225,N_1397,N_83);
nor U2226 (N_2226,N_1281,N_1072);
or U2227 (N_2227,N_806,N_1343);
nor U2228 (N_2228,N_991,N_236);
nor U2229 (N_2229,N_768,N_671);
and U2230 (N_2230,N_1131,N_1122);
or U2231 (N_2231,N_1364,N_708);
nor U2232 (N_2232,N_1189,N_955);
xor U2233 (N_2233,N_298,N_763);
and U2234 (N_2234,N_717,N_1301);
nand U2235 (N_2235,N_296,N_1490);
nand U2236 (N_2236,N_240,N_464);
nand U2237 (N_2237,N_34,N_723);
nand U2238 (N_2238,N_1048,N_1487);
nor U2239 (N_2239,N_550,N_1059);
or U2240 (N_2240,N_1269,N_669);
and U2241 (N_2241,N_788,N_399);
or U2242 (N_2242,N_971,N_945);
nor U2243 (N_2243,N_123,N_1419);
nand U2244 (N_2244,N_497,N_870);
nand U2245 (N_2245,N_1018,N_1115);
nor U2246 (N_2246,N_393,N_21);
or U2247 (N_2247,N_1244,N_580);
or U2248 (N_2248,N_1158,N_539);
xnor U2249 (N_2249,N_1266,N_110);
or U2250 (N_2250,N_8,N_504);
nor U2251 (N_2251,N_1113,N_1152);
xnor U2252 (N_2252,N_1364,N_52);
or U2253 (N_2253,N_922,N_1070);
or U2254 (N_2254,N_1420,N_939);
or U2255 (N_2255,N_723,N_1028);
or U2256 (N_2256,N_336,N_905);
and U2257 (N_2257,N_1402,N_109);
nand U2258 (N_2258,N_193,N_844);
nor U2259 (N_2259,N_243,N_892);
nor U2260 (N_2260,N_404,N_1199);
nand U2261 (N_2261,N_496,N_1166);
nor U2262 (N_2262,N_788,N_1028);
and U2263 (N_2263,N_1214,N_1056);
nor U2264 (N_2264,N_1072,N_1255);
nor U2265 (N_2265,N_823,N_1462);
nor U2266 (N_2266,N_1044,N_817);
and U2267 (N_2267,N_511,N_351);
nor U2268 (N_2268,N_48,N_438);
and U2269 (N_2269,N_988,N_325);
xor U2270 (N_2270,N_1435,N_10);
or U2271 (N_2271,N_1363,N_759);
nand U2272 (N_2272,N_57,N_497);
xor U2273 (N_2273,N_882,N_1203);
nand U2274 (N_2274,N_1110,N_61);
and U2275 (N_2275,N_50,N_1119);
nor U2276 (N_2276,N_690,N_876);
nand U2277 (N_2277,N_1498,N_586);
nand U2278 (N_2278,N_458,N_569);
nand U2279 (N_2279,N_149,N_266);
nand U2280 (N_2280,N_557,N_1195);
nand U2281 (N_2281,N_752,N_519);
nor U2282 (N_2282,N_825,N_785);
nor U2283 (N_2283,N_181,N_89);
nand U2284 (N_2284,N_396,N_517);
nor U2285 (N_2285,N_1457,N_1320);
or U2286 (N_2286,N_1282,N_267);
nor U2287 (N_2287,N_84,N_799);
nand U2288 (N_2288,N_1141,N_1390);
xnor U2289 (N_2289,N_1187,N_578);
nand U2290 (N_2290,N_578,N_1443);
and U2291 (N_2291,N_372,N_183);
nand U2292 (N_2292,N_1108,N_749);
or U2293 (N_2293,N_1477,N_653);
nor U2294 (N_2294,N_1013,N_671);
nor U2295 (N_2295,N_1141,N_954);
nor U2296 (N_2296,N_652,N_482);
and U2297 (N_2297,N_1199,N_1149);
nor U2298 (N_2298,N_332,N_1006);
and U2299 (N_2299,N_120,N_1345);
nor U2300 (N_2300,N_579,N_841);
or U2301 (N_2301,N_743,N_377);
or U2302 (N_2302,N_397,N_151);
and U2303 (N_2303,N_110,N_502);
nor U2304 (N_2304,N_869,N_1335);
nor U2305 (N_2305,N_1299,N_241);
nand U2306 (N_2306,N_650,N_1310);
nand U2307 (N_2307,N_1495,N_19);
nand U2308 (N_2308,N_438,N_661);
nor U2309 (N_2309,N_487,N_792);
nor U2310 (N_2310,N_166,N_508);
nand U2311 (N_2311,N_400,N_47);
and U2312 (N_2312,N_645,N_972);
nor U2313 (N_2313,N_296,N_1480);
xnor U2314 (N_2314,N_323,N_1153);
or U2315 (N_2315,N_401,N_927);
and U2316 (N_2316,N_251,N_287);
or U2317 (N_2317,N_327,N_86);
nor U2318 (N_2318,N_1380,N_1453);
nor U2319 (N_2319,N_1091,N_757);
nor U2320 (N_2320,N_699,N_1279);
xor U2321 (N_2321,N_968,N_88);
nand U2322 (N_2322,N_791,N_1230);
xnor U2323 (N_2323,N_875,N_640);
and U2324 (N_2324,N_201,N_1186);
nand U2325 (N_2325,N_1393,N_1248);
nand U2326 (N_2326,N_1276,N_1306);
or U2327 (N_2327,N_363,N_885);
and U2328 (N_2328,N_260,N_1087);
or U2329 (N_2329,N_1247,N_326);
or U2330 (N_2330,N_1419,N_954);
xor U2331 (N_2331,N_1144,N_529);
nand U2332 (N_2332,N_394,N_1057);
or U2333 (N_2333,N_184,N_672);
xnor U2334 (N_2334,N_781,N_1448);
and U2335 (N_2335,N_645,N_947);
and U2336 (N_2336,N_167,N_1166);
xor U2337 (N_2337,N_925,N_462);
or U2338 (N_2338,N_503,N_168);
and U2339 (N_2339,N_311,N_650);
nand U2340 (N_2340,N_842,N_1129);
nor U2341 (N_2341,N_652,N_339);
nand U2342 (N_2342,N_338,N_406);
and U2343 (N_2343,N_452,N_485);
nor U2344 (N_2344,N_77,N_1458);
xor U2345 (N_2345,N_931,N_1065);
nor U2346 (N_2346,N_1255,N_848);
or U2347 (N_2347,N_998,N_1017);
nor U2348 (N_2348,N_460,N_760);
nand U2349 (N_2349,N_1319,N_1020);
or U2350 (N_2350,N_672,N_854);
and U2351 (N_2351,N_1450,N_1269);
and U2352 (N_2352,N_1135,N_12);
xor U2353 (N_2353,N_461,N_710);
or U2354 (N_2354,N_583,N_630);
xnor U2355 (N_2355,N_862,N_972);
and U2356 (N_2356,N_282,N_60);
or U2357 (N_2357,N_892,N_374);
nor U2358 (N_2358,N_1171,N_1209);
or U2359 (N_2359,N_1425,N_946);
and U2360 (N_2360,N_1123,N_476);
and U2361 (N_2361,N_655,N_137);
nand U2362 (N_2362,N_1325,N_966);
nor U2363 (N_2363,N_399,N_533);
nand U2364 (N_2364,N_55,N_157);
or U2365 (N_2365,N_156,N_603);
or U2366 (N_2366,N_698,N_1120);
or U2367 (N_2367,N_802,N_1177);
nand U2368 (N_2368,N_831,N_1077);
nand U2369 (N_2369,N_229,N_976);
xor U2370 (N_2370,N_116,N_627);
nor U2371 (N_2371,N_193,N_609);
or U2372 (N_2372,N_278,N_1158);
nor U2373 (N_2373,N_1303,N_240);
xnor U2374 (N_2374,N_1236,N_1155);
nand U2375 (N_2375,N_110,N_1115);
nand U2376 (N_2376,N_459,N_1374);
and U2377 (N_2377,N_944,N_506);
nor U2378 (N_2378,N_1405,N_1399);
or U2379 (N_2379,N_1341,N_112);
nand U2380 (N_2380,N_229,N_1344);
or U2381 (N_2381,N_1087,N_1070);
or U2382 (N_2382,N_1401,N_52);
or U2383 (N_2383,N_409,N_270);
nor U2384 (N_2384,N_421,N_1092);
and U2385 (N_2385,N_636,N_698);
or U2386 (N_2386,N_44,N_378);
and U2387 (N_2387,N_432,N_1463);
and U2388 (N_2388,N_1380,N_328);
nor U2389 (N_2389,N_1107,N_996);
nor U2390 (N_2390,N_289,N_923);
and U2391 (N_2391,N_688,N_1067);
or U2392 (N_2392,N_849,N_996);
nand U2393 (N_2393,N_600,N_919);
or U2394 (N_2394,N_289,N_1055);
xnor U2395 (N_2395,N_550,N_1420);
or U2396 (N_2396,N_807,N_1358);
nand U2397 (N_2397,N_521,N_818);
nand U2398 (N_2398,N_930,N_1419);
and U2399 (N_2399,N_592,N_576);
or U2400 (N_2400,N_1292,N_475);
nor U2401 (N_2401,N_488,N_859);
nand U2402 (N_2402,N_718,N_118);
nor U2403 (N_2403,N_769,N_715);
and U2404 (N_2404,N_1459,N_1404);
nand U2405 (N_2405,N_316,N_3);
xor U2406 (N_2406,N_914,N_1405);
nor U2407 (N_2407,N_728,N_816);
nor U2408 (N_2408,N_202,N_200);
and U2409 (N_2409,N_179,N_128);
xnor U2410 (N_2410,N_177,N_1243);
nor U2411 (N_2411,N_425,N_521);
and U2412 (N_2412,N_666,N_49);
or U2413 (N_2413,N_1455,N_1202);
or U2414 (N_2414,N_535,N_745);
nor U2415 (N_2415,N_622,N_1066);
xnor U2416 (N_2416,N_1092,N_10);
nand U2417 (N_2417,N_208,N_1483);
and U2418 (N_2418,N_729,N_855);
nand U2419 (N_2419,N_285,N_1355);
or U2420 (N_2420,N_439,N_593);
and U2421 (N_2421,N_1058,N_21);
nor U2422 (N_2422,N_1215,N_1030);
xnor U2423 (N_2423,N_943,N_1264);
nor U2424 (N_2424,N_1482,N_1171);
and U2425 (N_2425,N_58,N_1034);
nand U2426 (N_2426,N_934,N_941);
and U2427 (N_2427,N_277,N_883);
and U2428 (N_2428,N_210,N_1405);
nor U2429 (N_2429,N_736,N_245);
nand U2430 (N_2430,N_335,N_259);
nor U2431 (N_2431,N_281,N_547);
or U2432 (N_2432,N_392,N_2);
nand U2433 (N_2433,N_606,N_1407);
and U2434 (N_2434,N_1394,N_1498);
nand U2435 (N_2435,N_747,N_1152);
and U2436 (N_2436,N_938,N_531);
xor U2437 (N_2437,N_1177,N_1084);
and U2438 (N_2438,N_1375,N_638);
xnor U2439 (N_2439,N_587,N_573);
nand U2440 (N_2440,N_844,N_1386);
and U2441 (N_2441,N_334,N_1099);
and U2442 (N_2442,N_1193,N_24);
and U2443 (N_2443,N_1215,N_198);
nand U2444 (N_2444,N_206,N_11);
nand U2445 (N_2445,N_895,N_1484);
or U2446 (N_2446,N_1204,N_265);
and U2447 (N_2447,N_863,N_607);
nor U2448 (N_2448,N_32,N_1410);
nor U2449 (N_2449,N_1346,N_964);
nor U2450 (N_2450,N_810,N_19);
and U2451 (N_2451,N_1037,N_567);
and U2452 (N_2452,N_1356,N_272);
nor U2453 (N_2453,N_211,N_323);
nand U2454 (N_2454,N_593,N_407);
and U2455 (N_2455,N_230,N_166);
or U2456 (N_2456,N_337,N_1380);
xnor U2457 (N_2457,N_230,N_1193);
nand U2458 (N_2458,N_1262,N_443);
nand U2459 (N_2459,N_928,N_801);
nor U2460 (N_2460,N_210,N_1073);
or U2461 (N_2461,N_843,N_353);
or U2462 (N_2462,N_1104,N_1235);
and U2463 (N_2463,N_103,N_968);
xor U2464 (N_2464,N_806,N_1016);
nand U2465 (N_2465,N_753,N_217);
nor U2466 (N_2466,N_1283,N_102);
or U2467 (N_2467,N_775,N_555);
or U2468 (N_2468,N_1467,N_857);
nor U2469 (N_2469,N_1322,N_148);
nor U2470 (N_2470,N_1432,N_683);
xnor U2471 (N_2471,N_58,N_762);
nand U2472 (N_2472,N_844,N_252);
nor U2473 (N_2473,N_444,N_22);
and U2474 (N_2474,N_32,N_1313);
and U2475 (N_2475,N_30,N_602);
and U2476 (N_2476,N_1021,N_1125);
and U2477 (N_2477,N_696,N_780);
and U2478 (N_2478,N_138,N_1417);
nor U2479 (N_2479,N_340,N_1409);
or U2480 (N_2480,N_55,N_546);
and U2481 (N_2481,N_1031,N_920);
nor U2482 (N_2482,N_126,N_1169);
nand U2483 (N_2483,N_1309,N_111);
nand U2484 (N_2484,N_454,N_1437);
nor U2485 (N_2485,N_127,N_1419);
nor U2486 (N_2486,N_12,N_1213);
nor U2487 (N_2487,N_198,N_1401);
and U2488 (N_2488,N_1166,N_1093);
nor U2489 (N_2489,N_611,N_329);
or U2490 (N_2490,N_1163,N_334);
and U2491 (N_2491,N_548,N_21);
and U2492 (N_2492,N_199,N_1227);
or U2493 (N_2493,N_556,N_606);
xnor U2494 (N_2494,N_652,N_615);
and U2495 (N_2495,N_301,N_137);
or U2496 (N_2496,N_915,N_1416);
or U2497 (N_2497,N_835,N_1259);
xnor U2498 (N_2498,N_1283,N_1135);
nor U2499 (N_2499,N_105,N_393);
nor U2500 (N_2500,N_995,N_843);
nor U2501 (N_2501,N_823,N_407);
and U2502 (N_2502,N_674,N_845);
xnor U2503 (N_2503,N_1256,N_1315);
nor U2504 (N_2504,N_799,N_1059);
xor U2505 (N_2505,N_706,N_1250);
and U2506 (N_2506,N_428,N_1183);
and U2507 (N_2507,N_1118,N_1414);
and U2508 (N_2508,N_627,N_1239);
or U2509 (N_2509,N_1455,N_1478);
nand U2510 (N_2510,N_248,N_1414);
or U2511 (N_2511,N_1485,N_636);
or U2512 (N_2512,N_293,N_852);
nor U2513 (N_2513,N_831,N_135);
and U2514 (N_2514,N_388,N_1386);
or U2515 (N_2515,N_1173,N_403);
or U2516 (N_2516,N_484,N_395);
and U2517 (N_2517,N_845,N_0);
nor U2518 (N_2518,N_1330,N_534);
xnor U2519 (N_2519,N_1135,N_139);
xnor U2520 (N_2520,N_651,N_681);
and U2521 (N_2521,N_504,N_1432);
nor U2522 (N_2522,N_613,N_126);
nand U2523 (N_2523,N_272,N_1163);
and U2524 (N_2524,N_1238,N_1357);
and U2525 (N_2525,N_783,N_1142);
and U2526 (N_2526,N_852,N_1264);
and U2527 (N_2527,N_66,N_1311);
or U2528 (N_2528,N_375,N_531);
or U2529 (N_2529,N_1433,N_96);
and U2530 (N_2530,N_1474,N_1328);
nand U2531 (N_2531,N_368,N_356);
and U2532 (N_2532,N_1080,N_1187);
xor U2533 (N_2533,N_197,N_1321);
or U2534 (N_2534,N_345,N_723);
or U2535 (N_2535,N_1216,N_525);
nand U2536 (N_2536,N_642,N_482);
nand U2537 (N_2537,N_808,N_652);
nand U2538 (N_2538,N_656,N_1069);
xor U2539 (N_2539,N_642,N_312);
or U2540 (N_2540,N_550,N_1134);
nand U2541 (N_2541,N_1054,N_593);
nor U2542 (N_2542,N_350,N_19);
nor U2543 (N_2543,N_975,N_52);
nand U2544 (N_2544,N_346,N_246);
nor U2545 (N_2545,N_613,N_1468);
nand U2546 (N_2546,N_954,N_835);
nand U2547 (N_2547,N_446,N_385);
nand U2548 (N_2548,N_723,N_627);
nor U2549 (N_2549,N_1314,N_1252);
nand U2550 (N_2550,N_588,N_898);
xnor U2551 (N_2551,N_1324,N_792);
nor U2552 (N_2552,N_957,N_533);
nor U2553 (N_2553,N_421,N_680);
nor U2554 (N_2554,N_152,N_883);
or U2555 (N_2555,N_224,N_291);
nand U2556 (N_2556,N_1012,N_895);
or U2557 (N_2557,N_1491,N_1390);
or U2558 (N_2558,N_808,N_1035);
or U2559 (N_2559,N_1327,N_1462);
and U2560 (N_2560,N_751,N_47);
xnor U2561 (N_2561,N_1410,N_1031);
or U2562 (N_2562,N_84,N_909);
nand U2563 (N_2563,N_180,N_688);
nor U2564 (N_2564,N_289,N_145);
and U2565 (N_2565,N_408,N_986);
and U2566 (N_2566,N_427,N_1054);
or U2567 (N_2567,N_153,N_1470);
or U2568 (N_2568,N_556,N_1231);
and U2569 (N_2569,N_382,N_1092);
and U2570 (N_2570,N_906,N_1301);
and U2571 (N_2571,N_109,N_1091);
nor U2572 (N_2572,N_1182,N_913);
and U2573 (N_2573,N_641,N_509);
nor U2574 (N_2574,N_764,N_1223);
and U2575 (N_2575,N_955,N_907);
nand U2576 (N_2576,N_52,N_564);
nand U2577 (N_2577,N_293,N_1146);
nor U2578 (N_2578,N_294,N_1288);
or U2579 (N_2579,N_1046,N_1462);
nand U2580 (N_2580,N_1040,N_456);
and U2581 (N_2581,N_1088,N_385);
or U2582 (N_2582,N_1489,N_257);
or U2583 (N_2583,N_715,N_1223);
and U2584 (N_2584,N_416,N_1392);
and U2585 (N_2585,N_32,N_1232);
nor U2586 (N_2586,N_386,N_1036);
and U2587 (N_2587,N_456,N_24);
and U2588 (N_2588,N_611,N_455);
and U2589 (N_2589,N_1332,N_157);
or U2590 (N_2590,N_1496,N_291);
and U2591 (N_2591,N_34,N_788);
xor U2592 (N_2592,N_320,N_508);
xnor U2593 (N_2593,N_881,N_586);
or U2594 (N_2594,N_1380,N_779);
and U2595 (N_2595,N_910,N_654);
nand U2596 (N_2596,N_902,N_678);
or U2597 (N_2597,N_605,N_905);
nor U2598 (N_2598,N_1247,N_1481);
or U2599 (N_2599,N_797,N_1313);
xor U2600 (N_2600,N_99,N_1212);
and U2601 (N_2601,N_317,N_1050);
nand U2602 (N_2602,N_1420,N_829);
and U2603 (N_2603,N_51,N_395);
nor U2604 (N_2604,N_310,N_722);
nand U2605 (N_2605,N_492,N_1341);
and U2606 (N_2606,N_65,N_649);
nand U2607 (N_2607,N_322,N_837);
nand U2608 (N_2608,N_692,N_683);
nor U2609 (N_2609,N_872,N_681);
xnor U2610 (N_2610,N_678,N_564);
nand U2611 (N_2611,N_1008,N_719);
nand U2612 (N_2612,N_137,N_1356);
or U2613 (N_2613,N_1215,N_1457);
nand U2614 (N_2614,N_697,N_869);
and U2615 (N_2615,N_385,N_53);
or U2616 (N_2616,N_195,N_370);
nand U2617 (N_2617,N_909,N_530);
and U2618 (N_2618,N_725,N_1469);
or U2619 (N_2619,N_548,N_940);
nand U2620 (N_2620,N_1401,N_68);
or U2621 (N_2621,N_810,N_1014);
nor U2622 (N_2622,N_485,N_682);
nor U2623 (N_2623,N_1254,N_402);
or U2624 (N_2624,N_644,N_1330);
or U2625 (N_2625,N_1334,N_876);
nand U2626 (N_2626,N_1067,N_64);
xnor U2627 (N_2627,N_397,N_342);
nor U2628 (N_2628,N_514,N_915);
and U2629 (N_2629,N_659,N_1463);
or U2630 (N_2630,N_1338,N_951);
and U2631 (N_2631,N_91,N_132);
nand U2632 (N_2632,N_383,N_1181);
nor U2633 (N_2633,N_183,N_628);
or U2634 (N_2634,N_1318,N_380);
and U2635 (N_2635,N_844,N_1238);
nor U2636 (N_2636,N_883,N_1344);
nor U2637 (N_2637,N_129,N_249);
nor U2638 (N_2638,N_412,N_1440);
and U2639 (N_2639,N_725,N_1237);
and U2640 (N_2640,N_1161,N_1391);
or U2641 (N_2641,N_439,N_261);
nor U2642 (N_2642,N_259,N_1201);
or U2643 (N_2643,N_1219,N_470);
nand U2644 (N_2644,N_617,N_628);
nor U2645 (N_2645,N_934,N_680);
and U2646 (N_2646,N_734,N_840);
and U2647 (N_2647,N_572,N_1453);
nor U2648 (N_2648,N_1382,N_1428);
nand U2649 (N_2649,N_815,N_662);
nor U2650 (N_2650,N_412,N_1469);
and U2651 (N_2651,N_134,N_409);
nor U2652 (N_2652,N_1015,N_428);
or U2653 (N_2653,N_827,N_1165);
and U2654 (N_2654,N_668,N_866);
nor U2655 (N_2655,N_477,N_1155);
and U2656 (N_2656,N_1058,N_462);
xnor U2657 (N_2657,N_1211,N_64);
and U2658 (N_2658,N_1457,N_345);
or U2659 (N_2659,N_630,N_225);
and U2660 (N_2660,N_1487,N_433);
or U2661 (N_2661,N_293,N_272);
and U2662 (N_2662,N_237,N_1467);
or U2663 (N_2663,N_740,N_792);
nand U2664 (N_2664,N_391,N_1151);
nand U2665 (N_2665,N_1042,N_1201);
xnor U2666 (N_2666,N_877,N_1125);
xnor U2667 (N_2667,N_1414,N_1351);
and U2668 (N_2668,N_678,N_17);
and U2669 (N_2669,N_1467,N_1275);
nand U2670 (N_2670,N_38,N_848);
nand U2671 (N_2671,N_781,N_1491);
or U2672 (N_2672,N_760,N_1137);
nor U2673 (N_2673,N_545,N_364);
or U2674 (N_2674,N_1012,N_953);
nor U2675 (N_2675,N_1318,N_163);
and U2676 (N_2676,N_755,N_1340);
nand U2677 (N_2677,N_1317,N_354);
nand U2678 (N_2678,N_1292,N_1169);
nand U2679 (N_2679,N_1451,N_782);
nor U2680 (N_2680,N_270,N_146);
or U2681 (N_2681,N_1148,N_1132);
nor U2682 (N_2682,N_563,N_1378);
nor U2683 (N_2683,N_1497,N_529);
or U2684 (N_2684,N_80,N_1090);
or U2685 (N_2685,N_331,N_1133);
or U2686 (N_2686,N_498,N_1039);
and U2687 (N_2687,N_1039,N_1182);
or U2688 (N_2688,N_365,N_444);
and U2689 (N_2689,N_407,N_386);
nor U2690 (N_2690,N_1353,N_816);
xor U2691 (N_2691,N_167,N_1454);
and U2692 (N_2692,N_767,N_1008);
nor U2693 (N_2693,N_826,N_781);
xnor U2694 (N_2694,N_460,N_189);
xnor U2695 (N_2695,N_780,N_64);
or U2696 (N_2696,N_481,N_787);
and U2697 (N_2697,N_1474,N_236);
or U2698 (N_2698,N_511,N_703);
xor U2699 (N_2699,N_385,N_1368);
xnor U2700 (N_2700,N_1091,N_1352);
or U2701 (N_2701,N_1187,N_405);
or U2702 (N_2702,N_395,N_1034);
and U2703 (N_2703,N_724,N_101);
nand U2704 (N_2704,N_773,N_663);
nand U2705 (N_2705,N_1206,N_680);
nand U2706 (N_2706,N_179,N_136);
nand U2707 (N_2707,N_430,N_385);
nand U2708 (N_2708,N_156,N_1158);
xor U2709 (N_2709,N_1306,N_6);
and U2710 (N_2710,N_1205,N_553);
nand U2711 (N_2711,N_670,N_1459);
xor U2712 (N_2712,N_1133,N_163);
nor U2713 (N_2713,N_277,N_823);
nor U2714 (N_2714,N_1460,N_818);
nand U2715 (N_2715,N_461,N_764);
xnor U2716 (N_2716,N_396,N_1207);
nor U2717 (N_2717,N_720,N_409);
nor U2718 (N_2718,N_1348,N_538);
nand U2719 (N_2719,N_522,N_691);
or U2720 (N_2720,N_215,N_469);
and U2721 (N_2721,N_1354,N_399);
nor U2722 (N_2722,N_936,N_523);
or U2723 (N_2723,N_522,N_781);
nor U2724 (N_2724,N_594,N_1286);
or U2725 (N_2725,N_1194,N_122);
xnor U2726 (N_2726,N_523,N_1007);
or U2727 (N_2727,N_629,N_670);
nand U2728 (N_2728,N_758,N_197);
or U2729 (N_2729,N_729,N_1442);
or U2730 (N_2730,N_1072,N_898);
and U2731 (N_2731,N_939,N_979);
or U2732 (N_2732,N_60,N_1032);
nand U2733 (N_2733,N_1268,N_550);
nor U2734 (N_2734,N_202,N_1497);
nor U2735 (N_2735,N_798,N_1439);
nand U2736 (N_2736,N_634,N_1446);
nand U2737 (N_2737,N_209,N_430);
nor U2738 (N_2738,N_1233,N_127);
or U2739 (N_2739,N_624,N_965);
nand U2740 (N_2740,N_147,N_1426);
or U2741 (N_2741,N_1486,N_379);
nor U2742 (N_2742,N_1372,N_891);
or U2743 (N_2743,N_833,N_850);
or U2744 (N_2744,N_445,N_249);
or U2745 (N_2745,N_651,N_813);
or U2746 (N_2746,N_1157,N_1176);
and U2747 (N_2747,N_191,N_288);
and U2748 (N_2748,N_827,N_1007);
and U2749 (N_2749,N_667,N_1344);
xor U2750 (N_2750,N_464,N_1441);
and U2751 (N_2751,N_1345,N_522);
nor U2752 (N_2752,N_1106,N_520);
and U2753 (N_2753,N_585,N_44);
nor U2754 (N_2754,N_267,N_1410);
and U2755 (N_2755,N_575,N_1168);
nand U2756 (N_2756,N_553,N_159);
xnor U2757 (N_2757,N_91,N_44);
or U2758 (N_2758,N_1456,N_538);
xor U2759 (N_2759,N_478,N_647);
nand U2760 (N_2760,N_1124,N_888);
nor U2761 (N_2761,N_74,N_826);
and U2762 (N_2762,N_1123,N_1189);
or U2763 (N_2763,N_996,N_885);
or U2764 (N_2764,N_1267,N_1366);
xnor U2765 (N_2765,N_655,N_481);
nand U2766 (N_2766,N_1391,N_516);
nor U2767 (N_2767,N_774,N_787);
xor U2768 (N_2768,N_921,N_416);
and U2769 (N_2769,N_265,N_1011);
nor U2770 (N_2770,N_364,N_1151);
or U2771 (N_2771,N_414,N_407);
or U2772 (N_2772,N_1131,N_780);
nor U2773 (N_2773,N_241,N_1360);
xor U2774 (N_2774,N_1366,N_483);
nand U2775 (N_2775,N_957,N_1409);
nor U2776 (N_2776,N_475,N_836);
xor U2777 (N_2777,N_639,N_1029);
nand U2778 (N_2778,N_637,N_1479);
and U2779 (N_2779,N_52,N_400);
and U2780 (N_2780,N_1073,N_930);
nand U2781 (N_2781,N_1194,N_803);
xor U2782 (N_2782,N_213,N_1424);
nor U2783 (N_2783,N_453,N_59);
and U2784 (N_2784,N_209,N_1243);
nand U2785 (N_2785,N_213,N_829);
nor U2786 (N_2786,N_1400,N_1490);
nor U2787 (N_2787,N_1318,N_559);
and U2788 (N_2788,N_297,N_1305);
nand U2789 (N_2789,N_995,N_1197);
nor U2790 (N_2790,N_982,N_1119);
xor U2791 (N_2791,N_648,N_52);
or U2792 (N_2792,N_1351,N_1252);
and U2793 (N_2793,N_1486,N_1241);
nor U2794 (N_2794,N_563,N_550);
nand U2795 (N_2795,N_281,N_613);
nor U2796 (N_2796,N_153,N_421);
nor U2797 (N_2797,N_79,N_237);
and U2798 (N_2798,N_204,N_844);
xnor U2799 (N_2799,N_193,N_23);
and U2800 (N_2800,N_1094,N_1332);
xor U2801 (N_2801,N_893,N_161);
and U2802 (N_2802,N_1273,N_1296);
and U2803 (N_2803,N_609,N_493);
or U2804 (N_2804,N_801,N_711);
nor U2805 (N_2805,N_1081,N_890);
or U2806 (N_2806,N_1156,N_619);
xor U2807 (N_2807,N_721,N_917);
and U2808 (N_2808,N_895,N_399);
and U2809 (N_2809,N_728,N_1443);
and U2810 (N_2810,N_1165,N_1090);
or U2811 (N_2811,N_1048,N_13);
nor U2812 (N_2812,N_222,N_177);
nand U2813 (N_2813,N_1419,N_990);
xnor U2814 (N_2814,N_376,N_45);
and U2815 (N_2815,N_537,N_1436);
nor U2816 (N_2816,N_518,N_592);
nand U2817 (N_2817,N_388,N_1112);
nor U2818 (N_2818,N_63,N_1371);
nand U2819 (N_2819,N_411,N_1393);
or U2820 (N_2820,N_51,N_651);
nor U2821 (N_2821,N_612,N_275);
nor U2822 (N_2822,N_651,N_668);
nor U2823 (N_2823,N_1238,N_722);
or U2824 (N_2824,N_1305,N_182);
and U2825 (N_2825,N_102,N_193);
nor U2826 (N_2826,N_91,N_1487);
nand U2827 (N_2827,N_544,N_1175);
nand U2828 (N_2828,N_451,N_613);
nand U2829 (N_2829,N_1243,N_1208);
and U2830 (N_2830,N_143,N_244);
and U2831 (N_2831,N_289,N_1177);
or U2832 (N_2832,N_762,N_1210);
nand U2833 (N_2833,N_1134,N_438);
or U2834 (N_2834,N_718,N_533);
nand U2835 (N_2835,N_1425,N_650);
and U2836 (N_2836,N_1298,N_1082);
nand U2837 (N_2837,N_788,N_1390);
nand U2838 (N_2838,N_781,N_793);
and U2839 (N_2839,N_1056,N_608);
nor U2840 (N_2840,N_764,N_1244);
nor U2841 (N_2841,N_201,N_631);
xor U2842 (N_2842,N_1288,N_809);
nand U2843 (N_2843,N_653,N_134);
nand U2844 (N_2844,N_915,N_988);
or U2845 (N_2845,N_534,N_1469);
nor U2846 (N_2846,N_1388,N_532);
or U2847 (N_2847,N_902,N_1155);
nor U2848 (N_2848,N_425,N_755);
nand U2849 (N_2849,N_872,N_1447);
nand U2850 (N_2850,N_659,N_848);
xor U2851 (N_2851,N_294,N_724);
nor U2852 (N_2852,N_394,N_1045);
nand U2853 (N_2853,N_834,N_449);
or U2854 (N_2854,N_790,N_45);
nor U2855 (N_2855,N_1137,N_1306);
nand U2856 (N_2856,N_1299,N_841);
nand U2857 (N_2857,N_1458,N_432);
and U2858 (N_2858,N_384,N_585);
nand U2859 (N_2859,N_719,N_457);
xor U2860 (N_2860,N_712,N_971);
nand U2861 (N_2861,N_292,N_883);
xnor U2862 (N_2862,N_125,N_843);
nand U2863 (N_2863,N_972,N_99);
or U2864 (N_2864,N_378,N_677);
and U2865 (N_2865,N_1267,N_49);
nor U2866 (N_2866,N_718,N_1027);
nor U2867 (N_2867,N_117,N_950);
nand U2868 (N_2868,N_547,N_1140);
nor U2869 (N_2869,N_109,N_105);
or U2870 (N_2870,N_309,N_1130);
nor U2871 (N_2871,N_556,N_80);
nor U2872 (N_2872,N_351,N_544);
and U2873 (N_2873,N_909,N_1310);
nand U2874 (N_2874,N_1482,N_104);
or U2875 (N_2875,N_325,N_102);
or U2876 (N_2876,N_462,N_400);
xor U2877 (N_2877,N_646,N_275);
xor U2878 (N_2878,N_213,N_402);
and U2879 (N_2879,N_322,N_149);
or U2880 (N_2880,N_845,N_152);
nor U2881 (N_2881,N_676,N_728);
or U2882 (N_2882,N_933,N_1253);
and U2883 (N_2883,N_931,N_10);
nor U2884 (N_2884,N_99,N_484);
or U2885 (N_2885,N_818,N_711);
and U2886 (N_2886,N_1495,N_362);
and U2887 (N_2887,N_1064,N_858);
or U2888 (N_2888,N_204,N_1310);
nor U2889 (N_2889,N_1017,N_156);
or U2890 (N_2890,N_1274,N_1418);
nand U2891 (N_2891,N_158,N_328);
or U2892 (N_2892,N_37,N_777);
nand U2893 (N_2893,N_1164,N_577);
and U2894 (N_2894,N_165,N_826);
nand U2895 (N_2895,N_608,N_1200);
or U2896 (N_2896,N_584,N_599);
nand U2897 (N_2897,N_1003,N_490);
or U2898 (N_2898,N_282,N_287);
nor U2899 (N_2899,N_1368,N_1137);
nor U2900 (N_2900,N_60,N_654);
or U2901 (N_2901,N_1037,N_1083);
nand U2902 (N_2902,N_232,N_1147);
nor U2903 (N_2903,N_1160,N_796);
or U2904 (N_2904,N_1454,N_1443);
xor U2905 (N_2905,N_1045,N_88);
or U2906 (N_2906,N_1103,N_706);
xor U2907 (N_2907,N_1116,N_842);
nor U2908 (N_2908,N_105,N_882);
nor U2909 (N_2909,N_827,N_383);
or U2910 (N_2910,N_804,N_933);
nor U2911 (N_2911,N_356,N_1229);
nand U2912 (N_2912,N_225,N_1498);
nor U2913 (N_2913,N_1065,N_1240);
nand U2914 (N_2914,N_1257,N_724);
nand U2915 (N_2915,N_332,N_1282);
nor U2916 (N_2916,N_680,N_299);
and U2917 (N_2917,N_517,N_1499);
and U2918 (N_2918,N_1109,N_1213);
and U2919 (N_2919,N_1467,N_1107);
nand U2920 (N_2920,N_852,N_666);
nand U2921 (N_2921,N_459,N_63);
or U2922 (N_2922,N_1346,N_523);
nor U2923 (N_2923,N_794,N_207);
and U2924 (N_2924,N_1477,N_1007);
and U2925 (N_2925,N_227,N_799);
or U2926 (N_2926,N_1224,N_16);
nor U2927 (N_2927,N_818,N_1402);
or U2928 (N_2928,N_176,N_1327);
and U2929 (N_2929,N_1421,N_852);
nand U2930 (N_2930,N_47,N_765);
nor U2931 (N_2931,N_843,N_1428);
nand U2932 (N_2932,N_48,N_14);
or U2933 (N_2933,N_301,N_639);
xor U2934 (N_2934,N_1179,N_124);
xor U2935 (N_2935,N_1391,N_1251);
nor U2936 (N_2936,N_273,N_877);
or U2937 (N_2937,N_1031,N_1423);
nand U2938 (N_2938,N_452,N_1310);
or U2939 (N_2939,N_98,N_862);
and U2940 (N_2940,N_468,N_1022);
nand U2941 (N_2941,N_925,N_1150);
and U2942 (N_2942,N_1088,N_1423);
and U2943 (N_2943,N_1142,N_140);
and U2944 (N_2944,N_1363,N_902);
or U2945 (N_2945,N_1025,N_546);
nand U2946 (N_2946,N_65,N_932);
nand U2947 (N_2947,N_1243,N_1085);
or U2948 (N_2948,N_326,N_968);
and U2949 (N_2949,N_1490,N_561);
xor U2950 (N_2950,N_1490,N_546);
nor U2951 (N_2951,N_547,N_1330);
xor U2952 (N_2952,N_930,N_737);
nor U2953 (N_2953,N_1341,N_851);
or U2954 (N_2954,N_1356,N_1487);
and U2955 (N_2955,N_637,N_443);
nor U2956 (N_2956,N_863,N_688);
and U2957 (N_2957,N_1414,N_1241);
and U2958 (N_2958,N_1084,N_1143);
or U2959 (N_2959,N_419,N_1181);
nand U2960 (N_2960,N_823,N_1153);
xor U2961 (N_2961,N_515,N_119);
or U2962 (N_2962,N_264,N_1170);
nand U2963 (N_2963,N_813,N_509);
xor U2964 (N_2964,N_880,N_343);
or U2965 (N_2965,N_261,N_80);
xnor U2966 (N_2966,N_596,N_88);
and U2967 (N_2967,N_386,N_925);
xnor U2968 (N_2968,N_170,N_1253);
nand U2969 (N_2969,N_964,N_813);
and U2970 (N_2970,N_558,N_1448);
or U2971 (N_2971,N_1244,N_777);
and U2972 (N_2972,N_763,N_1459);
nand U2973 (N_2973,N_1371,N_1035);
nand U2974 (N_2974,N_529,N_560);
xnor U2975 (N_2975,N_431,N_103);
xor U2976 (N_2976,N_766,N_1114);
or U2977 (N_2977,N_550,N_506);
or U2978 (N_2978,N_924,N_723);
or U2979 (N_2979,N_1191,N_1445);
nand U2980 (N_2980,N_837,N_1076);
or U2981 (N_2981,N_404,N_989);
nor U2982 (N_2982,N_398,N_170);
nand U2983 (N_2983,N_846,N_1454);
nor U2984 (N_2984,N_574,N_1211);
nor U2985 (N_2985,N_860,N_377);
nand U2986 (N_2986,N_795,N_631);
xnor U2987 (N_2987,N_1246,N_711);
or U2988 (N_2988,N_276,N_407);
and U2989 (N_2989,N_711,N_1477);
nand U2990 (N_2990,N_94,N_801);
or U2991 (N_2991,N_156,N_1425);
nand U2992 (N_2992,N_1192,N_77);
nand U2993 (N_2993,N_334,N_1100);
or U2994 (N_2994,N_1175,N_189);
nor U2995 (N_2995,N_1397,N_213);
or U2996 (N_2996,N_964,N_1171);
nand U2997 (N_2997,N_654,N_221);
and U2998 (N_2998,N_749,N_518);
xnor U2999 (N_2999,N_750,N_831);
and U3000 (N_3000,N_2580,N_2655);
nand U3001 (N_3001,N_2960,N_2067);
nand U3002 (N_3002,N_2123,N_2853);
and U3003 (N_3003,N_2203,N_2750);
and U3004 (N_3004,N_2245,N_2847);
or U3005 (N_3005,N_1627,N_1568);
nand U3006 (N_3006,N_1621,N_2554);
or U3007 (N_3007,N_1565,N_1768);
and U3008 (N_3008,N_2332,N_2392);
xor U3009 (N_3009,N_2244,N_1828);
and U3010 (N_3010,N_2482,N_2294);
or U3011 (N_3011,N_2445,N_2219);
nor U3012 (N_3012,N_2072,N_1873);
nor U3013 (N_3013,N_2191,N_1574);
or U3014 (N_3014,N_2930,N_2721);
or U3015 (N_3015,N_2848,N_1556);
or U3016 (N_3016,N_2080,N_2794);
nand U3017 (N_3017,N_2417,N_1634);
nor U3018 (N_3018,N_1653,N_1876);
and U3019 (N_3019,N_2321,N_2555);
nor U3020 (N_3020,N_2405,N_1712);
nor U3021 (N_3021,N_1667,N_2034);
nor U3022 (N_3022,N_2697,N_1524);
and U3023 (N_3023,N_1808,N_1756);
or U3024 (N_3024,N_2193,N_2315);
xor U3025 (N_3025,N_1536,N_1723);
and U3026 (N_3026,N_2781,N_2556);
and U3027 (N_3027,N_2728,N_1571);
nor U3028 (N_3028,N_2419,N_1937);
or U3029 (N_3029,N_1933,N_2626);
nor U3030 (N_3030,N_2044,N_2524);
nand U3031 (N_3031,N_2987,N_2282);
and U3032 (N_3032,N_1930,N_2166);
or U3033 (N_3033,N_2999,N_2260);
or U3034 (N_3034,N_2346,N_1781);
and U3035 (N_3035,N_2873,N_2195);
or U3036 (N_3036,N_2364,N_2478);
or U3037 (N_3037,N_2688,N_2581);
xnor U3038 (N_3038,N_2114,N_1842);
nand U3039 (N_3039,N_2192,N_2661);
nor U3040 (N_3040,N_1977,N_2190);
or U3041 (N_3041,N_2276,N_2514);
or U3042 (N_3042,N_2906,N_2736);
or U3043 (N_3043,N_2559,N_2352);
nor U3044 (N_3044,N_2569,N_1841);
and U3045 (N_3045,N_2110,N_2523);
nand U3046 (N_3046,N_2942,N_2105);
nand U3047 (N_3047,N_1908,N_1917);
or U3048 (N_3048,N_2571,N_1913);
xor U3049 (N_3049,N_2570,N_2924);
nor U3050 (N_3050,N_2611,N_2917);
or U3051 (N_3051,N_2052,N_1533);
and U3052 (N_3052,N_1625,N_1793);
and U3053 (N_3053,N_2995,N_1965);
and U3054 (N_3054,N_1877,N_1978);
xnor U3055 (N_3055,N_1825,N_2603);
xor U3056 (N_3056,N_1949,N_2936);
nor U3057 (N_3057,N_2645,N_1865);
nand U3058 (N_3058,N_2639,N_2991);
or U3059 (N_3059,N_2837,N_2948);
and U3060 (N_3060,N_2888,N_1716);
or U3061 (N_3061,N_2117,N_2631);
or U3062 (N_3062,N_2345,N_1747);
nor U3063 (N_3063,N_2579,N_1845);
and U3064 (N_3064,N_1696,N_2983);
or U3065 (N_3065,N_1889,N_1948);
and U3066 (N_3066,N_2157,N_2535);
or U3067 (N_3067,N_2823,N_2015);
nand U3068 (N_3068,N_2164,N_2676);
and U3069 (N_3069,N_2553,N_1931);
nand U3070 (N_3070,N_2507,N_2012);
or U3071 (N_3071,N_2429,N_2693);
nor U3072 (N_3072,N_2214,N_2342);
and U3073 (N_3073,N_2746,N_2996);
and U3074 (N_3074,N_2258,N_2143);
and U3075 (N_3075,N_2934,N_1882);
xnor U3076 (N_3076,N_2589,N_2098);
and U3077 (N_3077,N_2437,N_2869);
xor U3078 (N_3078,N_1671,N_2825);
nor U3079 (N_3079,N_1740,N_1640);
or U3080 (N_3080,N_1534,N_2403);
nand U3081 (N_3081,N_1733,N_2367);
and U3082 (N_3082,N_1602,N_2501);
nand U3083 (N_3083,N_1817,N_2247);
nand U3084 (N_3084,N_2707,N_2412);
and U3085 (N_3085,N_2544,N_2174);
nor U3086 (N_3086,N_2469,N_2726);
or U3087 (N_3087,N_2327,N_1871);
or U3088 (N_3088,N_2777,N_1938);
nand U3089 (N_3089,N_2086,N_2551);
nand U3090 (N_3090,N_2701,N_2497);
nand U3091 (N_3091,N_2729,N_2747);
and U3092 (N_3092,N_2604,N_1720);
nor U3093 (N_3093,N_1604,N_2939);
or U3094 (N_3094,N_1707,N_2209);
xnor U3095 (N_3095,N_1951,N_2703);
or U3096 (N_3096,N_1827,N_2952);
nor U3097 (N_3097,N_2973,N_2118);
nor U3098 (N_3098,N_2962,N_2685);
nor U3099 (N_3099,N_2040,N_2138);
or U3100 (N_3100,N_2454,N_2243);
nor U3101 (N_3101,N_2949,N_2055);
or U3102 (N_3102,N_1867,N_2019);
and U3103 (N_3103,N_1771,N_2031);
and U3104 (N_3104,N_2162,N_2986);
or U3105 (N_3105,N_2719,N_2388);
and U3106 (N_3106,N_2880,N_1940);
nand U3107 (N_3107,N_1925,N_1862);
or U3108 (N_3108,N_2439,N_2511);
or U3109 (N_3109,N_2773,N_2593);
nor U3110 (N_3110,N_2966,N_2506);
nand U3111 (N_3111,N_2222,N_2199);
nor U3112 (N_3112,N_1963,N_1750);
nor U3113 (N_3113,N_1852,N_1584);
and U3114 (N_3114,N_2850,N_2672);
and U3115 (N_3115,N_2979,N_2187);
nand U3116 (N_3116,N_1582,N_2749);
xnor U3117 (N_3117,N_2623,N_2084);
or U3118 (N_3118,N_2740,N_1754);
and U3119 (N_3119,N_1958,N_1526);
or U3120 (N_3120,N_2334,N_2664);
nor U3121 (N_3121,N_2009,N_2254);
or U3122 (N_3122,N_2658,N_2329);
and U3123 (N_3123,N_1911,N_2517);
xor U3124 (N_3124,N_2763,N_1893);
xnor U3125 (N_3125,N_1885,N_2834);
or U3126 (N_3126,N_1714,N_2430);
xnor U3127 (N_3127,N_2933,N_1559);
nand U3128 (N_3128,N_1833,N_2421);
and U3129 (N_3129,N_2946,N_2543);
xor U3130 (N_3130,N_2566,N_2365);
nor U3131 (N_3131,N_2499,N_1548);
nor U3132 (N_3132,N_2588,N_1799);
nand U3133 (N_3133,N_2826,N_2992);
nor U3134 (N_3134,N_1655,N_1832);
and U3135 (N_3135,N_1941,N_2185);
nor U3136 (N_3136,N_2926,N_1765);
and U3137 (N_3137,N_1989,N_2742);
or U3138 (N_3138,N_2680,N_2592);
nor U3139 (N_3139,N_2899,N_2638);
nand U3140 (N_3140,N_2265,N_1736);
and U3141 (N_3141,N_2753,N_2378);
xnor U3142 (N_3142,N_2882,N_1731);
or U3143 (N_3143,N_1920,N_2331);
nor U3144 (N_3144,N_2622,N_2158);
nand U3145 (N_3145,N_1557,N_2512);
xnor U3146 (N_3146,N_1957,N_2852);
nor U3147 (N_3147,N_2301,N_2528);
or U3148 (N_3148,N_2272,N_1814);
or U3149 (N_3149,N_1767,N_2772);
or U3150 (N_3150,N_1670,N_2024);
xnor U3151 (N_3151,N_2408,N_1848);
xnor U3152 (N_3152,N_2700,N_2017);
xnor U3153 (N_3153,N_2738,N_1981);
xor U3154 (N_3154,N_1947,N_2359);
nor U3155 (N_3155,N_2951,N_2128);
and U3156 (N_3156,N_1878,N_1782);
nand U3157 (N_3157,N_2731,N_2010);
nor U3158 (N_3158,N_2835,N_2533);
nor U3159 (N_3159,N_2165,N_2217);
xor U3160 (N_3160,N_1753,N_2255);
or U3161 (N_3161,N_1902,N_2238);
and U3162 (N_3162,N_2771,N_1821);
nand U3163 (N_3163,N_1628,N_2994);
and U3164 (N_3164,N_2526,N_2855);
or U3165 (N_3165,N_1928,N_2950);
nand U3166 (N_3166,N_2928,N_1773);
nor U3167 (N_3167,N_2197,N_2653);
xor U3168 (N_3168,N_1899,N_2093);
and U3169 (N_3169,N_2168,N_2492);
nor U3170 (N_3170,N_2572,N_2167);
or U3171 (N_3171,N_2038,N_2971);
nand U3172 (N_3172,N_2896,N_2250);
and U3173 (N_3173,N_1744,N_2505);
and U3174 (N_3174,N_2790,N_1769);
xor U3175 (N_3175,N_1783,N_1503);
or U3176 (N_3176,N_1974,N_2328);
nand U3177 (N_3177,N_1554,N_2586);
or U3178 (N_3178,N_1792,N_2576);
nor U3179 (N_3179,N_2182,N_2762);
or U3180 (N_3180,N_2377,N_1863);
nand U3181 (N_3181,N_1500,N_2807);
and U3182 (N_3182,N_1538,N_2865);
and U3183 (N_3183,N_2273,N_2641);
nor U3184 (N_3184,N_2479,N_2060);
nand U3185 (N_3185,N_2938,N_1654);
nand U3186 (N_3186,N_2724,N_1504);
or U3187 (N_3187,N_1727,N_2633);
or U3188 (N_3188,N_2816,N_2562);
nand U3189 (N_3189,N_2560,N_2287);
nor U3190 (N_3190,N_1562,N_1729);
and U3191 (N_3191,N_1607,N_2299);
nand U3192 (N_3192,N_2978,N_2532);
and U3193 (N_3193,N_1570,N_1888);
and U3194 (N_3194,N_2385,N_2285);
nand U3195 (N_3195,N_2401,N_2904);
or U3196 (N_3196,N_1830,N_1519);
nor U3197 (N_3197,N_2764,N_1718);
nand U3198 (N_3198,N_2754,N_1674);
xnor U3199 (N_3199,N_2616,N_2253);
or U3200 (N_3200,N_2968,N_2413);
nand U3201 (N_3201,N_1966,N_1944);
nor U3202 (N_3202,N_2360,N_2522);
nor U3203 (N_3203,N_2822,N_1587);
nor U3204 (N_3204,N_2607,N_2223);
or U3205 (N_3205,N_1840,N_2643);
nor U3206 (N_3206,N_2748,N_2220);
or U3207 (N_3207,N_1900,N_2859);
and U3208 (N_3208,N_2129,N_2974);
or U3209 (N_3209,N_1804,N_2884);
nor U3210 (N_3210,N_2844,N_2760);
and U3211 (N_3211,N_1800,N_1796);
or U3212 (N_3212,N_2494,N_1954);
or U3213 (N_3213,N_2268,N_1872);
nor U3214 (N_3214,N_2001,N_1521);
and U3215 (N_3215,N_2775,N_2887);
or U3216 (N_3216,N_1527,N_2786);
and U3217 (N_3217,N_2022,N_2070);
and U3218 (N_3218,N_2830,N_1778);
nor U3219 (N_3219,N_1818,N_2390);
nor U3220 (N_3220,N_2186,N_1580);
nand U3221 (N_3221,N_2350,N_2737);
nand U3222 (N_3222,N_2860,N_1860);
and U3223 (N_3223,N_1995,N_2879);
nand U3224 (N_3224,N_2578,N_2625);
nand U3225 (N_3225,N_1505,N_2043);
and U3226 (N_3226,N_1757,N_2281);
nand U3227 (N_3227,N_2539,N_2183);
xor U3228 (N_3228,N_2997,N_2954);
nand U3229 (N_3229,N_2805,N_2296);
or U3230 (N_3230,N_2196,N_2127);
nor U3231 (N_3231,N_2251,N_2373);
or U3232 (N_3232,N_2911,N_1886);
nor U3233 (N_3233,N_2319,N_2689);
nor U3234 (N_3234,N_2446,N_1784);
or U3235 (N_3235,N_2406,N_2915);
or U3236 (N_3236,N_2587,N_2914);
nand U3237 (N_3237,N_2466,N_1780);
xor U3238 (N_3238,N_1575,N_2139);
and U3239 (N_3239,N_1589,N_1661);
and U3240 (N_3240,N_2263,N_1598);
or U3241 (N_3241,N_2756,N_2134);
nor U3242 (N_3242,N_1766,N_2515);
or U3243 (N_3243,N_1857,N_2003);
nor U3244 (N_3244,N_2177,N_2104);
nand U3245 (N_3245,N_1528,N_2574);
nand U3246 (N_3246,N_1846,N_1961);
and U3247 (N_3247,N_2504,N_2142);
nand U3248 (N_3248,N_2152,N_2665);
and U3249 (N_3249,N_1724,N_1647);
and U3250 (N_3250,N_1578,N_1529);
or U3251 (N_3251,N_1903,N_1969);
and U3252 (N_3252,N_2155,N_2008);
and U3253 (N_3253,N_1929,N_2916);
nand U3254 (N_3254,N_2567,N_2344);
or U3255 (N_3255,N_2023,N_2905);
nand U3256 (N_3256,N_2782,N_1824);
nand U3257 (N_3257,N_2932,N_2981);
and U3258 (N_3258,N_1983,N_2881);
xor U3259 (N_3259,N_2982,N_2006);
and U3260 (N_3260,N_2690,N_1708);
nor U3261 (N_3261,N_1685,N_2371);
and U3262 (N_3262,N_1612,N_2460);
xor U3263 (N_3263,N_2189,N_2313);
and U3264 (N_3264,N_2351,N_2298);
and U3265 (N_3265,N_2425,N_2411);
nor U3266 (N_3266,N_2343,N_2767);
or U3267 (N_3267,N_1650,N_1638);
nand U3268 (N_3268,N_2037,N_2065);
nand U3269 (N_3269,N_2242,N_2005);
and U3270 (N_3270,N_2297,N_2396);
nor U3271 (N_3271,N_1516,N_1682);
nand U3272 (N_3272,N_1703,N_2096);
and U3273 (N_3273,N_2550,N_1734);
nor U3274 (N_3274,N_2434,N_2119);
and U3275 (N_3275,N_1525,N_2366);
or U3276 (N_3276,N_2667,N_2317);
nand U3277 (N_3277,N_2797,N_1791);
nor U3278 (N_3278,N_2453,N_1764);
and U3279 (N_3279,N_2670,N_2613);
and U3280 (N_3280,N_2941,N_2325);
nand U3281 (N_3281,N_1721,N_1681);
or U3282 (N_3282,N_1763,N_1659);
and U3283 (N_3283,N_1918,N_2462);
xor U3284 (N_3284,N_1835,N_2036);
and U3285 (N_3285,N_2432,N_1728);
nand U3286 (N_3286,N_2374,N_2259);
and U3287 (N_3287,N_1633,N_2791);
xnor U3288 (N_3288,N_1919,N_2277);
nand U3289 (N_3289,N_2868,N_2799);
xnor U3290 (N_3290,N_2789,N_2481);
or U3291 (N_3291,N_2839,N_2370);
nor U3292 (N_3292,N_2629,N_2452);
and U3293 (N_3293,N_2358,N_2500);
or U3294 (N_3294,N_2663,N_2598);
nor U3295 (N_3295,N_2188,N_1851);
nor U3296 (N_3296,N_2041,N_1770);
nand U3297 (N_3297,N_1749,N_2221);
nor U3298 (N_3298,N_2796,N_2180);
or U3299 (N_3299,N_2969,N_2929);
nand U3300 (N_3300,N_2699,N_1709);
or U3301 (N_3301,N_1615,N_2422);
or U3302 (N_3302,N_1591,N_2078);
or U3303 (N_3303,N_2716,N_2648);
nor U3304 (N_3304,N_2402,N_2326);
or U3305 (N_3305,N_2234,N_2475);
nand U3306 (N_3306,N_2606,N_1993);
and U3307 (N_3307,N_2488,N_2957);
nand U3308 (N_3308,N_2461,N_2675);
nand U3309 (N_3309,N_2780,N_2092);
xor U3310 (N_3310,N_2692,N_2863);
and U3311 (N_3311,N_2669,N_2521);
and U3312 (N_3312,N_2210,N_2278);
and U3313 (N_3313,N_1583,N_2115);
xnor U3314 (N_3314,N_2262,N_2459);
nor U3315 (N_3315,N_1547,N_2980);
and U3316 (N_3316,N_1713,N_2708);
or U3317 (N_3317,N_2927,N_2922);
xor U3318 (N_3318,N_2711,N_2901);
or U3319 (N_3319,N_2668,N_2612);
nand U3320 (N_3320,N_2102,N_2829);
nor U3321 (N_3321,N_2101,N_2694);
nor U3322 (N_3322,N_1738,N_2050);
xnor U3323 (N_3323,N_1997,N_1572);
or U3324 (N_3324,N_1946,N_2947);
or U3325 (N_3325,N_2564,N_1774);
nor U3326 (N_3326,N_2495,N_2069);
nand U3327 (N_3327,N_1614,N_2943);
nor U3328 (N_3328,N_2503,N_2874);
or U3329 (N_3329,N_1502,N_2998);
and U3330 (N_3330,N_1785,N_2380);
and U3331 (N_3331,N_2919,N_2279);
or U3332 (N_3332,N_1646,N_1866);
or U3333 (N_3333,N_2091,N_1610);
or U3334 (N_3334,N_2845,N_2473);
and U3335 (N_3335,N_1758,N_1535);
and U3336 (N_3336,N_1699,N_2843);
or U3337 (N_3337,N_2801,N_2369);
xnor U3338 (N_3338,N_2988,N_2135);
nand U3339 (N_3339,N_1726,N_1912);
xor U3340 (N_3340,N_2318,N_2290);
nor U3341 (N_3341,N_2608,N_2449);
xor U3342 (N_3342,N_2609,N_2745);
nor U3343 (N_3343,N_2307,N_2389);
nand U3344 (N_3344,N_1829,N_2382);
nor U3345 (N_3345,N_2071,N_1869);
nand U3346 (N_3346,N_1677,N_2508);
nor U3347 (N_3347,N_2025,N_1856);
nand U3348 (N_3348,N_1854,N_2595);
or U3349 (N_3349,N_2051,N_1987);
xnor U3350 (N_3350,N_1636,N_1904);
and U3351 (N_3351,N_2650,N_1608);
and U3352 (N_3352,N_1960,N_2150);
and U3353 (N_3353,N_2516,N_1711);
or U3354 (N_3354,N_2121,N_2891);
or U3355 (N_3355,N_2246,N_2619);
nor U3356 (N_3356,N_2838,N_2621);
nand U3357 (N_3357,N_2858,N_2815);
xnor U3358 (N_3358,N_1551,N_2467);
nand U3359 (N_3359,N_2458,N_2596);
and U3360 (N_3360,N_2103,N_1581);
or U3361 (N_3361,N_2184,N_1596);
nand U3362 (N_3362,N_2484,N_2083);
and U3363 (N_3363,N_1879,N_2678);
or U3364 (N_3364,N_2889,N_2818);
or U3365 (N_3365,N_2696,N_1595);
nor U3366 (N_3366,N_2733,N_1843);
nor U3367 (N_3367,N_1520,N_2575);
or U3368 (N_3368,N_1849,N_2540);
nand U3369 (N_3369,N_1701,N_1988);
nor U3370 (N_3370,N_2683,N_2026);
nor U3371 (N_3371,N_2033,N_2964);
and U3372 (N_3372,N_2257,N_2148);
nand U3373 (N_3373,N_2302,N_2176);
and U3374 (N_3374,N_2885,N_1950);
and U3375 (N_3375,N_2443,N_2206);
or U3376 (N_3376,N_2269,N_1805);
nand U3377 (N_3377,N_2339,N_2379);
or U3378 (N_3378,N_2963,N_1510);
and U3379 (N_3379,N_1730,N_2125);
and U3380 (N_3380,N_2679,N_2151);
or U3381 (N_3381,N_2248,N_2832);
nand U3382 (N_3382,N_1819,N_2349);
nand U3383 (N_3383,N_2907,N_1868);
nand U3384 (N_3384,N_1923,N_2857);
nor U3385 (N_3385,N_1586,N_2627);
nand U3386 (N_3386,N_2886,N_2491);
nor U3387 (N_3387,N_2471,N_1555);
and U3388 (N_3388,N_1656,N_2940);
nand U3389 (N_3389,N_2984,N_2013);
xnor U3390 (N_3390,N_2831,N_2713);
or U3391 (N_3391,N_2061,N_1725);
or U3392 (N_3392,N_2862,N_1537);
and U3393 (N_3393,N_2827,N_2808);
nor U3394 (N_3394,N_2144,N_1898);
nand U3395 (N_3395,N_2893,N_1984);
xor U3396 (N_3396,N_2836,N_2386);
or U3397 (N_3397,N_2787,N_1921);
and U3398 (N_3398,N_2741,N_2636);
or U3399 (N_3399,N_2635,N_2486);
nand U3400 (N_3400,N_2252,N_2876);
nor U3401 (N_3401,N_2323,N_2909);
or U3402 (N_3402,N_2730,N_2531);
and U3403 (N_3403,N_2046,N_2178);
and U3404 (N_3404,N_2424,N_2136);
nand U3405 (N_3405,N_2106,N_1687);
nor U3406 (N_3406,N_1569,N_2181);
nor U3407 (N_3407,N_2237,N_2368);
or U3408 (N_3408,N_2732,N_2601);
and U3409 (N_3409,N_1660,N_2856);
and U3410 (N_3410,N_1657,N_1890);
nand U3411 (N_3411,N_1970,N_2153);
xor U3412 (N_3412,N_1952,N_2356);
or U3413 (N_3413,N_1775,N_2039);
xnor U3414 (N_3414,N_2903,N_2520);
nor U3415 (N_3415,N_1684,N_2451);
and U3416 (N_3416,N_2878,N_2241);
nor U3417 (N_3417,N_1705,N_2225);
nor U3418 (N_3418,N_2718,N_2147);
or U3419 (N_3419,N_2124,N_2362);
or U3420 (N_3420,N_2493,N_1892);
or U3421 (N_3421,N_2892,N_2415);
and U3422 (N_3422,N_1838,N_1509);
or U3423 (N_3423,N_1539,N_1915);
nor U3424 (N_3424,N_1870,N_1563);
nor U3425 (N_3425,N_2972,N_2811);
nor U3426 (N_3426,N_1560,N_2045);
and U3427 (N_3427,N_2720,N_2058);
or U3428 (N_3428,N_1884,N_2530);
nor U3429 (N_3429,N_2812,N_1579);
or U3430 (N_3430,N_2759,N_1801);
nand U3431 (N_3431,N_1910,N_2602);
and U3432 (N_3432,N_2082,N_1577);
xor U3433 (N_3433,N_2854,N_2375);
nand U3434 (N_3434,N_1609,N_2057);
nor U3435 (N_3435,N_2895,N_2931);
or U3436 (N_3436,N_1945,N_2229);
and U3437 (N_3437,N_2310,N_1629);
nand U3438 (N_3438,N_2198,N_2712);
nand U3439 (N_3439,N_2813,N_2545);
nand U3440 (N_3440,N_1979,N_2099);
or U3441 (N_3441,N_2624,N_2549);
and U3442 (N_3442,N_1992,N_2395);
and U3443 (N_3443,N_1619,N_1743);
nand U3444 (N_3444,N_2646,N_1968);
nand U3445 (N_3445,N_2722,N_2537);
nor U3446 (N_3446,N_2630,N_2097);
nand U3447 (N_3447,N_2561,N_2894);
nor U3448 (N_3448,N_2577,N_2803);
nor U3449 (N_3449,N_2457,N_2814);
and U3450 (N_3450,N_2605,N_2674);
xnor U3451 (N_3451,N_1875,N_2075);
nor U3452 (N_3452,N_2267,N_2849);
and U3453 (N_3453,N_2765,N_2944);
nor U3454 (N_3454,N_2824,N_1901);
nand U3455 (N_3455,N_2049,N_1518);
xor U3456 (N_3456,N_2841,N_1996);
nor U3457 (N_3457,N_1861,N_2029);
nand U3458 (N_3458,N_1552,N_2465);
nor U3459 (N_3459,N_2109,N_2656);
nand U3460 (N_3460,N_1932,N_2074);
nor U3461 (N_3461,N_2387,N_1956);
and U3462 (N_3462,N_2231,N_1816);
and U3463 (N_3463,N_2383,N_2935);
and U3464 (N_3464,N_2160,N_1651);
or U3465 (N_3465,N_2568,N_2095);
xnor U3466 (N_3466,N_2977,N_2734);
nor U3467 (N_3467,N_2354,N_2890);
or U3468 (N_3468,N_2681,N_2447);
xnor U3469 (N_3469,N_1745,N_2582);
nor U3470 (N_3470,N_1632,N_1501);
or U3471 (N_3471,N_2428,N_1786);
or U3472 (N_3472,N_2423,N_2802);
nand U3473 (N_3473,N_2710,N_2840);
and U3474 (N_3474,N_1822,N_2751);
nand U3475 (N_3475,N_1836,N_2766);
nor U3476 (N_3476,N_1611,N_2291);
or U3477 (N_3477,N_2000,N_2032);
xor U3478 (N_3478,N_2207,N_1722);
xor U3479 (N_3479,N_1673,N_2918);
xor U3480 (N_3480,N_2666,N_1982);
or U3481 (N_3481,N_1631,N_2438);
xor U3482 (N_3482,N_2793,N_1916);
nand U3483 (N_3483,N_1688,N_2961);
and U3484 (N_3484,N_2806,N_2476);
and U3485 (N_3485,N_1760,N_1517);
or U3486 (N_3486,N_2159,N_2776);
and U3487 (N_3487,N_2081,N_2020);
or U3488 (N_3488,N_1588,N_2691);
or U3489 (N_3489,N_2394,N_2867);
or U3490 (N_3490,N_1967,N_2361);
or U3491 (N_3491,N_2662,N_1752);
nor U3492 (N_3492,N_1939,N_1839);
nand U3493 (N_3493,N_1797,N_1522);
and U3494 (N_3494,N_2615,N_2035);
nor U3495 (N_3495,N_2322,N_1635);
or U3496 (N_3496,N_1823,N_2030);
nand U3497 (N_3497,N_2308,N_1737);
nand U3498 (N_3498,N_2498,N_1812);
nand U3499 (N_3499,N_2739,N_2558);
or U3500 (N_3500,N_2100,N_1543);
and U3501 (N_3501,N_2011,N_2068);
and U3502 (N_3502,N_2088,N_1689);
or U3503 (N_3503,N_2817,N_2913);
or U3504 (N_3504,N_1742,N_2620);
and U3505 (N_3505,N_2054,N_1959);
nor U3506 (N_3506,N_2464,N_2420);
nor U3507 (N_3507,N_1593,N_2064);
or U3508 (N_3508,N_2427,N_1626);
or U3509 (N_3509,N_1666,N_1662);
and U3510 (N_3510,N_2407,N_1592);
or U3511 (N_3511,N_2218,N_2594);
nand U3512 (N_3512,N_1623,N_2821);
nor U3513 (N_3513,N_2965,N_2795);
xor U3514 (N_3514,N_2284,N_2744);
nand U3515 (N_3515,N_2779,N_2264);
nor U3516 (N_3516,N_2122,N_2959);
and U3517 (N_3517,N_2270,N_2489);
nand U3518 (N_3518,N_1735,N_2442);
and U3519 (N_3519,N_1693,N_1924);
nand U3520 (N_3520,N_1844,N_1971);
or U3521 (N_3521,N_1594,N_2912);
nor U3522 (N_3522,N_2792,N_2833);
or U3523 (N_3523,N_1532,N_1649);
nand U3524 (N_3524,N_2784,N_1855);
or U3525 (N_3525,N_2444,N_2659);
or U3526 (N_3526,N_2213,N_1972);
nor U3527 (N_3527,N_2426,N_2513);
and U3528 (N_3528,N_2953,N_2757);
or U3529 (N_3529,N_2141,N_2698);
and U3530 (N_3530,N_2431,N_2752);
or U3531 (N_3531,N_2585,N_2706);
or U3532 (N_3532,N_2416,N_2463);
nand U3533 (N_3533,N_2227,N_2989);
xor U3534 (N_3534,N_2778,N_2557);
nand U3535 (N_3535,N_2519,N_2363);
or U3536 (N_3536,N_1664,N_2133);
or U3537 (N_3537,N_2470,N_1759);
nor U3538 (N_3538,N_2314,N_1942);
nor U3539 (N_3539,N_2975,N_2695);
or U3540 (N_3540,N_2172,N_2487);
and U3541 (N_3541,N_2861,N_2509);
nand U3542 (N_3542,N_2063,N_2376);
nand U3543 (N_3543,N_2477,N_2534);
nor U3544 (N_3544,N_1700,N_2089);
nor U3545 (N_3545,N_2384,N_2723);
and U3546 (N_3546,N_2714,N_2283);
nor U3547 (N_3547,N_1648,N_2970);
and U3548 (N_3548,N_1934,N_2870);
nor U3549 (N_3549,N_2156,N_2316);
or U3550 (N_3550,N_2640,N_2048);
nand U3551 (N_3551,N_1544,N_2800);
xor U3552 (N_3552,N_2085,N_2654);
nand U3553 (N_3553,N_1909,N_2820);
or U3554 (N_3554,N_2145,N_2357);
nor U3555 (N_3555,N_2336,N_1605);
or U3556 (N_3556,N_1698,N_1906);
nand U3557 (N_3557,N_2783,N_2923);
and U3558 (N_3558,N_2021,N_1507);
or U3559 (N_3559,N_1999,N_2169);
nand U3560 (N_3560,N_2875,N_2397);
and U3561 (N_3561,N_2435,N_1834);
xnor U3562 (N_3562,N_2016,N_1837);
or U3563 (N_3563,N_1567,N_2441);
and U3564 (N_3564,N_2686,N_2275);
nor U3565 (N_3565,N_1601,N_2330);
or U3566 (N_3566,N_1788,N_2483);
and U3567 (N_3567,N_2341,N_2404);
and U3568 (N_3568,N_2565,N_2236);
and U3569 (N_3569,N_2828,N_2200);
and U3570 (N_3570,N_1669,N_2400);
nand U3571 (N_3571,N_1665,N_2090);
nor U3572 (N_3572,N_2684,N_1746);
and U3573 (N_3573,N_2637,N_2717);
xor U3574 (N_3574,N_2230,N_2014);
nor U3575 (N_3575,N_2902,N_1576);
or U3576 (N_3576,N_2925,N_2958);
nand U3577 (N_3577,N_1810,N_2705);
and U3578 (N_3578,N_1645,N_1973);
nor U3579 (N_3579,N_2455,N_2062);
or U3580 (N_3580,N_2130,N_1513);
xor U3581 (N_3581,N_2107,N_2274);
nor U3582 (N_3582,N_2266,N_1617);
nor U3583 (N_3583,N_2340,N_1694);
nor U3584 (N_3584,N_1620,N_2306);
nor U3585 (N_3585,N_2956,N_2614);
and U3586 (N_3586,N_2398,N_2338);
and U3587 (N_3587,N_2304,N_1881);
nand U3588 (N_3588,N_2399,N_2450);
and U3589 (N_3589,N_2215,N_1630);
nor U3590 (N_3590,N_1642,N_2126);
and U3591 (N_3591,N_2921,N_2216);
and U3592 (N_3592,N_2937,N_1643);
or U3593 (N_3593,N_2146,N_2440);
and U3594 (N_3594,N_2866,N_2414);
or U3595 (N_3595,N_2908,N_1603);
nor U3596 (N_3596,N_1658,N_2502);
nand U3597 (N_3597,N_1732,N_1523);
xnor U3598 (N_3598,N_2094,N_1772);
and U3599 (N_3599,N_1964,N_2249);
nand U3600 (N_3600,N_2320,N_2496);
or U3601 (N_3601,N_2289,N_1779);
and U3602 (N_3602,N_1820,N_2955);
nand U3603 (N_3603,N_2804,N_1678);
xor U3604 (N_3604,N_1706,N_2324);
nand U3605 (N_3605,N_2239,N_2743);
xnor U3606 (N_3606,N_2468,N_2293);
nand U3607 (N_3607,N_1686,N_2599);
nand U3608 (N_3608,N_2271,N_1692);
and U3609 (N_3609,N_2212,N_2993);
nor U3610 (N_3610,N_1540,N_1787);
nand U3611 (N_3611,N_2704,N_1585);
or U3612 (N_3612,N_2518,N_2671);
nor U3613 (N_3613,N_2073,N_2552);
or U3614 (N_3614,N_1719,N_2525);
nand U3615 (N_3615,N_2007,N_2233);
nor U3616 (N_3616,N_1790,N_2788);
nand U3617 (N_3617,N_2644,N_2632);
nand U3618 (N_3618,N_2657,N_2353);
nand U3619 (N_3619,N_2727,N_2131);
xnor U3620 (N_3620,N_1795,N_2967);
and U3621 (N_3621,N_1717,N_1546);
xnor U3622 (N_3622,N_1896,N_1874);
and U3623 (N_3623,N_2261,N_2175);
nor U3624 (N_3624,N_1809,N_2920);
or U3625 (N_3625,N_2642,N_1695);
nor U3626 (N_3626,N_1541,N_2137);
or U3627 (N_3627,N_2111,N_2303);
or U3628 (N_3628,N_2288,N_1530);
nand U3629 (N_3629,N_1690,N_2018);
xnor U3630 (N_3630,N_1755,N_2682);
nand U3631 (N_3631,N_2056,N_1624);
and U3632 (N_3632,N_1789,N_1613);
or U3633 (N_3633,N_1922,N_1675);
nand U3634 (N_3634,N_2652,N_2161);
nand U3635 (N_3635,N_1710,N_2785);
or U3636 (N_3636,N_1663,N_2179);
or U3637 (N_3637,N_1762,N_1858);
nor U3638 (N_3638,N_2409,N_2112);
nor U3639 (N_3639,N_2774,N_2347);
and U3640 (N_3640,N_1887,N_1561);
and U3641 (N_3641,N_1798,N_1751);
and U3642 (N_3642,N_1803,N_2871);
or U3643 (N_3643,N_2898,N_2809);
xnor U3644 (N_3644,N_1776,N_2610);
xor U3645 (N_3645,N_1927,N_2563);
or U3646 (N_3646,N_2660,N_1990);
nand U3647 (N_3647,N_2042,N_2224);
xnor U3648 (N_3648,N_2597,N_2628);
or U3649 (N_3649,N_1545,N_1986);
nor U3650 (N_3650,N_2132,N_1511);
nand U3651 (N_3651,N_1506,N_2583);
and U3652 (N_3652,N_1715,N_1668);
and U3653 (N_3653,N_1597,N_2677);
nor U3654 (N_3654,N_2077,N_1531);
and U3655 (N_3655,N_1553,N_2295);
and U3656 (N_3656,N_2333,N_1905);
or U3657 (N_3657,N_1691,N_1618);
or U3658 (N_3658,N_2702,N_2002);
nand U3659 (N_3659,N_2116,N_1697);
or U3660 (N_3660,N_2590,N_2715);
nor U3661 (N_3661,N_2761,N_2312);
or U3662 (N_3662,N_1550,N_2538);
and U3663 (N_3663,N_2755,N_2649);
or U3664 (N_3664,N_2573,N_2810);
or U3665 (N_3665,N_2309,N_1549);
nand U3666 (N_3666,N_1826,N_2226);
xor U3667 (N_3667,N_2735,N_2546);
and U3668 (N_3668,N_1975,N_1761);
xor U3669 (N_3669,N_2900,N_2300);
and U3670 (N_3670,N_2154,N_2536);
and U3671 (N_3671,N_1652,N_1616);
and U3672 (N_3672,N_2170,N_1641);
nand U3673 (N_3673,N_2171,N_1883);
nand U3674 (N_3674,N_2617,N_1813);
or U3675 (N_3675,N_2510,N_1639);
or U3676 (N_3676,N_1847,N_2240);
xnor U3677 (N_3677,N_2201,N_2108);
xor U3678 (N_3678,N_1622,N_2851);
or U3679 (N_3679,N_2348,N_2842);
nor U3680 (N_3680,N_2337,N_2618);
and U3681 (N_3681,N_2864,N_1566);
xnor U3682 (N_3682,N_2391,N_1564);
nor U3683 (N_3683,N_1683,N_2600);
nand U3684 (N_3684,N_2798,N_2472);
nor U3685 (N_3685,N_1953,N_1998);
nor U3686 (N_3686,N_2372,N_2204);
nor U3687 (N_3687,N_2945,N_2819);
or U3688 (N_3688,N_2872,N_2027);
and U3689 (N_3689,N_1590,N_2990);
nand U3690 (N_3690,N_2490,N_2355);
nand U3691 (N_3691,N_2768,N_2381);
and U3692 (N_3692,N_2066,N_1991);
or U3693 (N_3693,N_2211,N_1955);
xor U3694 (N_3694,N_2292,N_1514);
nor U3695 (N_3695,N_2311,N_2541);
nand U3696 (N_3696,N_2173,N_1815);
and U3697 (N_3697,N_2436,N_1508);
and U3698 (N_3698,N_2228,N_2456);
xnor U3699 (N_3699,N_2004,N_2205);
nor U3700 (N_3700,N_1739,N_2547);
or U3701 (N_3701,N_2673,N_1806);
nor U3702 (N_3702,N_1600,N_2877);
nor U3703 (N_3703,N_2897,N_1976);
nor U3704 (N_3704,N_2529,N_1891);
nand U3705 (N_3705,N_1811,N_2113);
nor U3706 (N_3706,N_1985,N_1914);
and U3707 (N_3707,N_1573,N_2256);
or U3708 (N_3708,N_1512,N_2758);
or U3709 (N_3709,N_1672,N_2709);
or U3710 (N_3710,N_2053,N_2591);
nor U3711 (N_3711,N_2140,N_1962);
or U3712 (N_3712,N_1907,N_2647);
and U3713 (N_3713,N_1943,N_2448);
nor U3714 (N_3714,N_1777,N_2208);
xnor U3715 (N_3715,N_2393,N_2527);
nor U3716 (N_3716,N_2076,N_2770);
nor U3717 (N_3717,N_1680,N_2232);
and U3718 (N_3718,N_1702,N_2079);
or U3719 (N_3719,N_2335,N_2910);
xor U3720 (N_3720,N_2149,N_2542);
nor U3721 (N_3721,N_1679,N_2548);
xor U3722 (N_3722,N_2286,N_2651);
nor U3723 (N_3723,N_1637,N_2474);
and U3724 (N_3724,N_1935,N_2883);
nand U3725 (N_3725,N_2235,N_1515);
nor U3726 (N_3726,N_2769,N_1676);
xnor U3727 (N_3727,N_2047,N_1850);
and U3728 (N_3728,N_2725,N_2163);
nor U3729 (N_3729,N_1897,N_2280);
and U3730 (N_3730,N_1704,N_1880);
nand U3731 (N_3731,N_1926,N_2059);
xnor U3732 (N_3732,N_1599,N_1748);
nor U3733 (N_3733,N_1831,N_2194);
nor U3734 (N_3734,N_2202,N_2418);
or U3735 (N_3735,N_1936,N_2410);
xor U3736 (N_3736,N_2584,N_2305);
xnor U3737 (N_3737,N_1980,N_1741);
or U3738 (N_3738,N_1802,N_2976);
and U3739 (N_3739,N_1859,N_2634);
and U3740 (N_3740,N_1542,N_1558);
and U3741 (N_3741,N_2985,N_2120);
nand U3742 (N_3742,N_1644,N_2028);
nand U3743 (N_3743,N_1794,N_1853);
and U3744 (N_3744,N_1895,N_2480);
nand U3745 (N_3745,N_1894,N_2687);
or U3746 (N_3746,N_2087,N_1606);
and U3747 (N_3747,N_2433,N_2485);
and U3748 (N_3748,N_1994,N_2846);
or U3749 (N_3749,N_1864,N_1807);
and U3750 (N_3750,N_1629,N_2269);
nand U3751 (N_3751,N_2008,N_2217);
and U3752 (N_3752,N_2757,N_1922);
or U3753 (N_3753,N_2399,N_1895);
or U3754 (N_3754,N_2656,N_2813);
and U3755 (N_3755,N_1808,N_1882);
nor U3756 (N_3756,N_1804,N_1561);
and U3757 (N_3757,N_1756,N_2123);
and U3758 (N_3758,N_2063,N_1692);
and U3759 (N_3759,N_2032,N_2346);
and U3760 (N_3760,N_2983,N_1716);
and U3761 (N_3761,N_2978,N_2756);
xnor U3762 (N_3762,N_1532,N_1716);
nand U3763 (N_3763,N_2773,N_2902);
nor U3764 (N_3764,N_2917,N_2003);
xnor U3765 (N_3765,N_1877,N_1522);
or U3766 (N_3766,N_2325,N_2863);
nand U3767 (N_3767,N_2854,N_1665);
nand U3768 (N_3768,N_2157,N_2798);
nand U3769 (N_3769,N_1783,N_2157);
xnor U3770 (N_3770,N_2144,N_1720);
xnor U3771 (N_3771,N_2210,N_2097);
and U3772 (N_3772,N_1622,N_2786);
and U3773 (N_3773,N_2158,N_1879);
and U3774 (N_3774,N_2453,N_2333);
xor U3775 (N_3775,N_2083,N_1522);
nand U3776 (N_3776,N_2693,N_2977);
xor U3777 (N_3777,N_2044,N_2804);
nand U3778 (N_3778,N_1981,N_2330);
xnor U3779 (N_3779,N_1709,N_2336);
nor U3780 (N_3780,N_1776,N_2257);
nand U3781 (N_3781,N_1581,N_1790);
nand U3782 (N_3782,N_2268,N_2770);
nor U3783 (N_3783,N_1787,N_2863);
nand U3784 (N_3784,N_1610,N_2040);
nor U3785 (N_3785,N_1679,N_2739);
and U3786 (N_3786,N_2143,N_1613);
nor U3787 (N_3787,N_2045,N_2317);
and U3788 (N_3788,N_2171,N_1552);
or U3789 (N_3789,N_1557,N_2716);
nor U3790 (N_3790,N_2686,N_2936);
nor U3791 (N_3791,N_2322,N_1537);
nor U3792 (N_3792,N_2806,N_1528);
nor U3793 (N_3793,N_1875,N_2199);
or U3794 (N_3794,N_2324,N_2112);
nor U3795 (N_3795,N_2370,N_2675);
or U3796 (N_3796,N_2893,N_2037);
nand U3797 (N_3797,N_2128,N_2411);
xor U3798 (N_3798,N_2119,N_2627);
or U3799 (N_3799,N_1801,N_1523);
xor U3800 (N_3800,N_1746,N_1948);
or U3801 (N_3801,N_2943,N_1596);
nand U3802 (N_3802,N_1533,N_2278);
or U3803 (N_3803,N_1567,N_2668);
nand U3804 (N_3804,N_1892,N_1966);
nor U3805 (N_3805,N_2621,N_2188);
nand U3806 (N_3806,N_2700,N_2296);
and U3807 (N_3807,N_2139,N_2644);
nor U3808 (N_3808,N_2498,N_2891);
or U3809 (N_3809,N_1718,N_1505);
xnor U3810 (N_3810,N_2608,N_2732);
and U3811 (N_3811,N_2935,N_2109);
nand U3812 (N_3812,N_1908,N_2586);
nor U3813 (N_3813,N_2822,N_2769);
or U3814 (N_3814,N_1852,N_1871);
nand U3815 (N_3815,N_2327,N_2061);
nor U3816 (N_3816,N_1929,N_2952);
nor U3817 (N_3817,N_1602,N_2353);
nor U3818 (N_3818,N_2934,N_2057);
and U3819 (N_3819,N_2611,N_1588);
or U3820 (N_3820,N_1687,N_2526);
and U3821 (N_3821,N_1667,N_1990);
or U3822 (N_3822,N_2056,N_2576);
and U3823 (N_3823,N_2655,N_2278);
and U3824 (N_3824,N_2903,N_2677);
nor U3825 (N_3825,N_2647,N_1671);
or U3826 (N_3826,N_2514,N_2721);
or U3827 (N_3827,N_2769,N_2048);
and U3828 (N_3828,N_2768,N_2919);
xor U3829 (N_3829,N_1852,N_2484);
and U3830 (N_3830,N_2137,N_2988);
or U3831 (N_3831,N_1862,N_1939);
and U3832 (N_3832,N_2555,N_2657);
or U3833 (N_3833,N_2014,N_2935);
or U3834 (N_3834,N_2325,N_2170);
nor U3835 (N_3835,N_1672,N_2936);
nand U3836 (N_3836,N_1750,N_2107);
nor U3837 (N_3837,N_2240,N_2902);
nand U3838 (N_3838,N_1510,N_1857);
nor U3839 (N_3839,N_2227,N_2488);
nor U3840 (N_3840,N_2623,N_1533);
nand U3841 (N_3841,N_2328,N_2284);
or U3842 (N_3842,N_1577,N_2606);
nand U3843 (N_3843,N_1771,N_1927);
nor U3844 (N_3844,N_2704,N_2724);
nor U3845 (N_3845,N_1910,N_1638);
nor U3846 (N_3846,N_2794,N_2782);
or U3847 (N_3847,N_1690,N_2567);
or U3848 (N_3848,N_2488,N_1978);
or U3849 (N_3849,N_2173,N_1794);
or U3850 (N_3850,N_2992,N_2498);
nand U3851 (N_3851,N_1675,N_2158);
nor U3852 (N_3852,N_1900,N_1573);
or U3853 (N_3853,N_1903,N_2159);
or U3854 (N_3854,N_1617,N_1515);
xnor U3855 (N_3855,N_1796,N_1704);
or U3856 (N_3856,N_1801,N_1857);
nor U3857 (N_3857,N_2561,N_2054);
nand U3858 (N_3858,N_2081,N_2575);
and U3859 (N_3859,N_2797,N_1653);
or U3860 (N_3860,N_2000,N_1842);
nand U3861 (N_3861,N_2708,N_2649);
xnor U3862 (N_3862,N_2114,N_2556);
nor U3863 (N_3863,N_2871,N_2067);
nand U3864 (N_3864,N_2230,N_2641);
nand U3865 (N_3865,N_1903,N_2891);
nand U3866 (N_3866,N_1760,N_1886);
or U3867 (N_3867,N_1663,N_1646);
and U3868 (N_3868,N_2814,N_2883);
and U3869 (N_3869,N_1874,N_1606);
nand U3870 (N_3870,N_1654,N_1875);
or U3871 (N_3871,N_2718,N_1916);
nand U3872 (N_3872,N_2193,N_2726);
or U3873 (N_3873,N_2505,N_2009);
or U3874 (N_3874,N_1688,N_1989);
and U3875 (N_3875,N_1609,N_1551);
nor U3876 (N_3876,N_2464,N_2064);
xnor U3877 (N_3877,N_2662,N_2303);
xnor U3878 (N_3878,N_2176,N_1591);
and U3879 (N_3879,N_2838,N_1797);
nand U3880 (N_3880,N_2002,N_2419);
nand U3881 (N_3881,N_2990,N_1531);
and U3882 (N_3882,N_2207,N_2676);
xnor U3883 (N_3883,N_1643,N_2664);
nand U3884 (N_3884,N_1829,N_1635);
nand U3885 (N_3885,N_2209,N_2212);
nand U3886 (N_3886,N_2139,N_1594);
nor U3887 (N_3887,N_1982,N_2527);
nand U3888 (N_3888,N_2451,N_2305);
xor U3889 (N_3889,N_1888,N_1789);
nor U3890 (N_3890,N_1734,N_1542);
nand U3891 (N_3891,N_2462,N_2477);
nand U3892 (N_3892,N_1639,N_2319);
nand U3893 (N_3893,N_2381,N_2630);
nor U3894 (N_3894,N_2218,N_2791);
nand U3895 (N_3895,N_2240,N_2386);
nor U3896 (N_3896,N_2265,N_1541);
nand U3897 (N_3897,N_2772,N_2802);
nor U3898 (N_3898,N_1982,N_2633);
and U3899 (N_3899,N_2789,N_2337);
and U3900 (N_3900,N_1781,N_1991);
nand U3901 (N_3901,N_2664,N_1830);
xor U3902 (N_3902,N_2500,N_2405);
or U3903 (N_3903,N_1507,N_1630);
nor U3904 (N_3904,N_2070,N_1989);
and U3905 (N_3905,N_2694,N_1554);
xor U3906 (N_3906,N_2842,N_2612);
nor U3907 (N_3907,N_2014,N_2532);
or U3908 (N_3908,N_1672,N_1834);
and U3909 (N_3909,N_1937,N_1518);
or U3910 (N_3910,N_2960,N_2179);
nor U3911 (N_3911,N_1959,N_1685);
nand U3912 (N_3912,N_2382,N_1735);
nand U3913 (N_3913,N_1602,N_2080);
nand U3914 (N_3914,N_2642,N_2392);
or U3915 (N_3915,N_2255,N_2587);
or U3916 (N_3916,N_2344,N_1951);
nor U3917 (N_3917,N_2721,N_2851);
and U3918 (N_3918,N_1804,N_2683);
nand U3919 (N_3919,N_2294,N_2371);
xor U3920 (N_3920,N_2400,N_2129);
or U3921 (N_3921,N_1502,N_2201);
and U3922 (N_3922,N_2087,N_1963);
or U3923 (N_3923,N_1601,N_1505);
nor U3924 (N_3924,N_2703,N_2807);
and U3925 (N_3925,N_1833,N_2201);
and U3926 (N_3926,N_2268,N_2358);
and U3927 (N_3927,N_2579,N_2927);
nand U3928 (N_3928,N_1512,N_2520);
and U3929 (N_3929,N_1559,N_2440);
nand U3930 (N_3930,N_2931,N_2340);
and U3931 (N_3931,N_2337,N_2285);
nand U3932 (N_3932,N_2626,N_2226);
or U3933 (N_3933,N_2974,N_2833);
and U3934 (N_3934,N_2970,N_2257);
nand U3935 (N_3935,N_1547,N_2785);
or U3936 (N_3936,N_2944,N_2811);
or U3937 (N_3937,N_2285,N_2714);
nand U3938 (N_3938,N_2867,N_2224);
or U3939 (N_3939,N_2870,N_1890);
and U3940 (N_3940,N_2860,N_1641);
or U3941 (N_3941,N_1742,N_2988);
nor U3942 (N_3942,N_1941,N_2261);
nand U3943 (N_3943,N_1997,N_2492);
or U3944 (N_3944,N_1792,N_2718);
or U3945 (N_3945,N_1810,N_2989);
nand U3946 (N_3946,N_2568,N_2188);
nand U3947 (N_3947,N_2252,N_2332);
or U3948 (N_3948,N_2988,N_2610);
or U3949 (N_3949,N_2622,N_1974);
nand U3950 (N_3950,N_2975,N_2330);
nor U3951 (N_3951,N_1619,N_2078);
or U3952 (N_3952,N_1682,N_2088);
xnor U3953 (N_3953,N_2178,N_2093);
xnor U3954 (N_3954,N_1914,N_2428);
or U3955 (N_3955,N_2064,N_2763);
and U3956 (N_3956,N_2266,N_2691);
nand U3957 (N_3957,N_2032,N_2051);
xnor U3958 (N_3958,N_1635,N_1919);
xnor U3959 (N_3959,N_2184,N_2955);
nand U3960 (N_3960,N_2733,N_2577);
nor U3961 (N_3961,N_2811,N_1690);
and U3962 (N_3962,N_2637,N_1867);
nor U3963 (N_3963,N_2516,N_2274);
or U3964 (N_3964,N_2899,N_2446);
and U3965 (N_3965,N_2038,N_1986);
nor U3966 (N_3966,N_1896,N_2023);
and U3967 (N_3967,N_2266,N_2037);
or U3968 (N_3968,N_2244,N_2328);
and U3969 (N_3969,N_2173,N_2301);
nand U3970 (N_3970,N_2367,N_1800);
or U3971 (N_3971,N_1998,N_2639);
or U3972 (N_3972,N_2815,N_2842);
nand U3973 (N_3973,N_1843,N_2550);
and U3974 (N_3974,N_1707,N_1569);
nor U3975 (N_3975,N_1987,N_2522);
nor U3976 (N_3976,N_1742,N_2206);
nor U3977 (N_3977,N_2883,N_1916);
and U3978 (N_3978,N_1600,N_2559);
and U3979 (N_3979,N_2826,N_2000);
or U3980 (N_3980,N_1917,N_1527);
or U3981 (N_3981,N_2891,N_2390);
nand U3982 (N_3982,N_2178,N_1550);
nor U3983 (N_3983,N_1912,N_1553);
and U3984 (N_3984,N_2122,N_2099);
nor U3985 (N_3985,N_1965,N_1560);
xor U3986 (N_3986,N_2819,N_2647);
nand U3987 (N_3987,N_2908,N_1996);
nand U3988 (N_3988,N_2037,N_1631);
nor U3989 (N_3989,N_2035,N_1968);
and U3990 (N_3990,N_2913,N_1831);
nand U3991 (N_3991,N_1655,N_2555);
nor U3992 (N_3992,N_2019,N_2078);
or U3993 (N_3993,N_2641,N_2214);
and U3994 (N_3994,N_1692,N_2337);
nand U3995 (N_3995,N_2917,N_2333);
nor U3996 (N_3996,N_1667,N_2759);
and U3997 (N_3997,N_2264,N_1695);
nor U3998 (N_3998,N_2274,N_2515);
or U3999 (N_3999,N_1621,N_2975);
and U4000 (N_4000,N_2908,N_2644);
or U4001 (N_4001,N_1796,N_1758);
nand U4002 (N_4002,N_1964,N_1838);
or U4003 (N_4003,N_2132,N_1823);
xnor U4004 (N_4004,N_1888,N_2697);
nand U4005 (N_4005,N_2304,N_2901);
nor U4006 (N_4006,N_1503,N_2313);
nor U4007 (N_4007,N_2081,N_1588);
nor U4008 (N_4008,N_2330,N_2214);
and U4009 (N_4009,N_2888,N_2074);
and U4010 (N_4010,N_1625,N_2578);
nor U4011 (N_4011,N_2397,N_1972);
or U4012 (N_4012,N_1552,N_2094);
or U4013 (N_4013,N_2282,N_1793);
nand U4014 (N_4014,N_2768,N_2004);
nor U4015 (N_4015,N_2300,N_2200);
and U4016 (N_4016,N_1870,N_2919);
and U4017 (N_4017,N_2877,N_1941);
nand U4018 (N_4018,N_1629,N_2560);
nor U4019 (N_4019,N_2675,N_1809);
or U4020 (N_4020,N_2253,N_1823);
and U4021 (N_4021,N_1776,N_2805);
or U4022 (N_4022,N_2165,N_2151);
or U4023 (N_4023,N_2946,N_1840);
xnor U4024 (N_4024,N_2065,N_2419);
and U4025 (N_4025,N_2850,N_2809);
or U4026 (N_4026,N_1904,N_1670);
or U4027 (N_4027,N_2882,N_1545);
nor U4028 (N_4028,N_2476,N_1917);
nor U4029 (N_4029,N_2429,N_2796);
nor U4030 (N_4030,N_2662,N_1833);
and U4031 (N_4031,N_2151,N_2150);
nor U4032 (N_4032,N_2364,N_1527);
and U4033 (N_4033,N_1607,N_1914);
nor U4034 (N_4034,N_2343,N_2966);
nor U4035 (N_4035,N_1516,N_2750);
nor U4036 (N_4036,N_1593,N_2728);
or U4037 (N_4037,N_2058,N_2293);
and U4038 (N_4038,N_2749,N_1779);
or U4039 (N_4039,N_2733,N_2646);
nand U4040 (N_4040,N_2517,N_2670);
or U4041 (N_4041,N_2986,N_1619);
nor U4042 (N_4042,N_2491,N_1591);
nand U4043 (N_4043,N_2134,N_2385);
nand U4044 (N_4044,N_2620,N_2984);
nor U4045 (N_4045,N_2320,N_1756);
and U4046 (N_4046,N_1834,N_2856);
and U4047 (N_4047,N_1840,N_2569);
or U4048 (N_4048,N_1898,N_1659);
and U4049 (N_4049,N_1675,N_1951);
and U4050 (N_4050,N_2674,N_2760);
xnor U4051 (N_4051,N_2246,N_2602);
or U4052 (N_4052,N_2203,N_1882);
nand U4053 (N_4053,N_2527,N_2844);
xnor U4054 (N_4054,N_1928,N_1842);
and U4055 (N_4055,N_1505,N_1697);
nor U4056 (N_4056,N_2169,N_1969);
xor U4057 (N_4057,N_2110,N_2035);
nor U4058 (N_4058,N_1809,N_2613);
nor U4059 (N_4059,N_1601,N_2852);
nor U4060 (N_4060,N_2750,N_2075);
and U4061 (N_4061,N_2417,N_2087);
xor U4062 (N_4062,N_1860,N_1878);
nor U4063 (N_4063,N_2609,N_1519);
and U4064 (N_4064,N_1582,N_1598);
nand U4065 (N_4065,N_1791,N_2710);
and U4066 (N_4066,N_2033,N_1739);
nor U4067 (N_4067,N_1723,N_2971);
and U4068 (N_4068,N_2182,N_2244);
or U4069 (N_4069,N_1947,N_2745);
nor U4070 (N_4070,N_2066,N_2650);
or U4071 (N_4071,N_2926,N_2245);
or U4072 (N_4072,N_2159,N_2591);
xor U4073 (N_4073,N_1918,N_2456);
and U4074 (N_4074,N_2328,N_2236);
and U4075 (N_4075,N_2613,N_2813);
or U4076 (N_4076,N_2447,N_1768);
xor U4077 (N_4077,N_1870,N_2995);
nand U4078 (N_4078,N_2956,N_2393);
and U4079 (N_4079,N_1781,N_2113);
nor U4080 (N_4080,N_2460,N_2467);
nor U4081 (N_4081,N_2698,N_2357);
or U4082 (N_4082,N_1956,N_2342);
nor U4083 (N_4083,N_2271,N_2547);
and U4084 (N_4084,N_1628,N_2418);
or U4085 (N_4085,N_2698,N_1837);
and U4086 (N_4086,N_1903,N_2486);
or U4087 (N_4087,N_2064,N_1617);
nor U4088 (N_4088,N_2493,N_2519);
xnor U4089 (N_4089,N_2697,N_2594);
nor U4090 (N_4090,N_2664,N_2370);
nand U4091 (N_4091,N_1700,N_2748);
nor U4092 (N_4092,N_2144,N_1515);
nand U4093 (N_4093,N_2658,N_2128);
or U4094 (N_4094,N_2442,N_1869);
nor U4095 (N_4095,N_2923,N_2164);
nand U4096 (N_4096,N_2487,N_1785);
or U4097 (N_4097,N_2706,N_2222);
nand U4098 (N_4098,N_2438,N_2862);
and U4099 (N_4099,N_2039,N_2537);
xnor U4100 (N_4100,N_2317,N_1894);
xnor U4101 (N_4101,N_1551,N_2837);
and U4102 (N_4102,N_1759,N_2195);
or U4103 (N_4103,N_1628,N_2656);
and U4104 (N_4104,N_2513,N_1516);
nand U4105 (N_4105,N_2369,N_1673);
nand U4106 (N_4106,N_2893,N_1741);
and U4107 (N_4107,N_1971,N_2837);
nand U4108 (N_4108,N_1597,N_1703);
nand U4109 (N_4109,N_2011,N_1679);
nand U4110 (N_4110,N_2644,N_2839);
nand U4111 (N_4111,N_1979,N_2928);
nor U4112 (N_4112,N_2141,N_1956);
or U4113 (N_4113,N_2151,N_2056);
xnor U4114 (N_4114,N_2120,N_2677);
nor U4115 (N_4115,N_1624,N_2571);
and U4116 (N_4116,N_2394,N_2916);
or U4117 (N_4117,N_2638,N_1609);
nor U4118 (N_4118,N_1506,N_2910);
and U4119 (N_4119,N_2223,N_2200);
nor U4120 (N_4120,N_1862,N_2845);
or U4121 (N_4121,N_2969,N_2210);
nand U4122 (N_4122,N_1854,N_2494);
nand U4123 (N_4123,N_1601,N_1545);
and U4124 (N_4124,N_2991,N_2702);
nand U4125 (N_4125,N_1801,N_2814);
or U4126 (N_4126,N_2475,N_1595);
and U4127 (N_4127,N_1801,N_2317);
xor U4128 (N_4128,N_1567,N_2894);
nand U4129 (N_4129,N_1505,N_2752);
nand U4130 (N_4130,N_1550,N_1535);
nor U4131 (N_4131,N_2869,N_1882);
nor U4132 (N_4132,N_2107,N_1570);
and U4133 (N_4133,N_2456,N_2649);
nand U4134 (N_4134,N_2424,N_2430);
nand U4135 (N_4135,N_2943,N_1962);
nand U4136 (N_4136,N_2589,N_1546);
xor U4137 (N_4137,N_1895,N_2597);
and U4138 (N_4138,N_1806,N_2982);
nor U4139 (N_4139,N_2117,N_2398);
nand U4140 (N_4140,N_2887,N_1832);
nand U4141 (N_4141,N_2298,N_2845);
or U4142 (N_4142,N_1773,N_2843);
or U4143 (N_4143,N_2473,N_2391);
nor U4144 (N_4144,N_2468,N_1510);
nor U4145 (N_4145,N_1984,N_2306);
nand U4146 (N_4146,N_2488,N_1530);
and U4147 (N_4147,N_2606,N_1621);
and U4148 (N_4148,N_1929,N_1615);
xnor U4149 (N_4149,N_2924,N_2870);
and U4150 (N_4150,N_2682,N_2608);
nand U4151 (N_4151,N_1527,N_1928);
nor U4152 (N_4152,N_2727,N_2273);
nor U4153 (N_4153,N_2632,N_2228);
nand U4154 (N_4154,N_1595,N_2987);
and U4155 (N_4155,N_2963,N_2057);
xor U4156 (N_4156,N_1944,N_2563);
xor U4157 (N_4157,N_1935,N_2974);
and U4158 (N_4158,N_1548,N_1596);
nor U4159 (N_4159,N_1882,N_2616);
and U4160 (N_4160,N_1748,N_2076);
nand U4161 (N_4161,N_1940,N_2543);
and U4162 (N_4162,N_2909,N_1761);
nand U4163 (N_4163,N_2528,N_2002);
xnor U4164 (N_4164,N_2954,N_2396);
and U4165 (N_4165,N_2622,N_1762);
or U4166 (N_4166,N_2446,N_1591);
or U4167 (N_4167,N_2291,N_2225);
nor U4168 (N_4168,N_1750,N_2558);
nor U4169 (N_4169,N_2268,N_2861);
nand U4170 (N_4170,N_1807,N_2331);
and U4171 (N_4171,N_2011,N_2480);
and U4172 (N_4172,N_2827,N_2333);
xnor U4173 (N_4173,N_2295,N_2326);
or U4174 (N_4174,N_1653,N_2821);
nand U4175 (N_4175,N_2505,N_2074);
nor U4176 (N_4176,N_2658,N_2788);
or U4177 (N_4177,N_2967,N_2360);
nor U4178 (N_4178,N_1664,N_1713);
nand U4179 (N_4179,N_1920,N_2622);
and U4180 (N_4180,N_2646,N_1631);
nand U4181 (N_4181,N_2191,N_2004);
xor U4182 (N_4182,N_2604,N_2496);
or U4183 (N_4183,N_2679,N_1669);
nand U4184 (N_4184,N_1637,N_2385);
nor U4185 (N_4185,N_1669,N_2353);
nand U4186 (N_4186,N_1588,N_1577);
nor U4187 (N_4187,N_1602,N_2289);
nor U4188 (N_4188,N_1575,N_1625);
nand U4189 (N_4189,N_2093,N_2802);
nor U4190 (N_4190,N_1732,N_2041);
nand U4191 (N_4191,N_1820,N_2206);
and U4192 (N_4192,N_2011,N_2147);
or U4193 (N_4193,N_2441,N_1603);
or U4194 (N_4194,N_2054,N_1605);
nand U4195 (N_4195,N_2137,N_2572);
nand U4196 (N_4196,N_2272,N_1739);
nand U4197 (N_4197,N_2294,N_1695);
or U4198 (N_4198,N_2253,N_2739);
or U4199 (N_4199,N_2002,N_2849);
and U4200 (N_4200,N_2414,N_2238);
nand U4201 (N_4201,N_2889,N_2020);
nor U4202 (N_4202,N_2106,N_2643);
nand U4203 (N_4203,N_2668,N_2759);
xnor U4204 (N_4204,N_2600,N_2415);
nor U4205 (N_4205,N_1663,N_1762);
nor U4206 (N_4206,N_2792,N_2872);
or U4207 (N_4207,N_2291,N_2236);
or U4208 (N_4208,N_2259,N_2357);
nand U4209 (N_4209,N_2943,N_2389);
or U4210 (N_4210,N_2406,N_2399);
nor U4211 (N_4211,N_2031,N_2222);
nand U4212 (N_4212,N_2603,N_2898);
and U4213 (N_4213,N_2672,N_2557);
nand U4214 (N_4214,N_1710,N_2229);
nand U4215 (N_4215,N_2709,N_2149);
nor U4216 (N_4216,N_1535,N_2883);
and U4217 (N_4217,N_2579,N_2107);
and U4218 (N_4218,N_2770,N_2503);
or U4219 (N_4219,N_2199,N_2596);
and U4220 (N_4220,N_2971,N_2471);
and U4221 (N_4221,N_1512,N_1819);
and U4222 (N_4222,N_2374,N_2003);
nor U4223 (N_4223,N_1849,N_1622);
or U4224 (N_4224,N_2716,N_1575);
or U4225 (N_4225,N_1751,N_1659);
nand U4226 (N_4226,N_2132,N_2718);
and U4227 (N_4227,N_2207,N_1697);
nor U4228 (N_4228,N_2388,N_2381);
nor U4229 (N_4229,N_1729,N_2376);
nand U4230 (N_4230,N_2473,N_1851);
xor U4231 (N_4231,N_2473,N_1893);
or U4232 (N_4232,N_2356,N_2921);
or U4233 (N_4233,N_2543,N_2971);
or U4234 (N_4234,N_2271,N_1656);
nand U4235 (N_4235,N_2771,N_2811);
nor U4236 (N_4236,N_1521,N_1634);
and U4237 (N_4237,N_1669,N_2668);
nand U4238 (N_4238,N_1663,N_2848);
nor U4239 (N_4239,N_2255,N_2718);
and U4240 (N_4240,N_2396,N_2874);
or U4241 (N_4241,N_1848,N_1732);
xor U4242 (N_4242,N_2302,N_1895);
nand U4243 (N_4243,N_2732,N_1611);
xor U4244 (N_4244,N_2722,N_1717);
nor U4245 (N_4245,N_2203,N_2798);
xor U4246 (N_4246,N_2334,N_2567);
nor U4247 (N_4247,N_2499,N_2385);
or U4248 (N_4248,N_1712,N_1603);
and U4249 (N_4249,N_2454,N_1889);
or U4250 (N_4250,N_1653,N_1655);
and U4251 (N_4251,N_1883,N_2936);
nor U4252 (N_4252,N_2217,N_2334);
and U4253 (N_4253,N_2269,N_2860);
nor U4254 (N_4254,N_2024,N_2056);
nor U4255 (N_4255,N_1954,N_2303);
nor U4256 (N_4256,N_2320,N_1670);
nor U4257 (N_4257,N_2554,N_2600);
or U4258 (N_4258,N_2724,N_2099);
nand U4259 (N_4259,N_1762,N_2728);
and U4260 (N_4260,N_2756,N_2472);
xnor U4261 (N_4261,N_1570,N_2807);
or U4262 (N_4262,N_1836,N_1657);
or U4263 (N_4263,N_1931,N_2335);
nor U4264 (N_4264,N_2782,N_2019);
nor U4265 (N_4265,N_2118,N_1805);
and U4266 (N_4266,N_1736,N_2823);
and U4267 (N_4267,N_1979,N_1810);
nor U4268 (N_4268,N_1656,N_2874);
nor U4269 (N_4269,N_2640,N_2550);
nand U4270 (N_4270,N_1847,N_2692);
or U4271 (N_4271,N_1609,N_1739);
nor U4272 (N_4272,N_2486,N_2008);
nand U4273 (N_4273,N_2600,N_2740);
nor U4274 (N_4274,N_1931,N_2437);
nor U4275 (N_4275,N_1796,N_2445);
nand U4276 (N_4276,N_1792,N_1622);
or U4277 (N_4277,N_2535,N_2241);
and U4278 (N_4278,N_1536,N_1542);
or U4279 (N_4279,N_2736,N_1607);
nand U4280 (N_4280,N_1530,N_2962);
nor U4281 (N_4281,N_1790,N_2031);
nand U4282 (N_4282,N_1931,N_2715);
nor U4283 (N_4283,N_2024,N_2473);
nor U4284 (N_4284,N_2695,N_1544);
nor U4285 (N_4285,N_2647,N_2013);
nand U4286 (N_4286,N_2489,N_1551);
or U4287 (N_4287,N_2112,N_2299);
or U4288 (N_4288,N_2724,N_2191);
and U4289 (N_4289,N_2305,N_2974);
nand U4290 (N_4290,N_1809,N_2874);
or U4291 (N_4291,N_2609,N_2661);
or U4292 (N_4292,N_2460,N_1978);
or U4293 (N_4293,N_2500,N_2702);
nor U4294 (N_4294,N_2252,N_2360);
or U4295 (N_4295,N_1889,N_2446);
and U4296 (N_4296,N_2381,N_2648);
xnor U4297 (N_4297,N_1951,N_2271);
or U4298 (N_4298,N_2785,N_2254);
and U4299 (N_4299,N_2128,N_2167);
xor U4300 (N_4300,N_2002,N_1998);
nor U4301 (N_4301,N_1813,N_2751);
nor U4302 (N_4302,N_2337,N_2674);
nand U4303 (N_4303,N_1733,N_1537);
or U4304 (N_4304,N_1517,N_1937);
and U4305 (N_4305,N_1913,N_1752);
and U4306 (N_4306,N_2748,N_1958);
nand U4307 (N_4307,N_1771,N_2016);
and U4308 (N_4308,N_2128,N_1560);
nor U4309 (N_4309,N_2204,N_2951);
nor U4310 (N_4310,N_2918,N_1572);
nor U4311 (N_4311,N_2787,N_2846);
nor U4312 (N_4312,N_2001,N_2953);
xor U4313 (N_4313,N_2572,N_2159);
nor U4314 (N_4314,N_2737,N_1520);
xnor U4315 (N_4315,N_1583,N_2142);
nor U4316 (N_4316,N_2513,N_2635);
xor U4317 (N_4317,N_1772,N_1922);
nand U4318 (N_4318,N_2592,N_2048);
nor U4319 (N_4319,N_2013,N_1802);
and U4320 (N_4320,N_1533,N_2656);
nor U4321 (N_4321,N_2704,N_1927);
nand U4322 (N_4322,N_2625,N_2076);
or U4323 (N_4323,N_1666,N_2452);
and U4324 (N_4324,N_1660,N_1883);
xor U4325 (N_4325,N_1590,N_2971);
nand U4326 (N_4326,N_2413,N_2997);
and U4327 (N_4327,N_2835,N_2819);
nor U4328 (N_4328,N_1809,N_1598);
and U4329 (N_4329,N_1925,N_2340);
nand U4330 (N_4330,N_1665,N_1640);
nand U4331 (N_4331,N_2346,N_1648);
and U4332 (N_4332,N_2888,N_2311);
or U4333 (N_4333,N_2760,N_2794);
or U4334 (N_4334,N_1800,N_2332);
or U4335 (N_4335,N_1910,N_1866);
or U4336 (N_4336,N_2924,N_2523);
nand U4337 (N_4337,N_2981,N_2505);
or U4338 (N_4338,N_2120,N_1910);
nand U4339 (N_4339,N_1891,N_1660);
nand U4340 (N_4340,N_1958,N_2979);
or U4341 (N_4341,N_2032,N_2459);
or U4342 (N_4342,N_1981,N_2435);
and U4343 (N_4343,N_1716,N_2933);
nor U4344 (N_4344,N_2337,N_2550);
nor U4345 (N_4345,N_2652,N_1917);
xnor U4346 (N_4346,N_1550,N_2752);
nand U4347 (N_4347,N_1939,N_2096);
or U4348 (N_4348,N_2902,N_1757);
nand U4349 (N_4349,N_2832,N_2062);
nor U4350 (N_4350,N_2314,N_1902);
nand U4351 (N_4351,N_2648,N_2494);
nor U4352 (N_4352,N_1973,N_2406);
and U4353 (N_4353,N_2005,N_2228);
and U4354 (N_4354,N_2496,N_1606);
or U4355 (N_4355,N_2679,N_1559);
nand U4356 (N_4356,N_1899,N_1964);
and U4357 (N_4357,N_2142,N_2984);
nor U4358 (N_4358,N_2278,N_1897);
and U4359 (N_4359,N_2454,N_1749);
and U4360 (N_4360,N_2556,N_2442);
or U4361 (N_4361,N_2100,N_2606);
or U4362 (N_4362,N_2269,N_1953);
nor U4363 (N_4363,N_1724,N_2727);
nand U4364 (N_4364,N_2186,N_1573);
nand U4365 (N_4365,N_2449,N_1561);
and U4366 (N_4366,N_1902,N_2847);
or U4367 (N_4367,N_1527,N_1674);
xnor U4368 (N_4368,N_1560,N_2153);
nor U4369 (N_4369,N_2990,N_2624);
nand U4370 (N_4370,N_1523,N_2848);
nor U4371 (N_4371,N_2396,N_2344);
and U4372 (N_4372,N_2382,N_2311);
nand U4373 (N_4373,N_2794,N_1674);
xor U4374 (N_4374,N_2066,N_2033);
and U4375 (N_4375,N_2149,N_2108);
nand U4376 (N_4376,N_2655,N_1679);
or U4377 (N_4377,N_2343,N_2336);
nor U4378 (N_4378,N_1704,N_2488);
nor U4379 (N_4379,N_2785,N_1937);
xor U4380 (N_4380,N_2053,N_1544);
or U4381 (N_4381,N_2438,N_2206);
or U4382 (N_4382,N_2644,N_1879);
nand U4383 (N_4383,N_2568,N_1809);
or U4384 (N_4384,N_2673,N_1870);
nor U4385 (N_4385,N_2142,N_2508);
nand U4386 (N_4386,N_1722,N_2192);
and U4387 (N_4387,N_1654,N_2211);
nor U4388 (N_4388,N_2064,N_2376);
or U4389 (N_4389,N_1721,N_2847);
nor U4390 (N_4390,N_2884,N_2655);
or U4391 (N_4391,N_2626,N_2544);
xnor U4392 (N_4392,N_1698,N_2238);
xor U4393 (N_4393,N_2681,N_2601);
or U4394 (N_4394,N_1634,N_1968);
and U4395 (N_4395,N_1803,N_1926);
and U4396 (N_4396,N_2864,N_2552);
or U4397 (N_4397,N_1820,N_1821);
and U4398 (N_4398,N_2581,N_2252);
and U4399 (N_4399,N_1740,N_1853);
nand U4400 (N_4400,N_2266,N_2516);
or U4401 (N_4401,N_2768,N_2457);
nand U4402 (N_4402,N_1802,N_2063);
nor U4403 (N_4403,N_1700,N_1958);
xnor U4404 (N_4404,N_2077,N_2053);
or U4405 (N_4405,N_2820,N_1695);
nor U4406 (N_4406,N_2685,N_2690);
xor U4407 (N_4407,N_2249,N_1604);
nand U4408 (N_4408,N_2881,N_2047);
nand U4409 (N_4409,N_1743,N_2956);
nand U4410 (N_4410,N_2250,N_2504);
xnor U4411 (N_4411,N_1562,N_2282);
and U4412 (N_4412,N_1950,N_1584);
and U4413 (N_4413,N_2368,N_1616);
nor U4414 (N_4414,N_2238,N_1860);
and U4415 (N_4415,N_2672,N_2169);
and U4416 (N_4416,N_2595,N_1695);
and U4417 (N_4417,N_2048,N_1677);
nor U4418 (N_4418,N_1718,N_2889);
or U4419 (N_4419,N_2519,N_1635);
nor U4420 (N_4420,N_2787,N_2005);
nand U4421 (N_4421,N_1842,N_2315);
or U4422 (N_4422,N_1502,N_2882);
nor U4423 (N_4423,N_1869,N_1662);
or U4424 (N_4424,N_1546,N_2107);
xor U4425 (N_4425,N_2001,N_1854);
nand U4426 (N_4426,N_2918,N_2922);
and U4427 (N_4427,N_2292,N_2897);
nand U4428 (N_4428,N_2213,N_1901);
xor U4429 (N_4429,N_1976,N_1588);
nand U4430 (N_4430,N_1863,N_2967);
or U4431 (N_4431,N_2850,N_2428);
nor U4432 (N_4432,N_2647,N_1543);
or U4433 (N_4433,N_2592,N_2428);
and U4434 (N_4434,N_1784,N_2992);
and U4435 (N_4435,N_1793,N_2637);
nor U4436 (N_4436,N_1506,N_2045);
nor U4437 (N_4437,N_2156,N_2583);
nor U4438 (N_4438,N_1882,N_2221);
nand U4439 (N_4439,N_2036,N_2959);
and U4440 (N_4440,N_1800,N_2940);
nand U4441 (N_4441,N_1653,N_1609);
or U4442 (N_4442,N_2453,N_2290);
nor U4443 (N_4443,N_2091,N_1603);
nor U4444 (N_4444,N_2050,N_2452);
nor U4445 (N_4445,N_2418,N_1654);
and U4446 (N_4446,N_1749,N_1649);
nor U4447 (N_4447,N_2101,N_1621);
or U4448 (N_4448,N_2324,N_1660);
or U4449 (N_4449,N_2213,N_2275);
nor U4450 (N_4450,N_2148,N_1965);
and U4451 (N_4451,N_2572,N_2720);
and U4452 (N_4452,N_2819,N_2842);
and U4453 (N_4453,N_1962,N_1747);
nand U4454 (N_4454,N_1668,N_1573);
nor U4455 (N_4455,N_2641,N_2042);
nand U4456 (N_4456,N_2063,N_1596);
xor U4457 (N_4457,N_2082,N_2554);
or U4458 (N_4458,N_2502,N_1605);
nand U4459 (N_4459,N_2739,N_2304);
or U4460 (N_4460,N_2211,N_2302);
and U4461 (N_4461,N_2124,N_2464);
nor U4462 (N_4462,N_2914,N_1724);
and U4463 (N_4463,N_1528,N_2053);
xnor U4464 (N_4464,N_2798,N_2530);
and U4465 (N_4465,N_2156,N_2311);
nand U4466 (N_4466,N_2619,N_1996);
nor U4467 (N_4467,N_2646,N_1589);
nor U4468 (N_4468,N_2043,N_1648);
nor U4469 (N_4469,N_2749,N_1532);
and U4470 (N_4470,N_1960,N_1856);
and U4471 (N_4471,N_2181,N_1627);
and U4472 (N_4472,N_2117,N_2244);
xnor U4473 (N_4473,N_2460,N_2237);
nor U4474 (N_4474,N_1542,N_2356);
or U4475 (N_4475,N_2334,N_2647);
and U4476 (N_4476,N_2596,N_1562);
or U4477 (N_4477,N_1805,N_1919);
or U4478 (N_4478,N_2896,N_2963);
nand U4479 (N_4479,N_1913,N_1813);
nand U4480 (N_4480,N_2118,N_2383);
nand U4481 (N_4481,N_2792,N_1718);
nand U4482 (N_4482,N_2429,N_2244);
and U4483 (N_4483,N_2708,N_2379);
nand U4484 (N_4484,N_1791,N_2071);
xnor U4485 (N_4485,N_2580,N_2967);
xor U4486 (N_4486,N_2035,N_1859);
or U4487 (N_4487,N_1890,N_2487);
and U4488 (N_4488,N_1744,N_2858);
nand U4489 (N_4489,N_2529,N_2531);
nor U4490 (N_4490,N_2799,N_1971);
nor U4491 (N_4491,N_2448,N_1549);
nand U4492 (N_4492,N_2523,N_1746);
and U4493 (N_4493,N_2084,N_1814);
nand U4494 (N_4494,N_1945,N_2202);
nor U4495 (N_4495,N_2039,N_2715);
or U4496 (N_4496,N_1746,N_2036);
or U4497 (N_4497,N_2989,N_1918);
and U4498 (N_4498,N_2119,N_2935);
and U4499 (N_4499,N_2141,N_1728);
nand U4500 (N_4500,N_3093,N_3116);
or U4501 (N_4501,N_3785,N_3700);
and U4502 (N_4502,N_3332,N_3582);
nand U4503 (N_4503,N_3171,N_3425);
xnor U4504 (N_4504,N_3967,N_3643);
nand U4505 (N_4505,N_4414,N_4429);
nor U4506 (N_4506,N_3729,N_4196);
nor U4507 (N_4507,N_3519,N_3597);
nor U4508 (N_4508,N_3496,N_4333);
nand U4509 (N_4509,N_3874,N_3500);
or U4510 (N_4510,N_3288,N_3907);
nand U4511 (N_4511,N_3055,N_4206);
nand U4512 (N_4512,N_3654,N_4395);
or U4513 (N_4513,N_3339,N_3109);
xnor U4514 (N_4514,N_4229,N_3992);
or U4515 (N_4515,N_3948,N_4147);
xnor U4516 (N_4516,N_3150,N_3598);
and U4517 (N_4517,N_3124,N_4065);
or U4518 (N_4518,N_4305,N_3819);
nor U4519 (N_4519,N_3843,N_3179);
and U4520 (N_4520,N_3174,N_3004);
or U4521 (N_4521,N_4366,N_3899);
nor U4522 (N_4522,N_3075,N_3138);
nor U4523 (N_4523,N_3790,N_3195);
nor U4524 (N_4524,N_4084,N_3498);
and U4525 (N_4525,N_3632,N_3471);
and U4526 (N_4526,N_3151,N_4054);
and U4527 (N_4527,N_4111,N_3104);
nor U4528 (N_4528,N_4345,N_4160);
and U4529 (N_4529,N_3927,N_3275);
or U4530 (N_4530,N_3086,N_3634);
xor U4531 (N_4531,N_4478,N_4476);
xor U4532 (N_4532,N_3238,N_3715);
nor U4533 (N_4533,N_3367,N_4280);
nand U4534 (N_4534,N_3551,N_4039);
and U4535 (N_4535,N_3812,N_3581);
or U4536 (N_4536,N_3388,N_4415);
nor U4537 (N_4537,N_3144,N_3474);
nand U4538 (N_4538,N_4364,N_3697);
nor U4539 (N_4539,N_3832,N_3123);
nand U4540 (N_4540,N_3111,N_3949);
xnor U4541 (N_4541,N_4471,N_3739);
or U4542 (N_4542,N_3334,N_3090);
nor U4543 (N_4543,N_4473,N_3724);
nor U4544 (N_4544,N_4190,N_3943);
nand U4545 (N_4545,N_3403,N_3497);
or U4546 (N_4546,N_4324,N_4342);
or U4547 (N_4547,N_4393,N_3526);
and U4548 (N_4548,N_3894,N_3390);
nor U4549 (N_4549,N_3505,N_3869);
or U4550 (N_4550,N_3568,N_3987);
nand U4551 (N_4551,N_4254,N_4266);
or U4552 (N_4552,N_3616,N_3001);
and U4553 (N_4553,N_4468,N_3107);
nand U4554 (N_4554,N_3263,N_4083);
nor U4555 (N_4555,N_3098,N_3272);
and U4556 (N_4556,N_3589,N_3572);
and U4557 (N_4557,N_4030,N_3145);
and U4558 (N_4558,N_4077,N_4303);
or U4559 (N_4559,N_3296,N_4340);
nor U4560 (N_4560,N_4269,N_4316);
or U4561 (N_4561,N_3108,N_4390);
and U4562 (N_4562,N_4011,N_3932);
or U4563 (N_4563,N_4347,N_4377);
or U4564 (N_4564,N_3995,N_3845);
nand U4565 (N_4565,N_4056,N_3695);
and U4566 (N_4566,N_4201,N_4355);
and U4567 (N_4567,N_4026,N_4145);
or U4568 (N_4568,N_3494,N_3882);
or U4569 (N_4569,N_3514,N_3596);
nor U4570 (N_4570,N_4219,N_3336);
xor U4571 (N_4571,N_3838,N_4464);
nor U4572 (N_4572,N_3374,N_4365);
nand U4573 (N_4573,N_4226,N_3089);
nor U4574 (N_4574,N_4223,N_4282);
nor U4575 (N_4575,N_3127,N_4463);
and U4576 (N_4576,N_3590,N_3599);
nand U4577 (N_4577,N_3661,N_3017);
nor U4578 (N_4578,N_3342,N_3051);
and U4579 (N_4579,N_3506,N_3659);
nor U4580 (N_4580,N_3372,N_3189);
xor U4581 (N_4581,N_4491,N_3214);
or U4582 (N_4582,N_3522,N_3457);
nor U4583 (N_4583,N_3564,N_4210);
or U4584 (N_4584,N_3278,N_3330);
nand U4585 (N_4585,N_3593,N_3397);
or U4586 (N_4586,N_3938,N_4126);
nand U4587 (N_4587,N_3997,N_4410);
nor U4588 (N_4588,N_3893,N_3934);
nand U4589 (N_4589,N_4300,N_3553);
or U4590 (N_4590,N_4446,N_3312);
nor U4591 (N_4591,N_3813,N_3772);
nor U4592 (N_4592,N_4096,N_4370);
nor U4593 (N_4593,N_3381,N_4297);
or U4594 (N_4594,N_4154,N_3606);
or U4595 (N_4595,N_4214,N_3981);
nor U4596 (N_4596,N_3033,N_4171);
nand U4597 (N_4597,N_4045,N_3576);
nor U4598 (N_4598,N_4010,N_3942);
nor U4599 (N_4599,N_3623,N_3243);
nand U4600 (N_4600,N_4179,N_3972);
or U4601 (N_4601,N_4136,N_3018);
or U4602 (N_4602,N_3102,N_3473);
and U4603 (N_4603,N_3613,N_3309);
or U4604 (N_4604,N_4057,N_4492);
and U4605 (N_4605,N_3765,N_4128);
nand U4606 (N_4606,N_3706,N_4462);
nor U4607 (N_4607,N_3253,N_3904);
nand U4608 (N_4608,N_3610,N_4293);
nand U4609 (N_4609,N_3010,N_4406);
and U4610 (N_4610,N_3698,N_4443);
or U4611 (N_4611,N_3088,N_3207);
nor U4612 (N_4612,N_3852,N_3082);
nand U4613 (N_4613,N_3242,N_4287);
nor U4614 (N_4614,N_3511,N_3476);
nor U4615 (N_4615,N_3683,N_3415);
nand U4616 (N_4616,N_3656,N_4498);
xnor U4617 (N_4617,N_4389,N_3657);
and U4618 (N_4618,N_4115,N_3463);
nand U4619 (N_4619,N_4381,N_4360);
nand U4620 (N_4620,N_3280,N_4367);
nor U4621 (N_4621,N_3912,N_3244);
nand U4622 (N_4622,N_3410,N_4352);
nand U4623 (N_4623,N_4312,N_4213);
nor U4624 (N_4624,N_3628,N_4296);
and U4625 (N_4625,N_3059,N_3226);
xnor U4626 (N_4626,N_4198,N_4022);
and U4627 (N_4627,N_3538,N_4426);
nor U4628 (N_4628,N_3169,N_3071);
and U4629 (N_4629,N_3053,N_3675);
nand U4630 (N_4630,N_3031,N_3173);
or U4631 (N_4631,N_3327,N_3957);
and U4632 (N_4632,N_3513,N_3585);
nor U4633 (N_4633,N_3985,N_3200);
and U4634 (N_4634,N_3629,N_4194);
nor U4635 (N_4635,N_3114,N_3348);
and U4636 (N_4636,N_3741,N_3548);
and U4637 (N_4637,N_3614,N_3639);
nand U4638 (N_4638,N_4442,N_3084);
nor U4639 (N_4639,N_4221,N_3959);
nor U4640 (N_4640,N_3255,N_3557);
or U4641 (N_4641,N_3117,N_3544);
nand U4642 (N_4642,N_3465,N_4187);
or U4643 (N_4643,N_3917,N_4209);
and U4644 (N_4644,N_3023,N_3998);
xor U4645 (N_4645,N_4373,N_4167);
or U4646 (N_4646,N_4341,N_3205);
nand U4647 (N_4647,N_3350,N_4175);
nand U4648 (N_4648,N_4016,N_3445);
and U4649 (N_4649,N_3591,N_3773);
nor U4650 (N_4650,N_3830,N_3196);
nand U4651 (N_4651,N_3693,N_4285);
or U4652 (N_4652,N_3802,N_4088);
xor U4653 (N_4653,N_3543,N_4052);
xnor U4654 (N_4654,N_3925,N_4231);
or U4655 (N_4655,N_3443,N_3218);
and U4656 (N_4656,N_3615,N_4158);
or U4657 (N_4657,N_4397,N_4163);
nand U4658 (N_4658,N_3185,N_3187);
and U4659 (N_4659,N_3328,N_4174);
or U4660 (N_4660,N_3920,N_3627);
nor U4661 (N_4661,N_3274,N_3964);
xnor U4662 (N_4662,N_4104,N_3021);
nor U4663 (N_4663,N_4465,N_3501);
xnor U4664 (N_4664,N_3862,N_3745);
or U4665 (N_4665,N_4081,N_3022);
nand U4666 (N_4666,N_3008,N_4202);
or U4667 (N_4667,N_3820,N_3670);
nor U4668 (N_4668,N_4161,N_3190);
nand U4669 (N_4669,N_4384,N_3736);
and U4670 (N_4670,N_3481,N_4396);
or U4671 (N_4671,N_4286,N_4024);
nor U4672 (N_4672,N_3110,N_3143);
nand U4673 (N_4673,N_3958,N_4078);
nand U4674 (N_4674,N_3137,N_3245);
xor U4675 (N_4675,N_3295,N_3421);
and U4676 (N_4676,N_3678,N_3879);
xnor U4677 (N_4677,N_3666,N_3326);
and U4678 (N_4678,N_4146,N_3735);
and U4679 (N_4679,N_3261,N_4494);
nand U4680 (N_4680,N_3527,N_3704);
and U4681 (N_4681,N_3121,N_4278);
or U4682 (N_4682,N_4449,N_3000);
nor U4683 (N_4683,N_3963,N_3277);
nor U4684 (N_4684,N_3215,N_3989);
nor U4685 (N_4685,N_3645,N_3224);
nor U4686 (N_4686,N_3939,N_3674);
nor U4687 (N_4687,N_3167,N_3779);
nand U4688 (N_4688,N_3106,N_4268);
or U4689 (N_4689,N_4034,N_3573);
nor U4690 (N_4690,N_3699,N_4466);
xor U4691 (N_4691,N_4257,N_3076);
or U4692 (N_4692,N_4317,N_4362);
xnor U4693 (N_4693,N_3132,N_3923);
nand U4694 (N_4694,N_4434,N_4127);
nor U4695 (N_4695,N_3508,N_3234);
nor U4696 (N_4696,N_3152,N_3298);
or U4697 (N_4697,N_4431,N_3030);
nor U4698 (N_4698,N_4421,N_4073);
or U4699 (N_4699,N_4108,N_3754);
xnor U4700 (N_4700,N_3755,N_3032);
xor U4701 (N_4701,N_4181,N_3847);
nor U4702 (N_4702,N_3391,N_3883);
nor U4703 (N_4703,N_4467,N_3436);
nor U4704 (N_4704,N_4448,N_3947);
nor U4705 (N_4705,N_3870,N_4404);
or U4706 (N_4706,N_3133,N_4114);
xnor U4707 (N_4707,N_3447,N_3404);
and U4708 (N_4708,N_4186,N_3836);
or U4709 (N_4709,N_4119,N_3753);
or U4710 (N_4710,N_4197,N_4180);
nor U4711 (N_4711,N_3687,N_3448);
or U4712 (N_4712,N_3530,N_3878);
xor U4713 (N_4713,N_4375,N_4170);
nor U4714 (N_4714,N_3180,N_3141);
nand U4715 (N_4715,N_3746,N_4403);
or U4716 (N_4716,N_4118,N_3147);
or U4717 (N_4717,N_3118,N_4452);
nor U4718 (N_4718,N_4261,N_3077);
xnor U4719 (N_4719,N_4332,N_3814);
nand U4720 (N_4720,N_3913,N_3079);
and U4721 (N_4721,N_3279,N_3542);
nor U4722 (N_4722,N_3554,N_3766);
xor U4723 (N_4723,N_3545,N_3915);
or U4724 (N_4724,N_3744,N_3129);
and U4725 (N_4725,N_4318,N_3094);
nor U4726 (N_4726,N_3284,N_3731);
or U4727 (N_4727,N_3521,N_3398);
nand U4728 (N_4728,N_4242,N_3499);
and U4729 (N_4729,N_3160,N_3536);
xnor U4730 (N_4730,N_4246,N_3502);
and U4731 (N_4731,N_3982,N_3281);
nand U4732 (N_4732,N_3241,N_3461);
or U4733 (N_4733,N_4288,N_4418);
xnor U4734 (N_4734,N_4123,N_3426);
or U4735 (N_4735,N_4255,N_3567);
xnor U4736 (N_4736,N_3440,N_3767);
nor U4737 (N_4737,N_3588,N_4372);
nor U4738 (N_4738,N_3895,N_3113);
xnor U4739 (N_4739,N_3604,N_4249);
or U4740 (N_4740,N_4241,N_4049);
nor U4741 (N_4741,N_3607,N_3125);
xnor U4742 (N_4742,N_3362,N_3120);
and U4743 (N_4743,N_3911,N_4361);
or U4744 (N_4744,N_3087,N_3345);
nor U4745 (N_4745,N_3854,N_3918);
nand U4746 (N_4746,N_3297,N_3069);
nor U4747 (N_4747,N_4250,N_3702);
and U4748 (N_4748,N_3660,N_3701);
nor U4749 (N_4749,N_3406,N_3999);
nand U4750 (N_4750,N_4315,N_4263);
and U4751 (N_4751,N_3592,N_4330);
or U4752 (N_4752,N_4445,N_3317);
or U4753 (N_4753,N_3346,N_4217);
nor U4754 (N_4754,N_4131,N_3617);
xor U4755 (N_4755,N_3561,N_4349);
and U4756 (N_4756,N_3413,N_3338);
xor U4757 (N_4757,N_3763,N_3454);
and U4758 (N_4758,N_3827,N_3050);
or U4759 (N_4759,N_3877,N_3399);
and U4760 (N_4760,N_3323,N_3863);
nor U4761 (N_4761,N_3163,N_3475);
nand U4762 (N_4762,N_3953,N_4433);
nand U4763 (N_4763,N_3844,N_3266);
and U4764 (N_4764,N_4041,N_4321);
nor U4765 (N_4765,N_3751,N_4178);
nand U4766 (N_4766,N_3029,N_3438);
or U4767 (N_4767,N_3624,N_3482);
and U4768 (N_4768,N_3546,N_4405);
nand U4769 (N_4769,N_3377,N_3914);
or U4770 (N_4770,N_4172,N_4038);
nor U4771 (N_4771,N_3733,N_4006);
and U4772 (N_4772,N_4251,N_3770);
xnor U4773 (N_4773,N_3096,N_3209);
or U4774 (N_4774,N_3091,N_4374);
and U4775 (N_4775,N_4139,N_3192);
nand U4776 (N_4776,N_4107,N_4234);
and U4777 (N_4777,N_3804,N_3193);
or U4778 (N_4778,N_3432,N_3191);
nor U4779 (N_4779,N_3864,N_4336);
or U4780 (N_4780,N_3710,N_3930);
and U4781 (N_4781,N_3831,N_3853);
and U4782 (N_4782,N_4053,N_3054);
xor U4783 (N_4783,N_4247,N_3709);
nand U4784 (N_4784,N_3638,N_3100);
xnor U4785 (N_4785,N_3525,N_3928);
nand U4786 (N_4786,N_3198,N_4301);
nand U4787 (N_4787,N_4400,N_4295);
and U4788 (N_4788,N_3762,N_3991);
nand U4789 (N_4789,N_3304,N_4351);
nor U4790 (N_4790,N_3716,N_3756);
or U4791 (N_4791,N_3043,N_3618);
nor U4792 (N_4792,N_4149,N_4066);
and U4793 (N_4793,N_3041,N_3752);
and U4794 (N_4794,N_3287,N_3778);
and U4795 (N_4795,N_3584,N_3386);
or U4796 (N_4796,N_3034,N_4029);
or U4797 (N_4797,N_3897,N_3306);
nand U4798 (N_4798,N_3016,N_3028);
or U4799 (N_4799,N_3423,N_3483);
nand U4800 (N_4800,N_3574,N_3219);
nor U4801 (N_4801,N_3265,N_4132);
and U4802 (N_4802,N_3605,N_4398);
and U4803 (N_4803,N_4094,N_3449);
and U4804 (N_4804,N_3726,N_3974);
and U4805 (N_4805,N_3083,N_3202);
nand U4806 (N_4806,N_3961,N_3504);
and U4807 (N_4807,N_4307,N_3301);
or U4808 (N_4808,N_4207,N_3040);
or U4809 (N_4809,N_4152,N_3650);
and U4810 (N_4810,N_3905,N_4328);
nand U4811 (N_4811,N_3718,N_3216);
nor U4812 (N_4812,N_3990,N_3728);
nand U4813 (N_4813,N_3154,N_3555);
and U4814 (N_4814,N_3886,N_3453);
and U4815 (N_4815,N_4289,N_3042);
nand U4816 (N_4816,N_3227,N_4325);
nor U4817 (N_4817,N_3896,N_3705);
nand U4818 (N_4818,N_3774,N_3612);
nor U4819 (N_4819,N_4382,N_4379);
xor U4820 (N_4820,N_4211,N_4256);
and U4821 (N_4821,N_4051,N_4124);
and U4822 (N_4822,N_3823,N_3601);
nor U4823 (N_4823,N_4479,N_4121);
nor U4824 (N_4824,N_3258,N_3441);
nor U4825 (N_4825,N_3364,N_3149);
or U4826 (N_4826,N_3026,N_3063);
xor U4827 (N_4827,N_3722,N_4125);
nand U4828 (N_4828,N_3865,N_4183);
nand U4829 (N_4829,N_3669,N_4070);
or U4830 (N_4830,N_4290,N_4122);
nor U4831 (N_4831,N_3349,N_3247);
nor U4832 (N_4832,N_4116,N_3800);
nor U4833 (N_4833,N_3455,N_3460);
nand U4834 (N_4834,N_4248,N_4080);
or U4835 (N_4835,N_4168,N_3651);
nand U4836 (N_4836,N_4490,N_4407);
and U4837 (N_4837,N_3383,N_3652);
or U4838 (N_4838,N_3402,N_3062);
or U4839 (N_4839,N_3013,N_3556);
or U4840 (N_4840,N_4032,N_4164);
or U4841 (N_4841,N_4424,N_3369);
and U4842 (N_4842,N_3065,N_4311);
nand U4843 (N_4843,N_4093,N_3045);
nand U4844 (N_4844,N_3437,N_3648);
and U4845 (N_4845,N_4237,N_3305);
and U4846 (N_4846,N_3231,N_4177);
and U4847 (N_4847,N_4157,N_3368);
nor U4848 (N_4848,N_3595,N_3841);
or U4849 (N_4849,N_3560,N_3620);
xor U4850 (N_4850,N_3840,N_3552);
nor U4851 (N_4851,N_3409,N_4117);
or U4852 (N_4852,N_3811,N_3462);
nor U4853 (N_4853,N_4208,N_3230);
and U4854 (N_4854,N_4259,N_3126);
nor U4855 (N_4855,N_3663,N_3818);
nand U4856 (N_4856,N_3725,N_4060);
nand U4857 (N_4857,N_4143,N_3806);
and U4858 (N_4858,N_4033,N_3952);
and U4859 (N_4859,N_3396,N_3846);
nand U4860 (N_4860,N_3837,N_3153);
nor U4861 (N_4861,N_3988,N_3380);
nand U4862 (N_4862,N_3732,N_3518);
nor U4863 (N_4863,N_4275,N_3428);
or U4864 (N_4864,N_3781,N_3512);
nor U4865 (N_4865,N_3792,N_3569);
nor U4866 (N_4866,N_3470,N_3220);
nand U4867 (N_4867,N_4140,N_3039);
xor U4868 (N_4868,N_3533,N_4031);
and U4869 (N_4869,N_3048,N_4264);
xnor U4870 (N_4870,N_3980,N_4142);
and U4871 (N_4871,N_4189,N_4314);
nor U4872 (N_4872,N_4460,N_3450);
and U4873 (N_4873,N_3464,N_3066);
nand U4874 (N_4874,N_4294,N_3922);
nor U4875 (N_4875,N_3801,N_3810);
xor U4876 (N_4876,N_3749,N_3300);
or U4877 (N_4877,N_3035,N_3662);
and U4878 (N_4878,N_4091,N_3851);
nor U4879 (N_4879,N_4169,N_3135);
nor U4880 (N_4880,N_4383,N_3714);
nor U4881 (N_4881,N_4138,N_4222);
and U4882 (N_4882,N_4000,N_3064);
or U4883 (N_4883,N_3472,N_3492);
and U4884 (N_4884,N_4044,N_4099);
xnor U4885 (N_4885,N_3047,N_3290);
or U4886 (N_4886,N_4376,N_3873);
xor U4887 (N_4887,N_3822,N_3320);
nor U4888 (N_4888,N_3510,N_4192);
nor U4889 (N_4889,N_4193,N_4068);
nand U4890 (N_4890,N_4354,N_4310);
nor U4891 (N_4891,N_3337,N_4470);
nor U4892 (N_4892,N_3758,N_3439);
nand U4893 (N_4893,N_3644,N_4244);
nor U4894 (N_4894,N_3547,N_3155);
or U4895 (N_4895,N_3962,N_3252);
or U4896 (N_4896,N_4469,N_3264);
xor U4897 (N_4897,N_3408,N_4428);
xor U4898 (N_4898,N_3467,N_3528);
or U4899 (N_4899,N_4348,N_3641);
xnor U4900 (N_4900,N_3757,N_3427);
nor U4901 (N_4901,N_4475,N_3789);
or U4902 (N_4902,N_3184,N_3405);
xor U4903 (N_4903,N_4474,N_3690);
or U4904 (N_4904,N_3688,N_3433);
and U4905 (N_4905,N_3478,N_3469);
nand U4906 (N_4906,N_3868,N_3771);
and U4907 (N_4907,N_3203,N_3692);
nor U4908 (N_4908,N_3019,N_3575);
or U4909 (N_4909,N_3608,N_3602);
nor U4910 (N_4910,N_4417,N_4074);
nand U4911 (N_4911,N_3260,N_3122);
nand U4912 (N_4912,N_3049,N_3250);
or U4913 (N_4913,N_3855,N_3480);
and U4914 (N_4914,N_3456,N_3983);
xnor U4915 (N_4915,N_3416,N_3668);
nor U4916 (N_4916,N_3080,N_3908);
nor U4917 (N_4917,N_4188,N_3003);
nand U4918 (N_4918,N_3808,N_3024);
nor U4919 (N_4919,N_3929,N_3694);
or U4920 (N_4920,N_3833,N_3681);
xor U4921 (N_4921,N_3935,N_4028);
nor U4922 (N_4922,N_4299,N_3112);
xnor U4923 (N_4923,N_4085,N_4276);
and U4924 (N_4924,N_3468,N_4228);
nor U4925 (N_4925,N_3074,N_4245);
and U4926 (N_4926,N_4399,N_3293);
or U4927 (N_4927,N_4267,N_3027);
nand U4928 (N_4928,N_3849,N_3036);
nor U4929 (N_4929,N_4363,N_3815);
nor U4930 (N_4930,N_4419,N_4040);
xnor U4931 (N_4931,N_3816,N_3887);
nor U4932 (N_4932,N_3523,N_3236);
nor U4933 (N_4933,N_4482,N_3006);
nor U4934 (N_4934,N_3535,N_3228);
nand U4935 (N_4935,N_4042,N_3384);
and U4936 (N_4936,N_3392,N_3696);
or U4937 (N_4937,N_3933,N_3378);
and U4938 (N_4938,N_3148,N_4236);
and U4939 (N_4939,N_3303,N_3186);
and U4940 (N_4940,N_3232,N_3797);
nor U4941 (N_4941,N_4409,N_4082);
nand U4942 (N_4942,N_3037,N_3677);
or U4943 (N_4943,N_3703,N_3177);
xnor U4944 (N_4944,N_3748,N_3960);
and U4945 (N_4945,N_3994,N_4112);
nor U4946 (N_4946,N_4191,N_3044);
nand U4947 (N_4947,N_4027,N_3344);
and U4948 (N_4948,N_3365,N_4037);
and U4949 (N_4949,N_4205,N_3257);
nor U4950 (N_4950,N_3549,N_4013);
nor U4951 (N_4951,N_4343,N_4485);
nor U4952 (N_4952,N_4166,N_3078);
or U4953 (N_4953,N_3316,N_3689);
and U4954 (N_4954,N_3826,N_3529);
and U4955 (N_4955,N_3509,N_4008);
and U4956 (N_4956,N_3128,N_3009);
and U4957 (N_4957,N_3070,N_3676);
nor U4958 (N_4958,N_3359,N_3164);
nand U4959 (N_4959,N_4279,N_3978);
nor U4960 (N_4960,N_3283,N_3210);
xor U4961 (N_4961,N_3977,N_4155);
xor U4962 (N_4962,N_4133,N_3871);
nor U4963 (N_4963,N_3955,N_4481);
nand U4964 (N_4964,N_4141,N_3562);
or U4965 (N_4965,N_3420,N_3212);
and U4966 (N_4966,N_3619,N_3435);
nor U4967 (N_4967,N_4120,N_3626);
and U4968 (N_4968,N_3311,N_3750);
or U4969 (N_4969,N_4453,N_4165);
xor U4970 (N_4970,N_3916,N_3780);
or U4971 (N_4971,N_3056,N_3531);
nand U4972 (N_4972,N_4069,N_3014);
nor U4973 (N_4973,N_3673,N_4487);
and U4974 (N_4974,N_4062,N_3223);
nor U4975 (N_4975,N_4014,N_4392);
and U4976 (N_4976,N_3537,N_3343);
nor U4977 (N_4977,N_3168,N_3322);
nand U4978 (N_4978,N_3131,N_3158);
nor U4979 (N_4979,N_3188,N_3161);
and U4980 (N_4980,N_3370,N_3769);
and U4981 (N_4981,N_3875,N_3885);
nand U4982 (N_4982,N_3060,N_3817);
nand U4983 (N_4983,N_4230,N_4308);
nor U4984 (N_4984,N_4156,N_3211);
or U4985 (N_4985,N_3777,N_3727);
nor U4986 (N_4986,N_3289,N_3341);
or U4987 (N_4987,N_3422,N_4493);
or U4988 (N_4988,N_3134,N_3313);
nand U4989 (N_4989,N_3431,N_4021);
nor U4990 (N_4990,N_4440,N_3354);
nand U4991 (N_4991,N_4270,N_3940);
nand U4992 (N_4992,N_3828,N_3206);
nor U4993 (N_4993,N_4337,N_3571);
or U4994 (N_4994,N_3273,N_3351);
and U4995 (N_4995,N_4129,N_3876);
nor U4996 (N_4996,N_4277,N_4369);
nor U4997 (N_4997,N_3642,N_3532);
nor U4998 (N_4998,N_3237,N_3761);
and U4999 (N_4999,N_4484,N_4262);
xnor U5000 (N_5000,N_3307,N_3493);
nand U5001 (N_5001,N_4182,N_4339);
xnor U5002 (N_5002,N_4323,N_3796);
nand U5003 (N_5003,N_4402,N_3708);
nor U5004 (N_5004,N_3495,N_4371);
or U5005 (N_5005,N_4159,N_4019);
xor U5006 (N_5006,N_4436,N_3418);
nor U5007 (N_5007,N_3734,N_3565);
nand U5008 (N_5008,N_3931,N_4130);
nor U5009 (N_5009,N_3361,N_3637);
and U5010 (N_5010,N_3782,N_3966);
and U5011 (N_5011,N_3788,N_4358);
xnor U5012 (N_5012,N_3156,N_4292);
and U5013 (N_5013,N_3594,N_4047);
nand U5014 (N_5014,N_3577,N_3046);
nand U5015 (N_5015,N_4331,N_3524);
or U5016 (N_5016,N_3711,N_3892);
and U5017 (N_5017,N_4329,N_4416);
and U5018 (N_5018,N_3254,N_4058);
nand U5019 (N_5019,N_4017,N_4018);
and U5020 (N_5020,N_4204,N_3805);
and U5021 (N_5021,N_3635,N_4015);
nand U5022 (N_5022,N_3759,N_3829);
and U5023 (N_5023,N_4408,N_3130);
nand U5024 (N_5024,N_4391,N_3946);
or U5025 (N_5025,N_3020,N_3965);
or U5026 (N_5026,N_3329,N_4427);
or U5027 (N_5027,N_3636,N_4106);
or U5028 (N_5028,N_4103,N_4227);
nor U5029 (N_5029,N_4090,N_4425);
and U5030 (N_5030,N_4271,N_3850);
nor U5031 (N_5031,N_3720,N_3146);
nor U5032 (N_5032,N_3956,N_3884);
xor U5033 (N_5033,N_3101,N_3737);
and U5034 (N_5034,N_3880,N_4109);
xnor U5035 (N_5035,N_3507,N_3941);
or U5036 (N_5036,N_3488,N_3285);
nand U5037 (N_5037,N_3921,N_3314);
nor U5038 (N_5038,N_3649,N_4488);
or U5039 (N_5039,N_3299,N_4368);
or U5040 (N_5040,N_3201,N_4477);
nand U5041 (N_5041,N_3360,N_3976);
nor U5042 (N_5042,N_3159,N_3859);
nand U5043 (N_5043,N_4253,N_4411);
nand U5044 (N_5044,N_3647,N_4298);
or U5045 (N_5045,N_3633,N_3356);
nor U5046 (N_5046,N_4043,N_3760);
and U5047 (N_5047,N_3225,N_3587);
nand U5048 (N_5048,N_3611,N_3385);
xnor U5049 (N_5049,N_3784,N_4437);
nand U5050 (N_5050,N_4458,N_3487);
nand U5051 (N_5051,N_4387,N_3586);
or U5052 (N_5052,N_3559,N_3740);
nand U5053 (N_5053,N_4185,N_3858);
and U5054 (N_5054,N_3566,N_4220);
nor U5055 (N_5055,N_4309,N_3057);
nor U5056 (N_5056,N_3376,N_3890);
and U5057 (N_5057,N_3516,N_3085);
nor U5058 (N_5058,N_3315,N_3401);
xnor U5059 (N_5059,N_3490,N_3621);
nand U5060 (N_5060,N_3318,N_3095);
and U5061 (N_5061,N_4459,N_3489);
nor U5062 (N_5062,N_3058,N_3068);
and U5063 (N_5063,N_3452,N_3867);
nor U5064 (N_5064,N_3194,N_4097);
nand U5065 (N_5065,N_3451,N_3550);
nand U5066 (N_5066,N_3262,N_3609);
or U5067 (N_5067,N_3951,N_3157);
nor U5068 (N_5068,N_3373,N_3541);
and U5069 (N_5069,N_3199,N_3333);
or U5070 (N_5070,N_3375,N_3176);
xor U5071 (N_5071,N_4243,N_3835);
nand U5072 (N_5072,N_3007,N_3442);
or U5073 (N_5073,N_4144,N_3012);
and U5074 (N_5074,N_4232,N_3857);
nand U5075 (N_5075,N_3379,N_3888);
or U5076 (N_5076,N_3038,N_3208);
nor U5077 (N_5077,N_3866,N_3856);
nor U5078 (N_5078,N_4061,N_4059);
and U5079 (N_5079,N_3764,N_3286);
nor U5080 (N_5080,N_3229,N_4350);
or U5081 (N_5081,N_3353,N_4455);
nor U5082 (N_5082,N_3271,N_3011);
and U5083 (N_5083,N_3485,N_4003);
and U5084 (N_5084,N_4495,N_3430);
nor U5085 (N_5085,N_3971,N_4274);
and U5086 (N_5086,N_4394,N_3424);
nand U5087 (N_5087,N_3848,N_3276);
nand U5088 (N_5088,N_3680,N_4020);
nand U5089 (N_5089,N_3092,N_3839);
nand U5090 (N_5090,N_4009,N_3906);
nand U5091 (N_5091,N_3259,N_3105);
and U5092 (N_5092,N_4153,N_4344);
or U5093 (N_5093,N_3534,N_3411);
and U5094 (N_5094,N_4451,N_4258);
and U5095 (N_5095,N_4050,N_4216);
and U5096 (N_5096,N_3387,N_3799);
or U5097 (N_5097,N_3954,N_3834);
and U5098 (N_5098,N_4086,N_3240);
nand U5099 (N_5099,N_3950,N_3664);
nor U5100 (N_5100,N_4335,N_3366);
xor U5101 (N_5101,N_4413,N_4007);
xnor U5102 (N_5102,N_3898,N_3357);
and U5103 (N_5103,N_4378,N_3580);
nand U5104 (N_5104,N_3903,N_3979);
xor U5105 (N_5105,N_3803,N_4148);
nand U5106 (N_5106,N_3717,N_3395);
xnor U5107 (N_5107,N_4046,N_3631);
nor U5108 (N_5108,N_4076,N_3081);
and U5109 (N_5109,N_3477,N_3371);
xor U5110 (N_5110,N_3970,N_4385);
and U5111 (N_5111,N_4260,N_3419);
or U5112 (N_5112,N_4184,N_3973);
or U5113 (N_5113,N_3331,N_3358);
and U5114 (N_5114,N_4435,N_3787);
and U5115 (N_5115,N_3466,N_4388);
nor U5116 (N_5116,N_4240,N_4064);
nor U5117 (N_5117,N_4203,N_3072);
nor U5118 (N_5118,N_4483,N_3684);
nor U5119 (N_5119,N_3015,N_3382);
nand U5120 (N_5120,N_4444,N_4356);
xnor U5121 (N_5121,N_3807,N_4095);
and U5122 (N_5122,N_4134,N_3794);
and U5123 (N_5123,N_3686,N_4380);
or U5124 (N_5124,N_3768,N_3197);
and U5125 (N_5125,N_3233,N_4412);
and U5126 (N_5126,N_3793,N_3578);
and U5127 (N_5127,N_3515,N_3217);
nand U5128 (N_5128,N_3239,N_3719);
nand U5129 (N_5129,N_3713,N_4023);
and U5130 (N_5130,N_4423,N_4472);
and U5131 (N_5131,N_3140,N_3671);
nand U5132 (N_5132,N_4265,N_4075);
nand U5133 (N_5133,N_4353,N_4151);
or U5134 (N_5134,N_3809,N_3667);
nor U5135 (N_5135,N_3881,N_3910);
and U5136 (N_5136,N_3324,N_3539);
and U5137 (N_5137,N_4496,N_3712);
nand U5138 (N_5138,N_4004,N_3646);
or U5139 (N_5139,N_4195,N_4338);
nor U5140 (N_5140,N_3052,N_4489);
nor U5141 (N_5141,N_3099,N_3919);
nand U5142 (N_5142,N_3891,N_3222);
and U5143 (N_5143,N_3414,N_3417);
nor U5144 (N_5144,N_3579,N_3335);
nand U5145 (N_5145,N_3347,N_4386);
and U5146 (N_5146,N_3842,N_3821);
or U5147 (N_5147,N_4281,N_4001);
and U5148 (N_5148,N_3256,N_3294);
nand U5149 (N_5149,N_4432,N_3570);
nand U5150 (N_5150,N_3658,N_3968);
or U5151 (N_5151,N_4430,N_3900);
or U5152 (N_5152,N_3783,N_3902);
nor U5153 (N_5153,N_3268,N_3672);
nand U5154 (N_5154,N_3655,N_3407);
nand U5155 (N_5155,N_3986,N_3434);
or U5156 (N_5156,N_4135,N_3269);
or U5157 (N_5157,N_3119,N_3183);
nand U5158 (N_5158,N_4283,N_3325);
and U5159 (N_5159,N_3520,N_3909);
or U5160 (N_5160,N_3393,N_3563);
nor U5161 (N_5161,N_4012,N_3825);
nand U5162 (N_5162,N_3319,N_3926);
and U5163 (N_5163,N_3486,N_4233);
nand U5164 (N_5164,N_3270,N_4071);
nor U5165 (N_5165,N_3975,N_4235);
nand U5166 (N_5166,N_3412,N_3204);
xnor U5167 (N_5167,N_4326,N_3691);
or U5168 (N_5168,N_3115,N_3446);
and U5169 (N_5169,N_4102,N_4199);
and U5170 (N_5170,N_3097,N_4327);
nand U5171 (N_5171,N_4422,N_4441);
and U5172 (N_5172,N_3517,N_4439);
and U5173 (N_5173,N_4320,N_3491);
and U5174 (N_5174,N_4176,N_3340);
and U5175 (N_5175,N_3984,N_4322);
nor U5176 (N_5176,N_4087,N_3742);
and U5177 (N_5177,N_3073,N_4055);
nor U5178 (N_5178,N_3969,N_3394);
nand U5179 (N_5179,N_4113,N_4291);
nand U5180 (N_5180,N_3025,N_4067);
nor U5181 (N_5181,N_3139,N_4304);
nor U5182 (N_5182,N_4025,N_4357);
or U5183 (N_5183,N_4420,N_3251);
or U5184 (N_5184,N_3924,N_3860);
and U5185 (N_5185,N_3458,N_4162);
and U5186 (N_5186,N_4002,N_3625);
or U5187 (N_5187,N_3945,N_3221);
and U5188 (N_5188,N_3172,N_3103);
or U5189 (N_5189,N_3292,N_3249);
nand U5190 (N_5190,N_3679,N_3166);
xnor U5191 (N_5191,N_3786,N_3685);
nand U5192 (N_5192,N_3321,N_3872);
nor U5193 (N_5193,N_3653,N_3630);
nor U5194 (N_5194,N_3352,N_4225);
nand U5195 (N_5195,N_3248,N_4438);
and U5196 (N_5196,N_4079,N_3540);
xor U5197 (N_5197,N_3142,N_3996);
nand U5198 (N_5198,N_4272,N_4461);
nand U5199 (N_5199,N_4486,N_3795);
nor U5200 (N_5200,N_3640,N_3682);
xor U5201 (N_5201,N_3282,N_3558);
nand U5202 (N_5202,N_3600,N_3291);
and U5203 (N_5203,N_3429,N_4150);
and U5204 (N_5204,N_3400,N_3389);
or U5205 (N_5205,N_3622,N_3738);
nand U5206 (N_5206,N_3775,N_3503);
nand U5207 (N_5207,N_3136,N_3824);
or U5208 (N_5208,N_3061,N_3162);
nand U5209 (N_5209,N_3791,N_3005);
nor U5210 (N_5210,N_3310,N_3178);
and U5211 (N_5211,N_4284,N_4497);
nor U5212 (N_5212,N_3459,N_4346);
nand U5213 (N_5213,N_3937,N_4035);
and U5214 (N_5214,N_3721,N_4089);
nand U5215 (N_5215,N_3182,N_4334);
xor U5216 (N_5216,N_4450,N_3165);
and U5217 (N_5217,N_4401,N_4218);
nand U5218 (N_5218,N_3355,N_4319);
xnor U5219 (N_5219,N_3484,N_4063);
and U5220 (N_5220,N_4457,N_4092);
nand U5221 (N_5221,N_4238,N_3861);
nor U5222 (N_5222,N_4173,N_4447);
nand U5223 (N_5223,N_4454,N_3944);
or U5224 (N_5224,N_3302,N_4048);
and U5225 (N_5225,N_3246,N_3936);
and U5226 (N_5226,N_3723,N_3235);
nor U5227 (N_5227,N_4252,N_4456);
and U5228 (N_5228,N_3213,N_3798);
and U5229 (N_5229,N_4359,N_4215);
and U5230 (N_5230,N_4200,N_3776);
xnor U5231 (N_5231,N_4100,N_3665);
and U5232 (N_5232,N_3743,N_3603);
nand U5233 (N_5233,N_4005,N_4224);
or U5234 (N_5234,N_4273,N_3889);
nand U5235 (N_5235,N_4110,N_4499);
nor U5236 (N_5236,N_3267,N_3067);
and U5237 (N_5237,N_4101,N_4480);
or U5238 (N_5238,N_3308,N_3363);
nand U5239 (N_5239,N_3707,N_4137);
or U5240 (N_5240,N_3479,N_3444);
nor U5241 (N_5241,N_4306,N_4098);
xor U5242 (N_5242,N_4302,N_4212);
nand U5243 (N_5243,N_3181,N_3747);
nor U5244 (N_5244,N_3583,N_4105);
nor U5245 (N_5245,N_4036,N_3993);
and U5246 (N_5246,N_3730,N_4072);
nand U5247 (N_5247,N_3901,N_3175);
nand U5248 (N_5248,N_4313,N_3002);
nor U5249 (N_5249,N_4239,N_3170);
or U5250 (N_5250,N_3127,N_4309);
or U5251 (N_5251,N_4285,N_3834);
nand U5252 (N_5252,N_3375,N_4113);
nand U5253 (N_5253,N_4142,N_3817);
nand U5254 (N_5254,N_3565,N_3796);
xor U5255 (N_5255,N_3448,N_4488);
xnor U5256 (N_5256,N_3529,N_4215);
nor U5257 (N_5257,N_4274,N_4049);
nor U5258 (N_5258,N_3385,N_3051);
nor U5259 (N_5259,N_4377,N_3757);
xor U5260 (N_5260,N_3947,N_3091);
and U5261 (N_5261,N_4129,N_3789);
or U5262 (N_5262,N_3823,N_4415);
or U5263 (N_5263,N_3846,N_3313);
and U5264 (N_5264,N_4307,N_4406);
and U5265 (N_5265,N_3684,N_3821);
nor U5266 (N_5266,N_4125,N_3813);
or U5267 (N_5267,N_3346,N_3389);
and U5268 (N_5268,N_3592,N_3962);
and U5269 (N_5269,N_4040,N_3064);
and U5270 (N_5270,N_3821,N_4269);
and U5271 (N_5271,N_3490,N_3830);
nor U5272 (N_5272,N_3303,N_3565);
and U5273 (N_5273,N_3026,N_3856);
nand U5274 (N_5274,N_3749,N_3998);
nor U5275 (N_5275,N_3393,N_3138);
or U5276 (N_5276,N_3808,N_4091);
nor U5277 (N_5277,N_4489,N_3915);
and U5278 (N_5278,N_3041,N_4098);
and U5279 (N_5279,N_4423,N_4082);
or U5280 (N_5280,N_3335,N_4328);
xnor U5281 (N_5281,N_4154,N_4429);
and U5282 (N_5282,N_3861,N_3235);
xor U5283 (N_5283,N_4373,N_3559);
and U5284 (N_5284,N_3988,N_3128);
or U5285 (N_5285,N_3121,N_4305);
nand U5286 (N_5286,N_3504,N_4306);
and U5287 (N_5287,N_4285,N_3324);
and U5288 (N_5288,N_3919,N_3868);
or U5289 (N_5289,N_4034,N_3039);
nand U5290 (N_5290,N_4273,N_3871);
nand U5291 (N_5291,N_4411,N_3257);
xnor U5292 (N_5292,N_3400,N_4045);
and U5293 (N_5293,N_3571,N_3948);
nor U5294 (N_5294,N_3229,N_3994);
xnor U5295 (N_5295,N_4470,N_3801);
nor U5296 (N_5296,N_3895,N_4012);
nand U5297 (N_5297,N_3086,N_3871);
and U5298 (N_5298,N_3381,N_4105);
and U5299 (N_5299,N_4286,N_3542);
or U5300 (N_5300,N_3962,N_4334);
nor U5301 (N_5301,N_4365,N_3511);
or U5302 (N_5302,N_4491,N_3135);
nand U5303 (N_5303,N_3477,N_4223);
nand U5304 (N_5304,N_4314,N_4122);
nor U5305 (N_5305,N_3514,N_3523);
nand U5306 (N_5306,N_3435,N_4286);
nand U5307 (N_5307,N_3157,N_4492);
nand U5308 (N_5308,N_3582,N_3951);
nor U5309 (N_5309,N_4224,N_4253);
nor U5310 (N_5310,N_4334,N_3540);
xor U5311 (N_5311,N_3965,N_4399);
nor U5312 (N_5312,N_4460,N_4447);
nand U5313 (N_5313,N_3611,N_3227);
or U5314 (N_5314,N_3706,N_3868);
and U5315 (N_5315,N_3295,N_3662);
nor U5316 (N_5316,N_3252,N_3657);
nor U5317 (N_5317,N_4409,N_3615);
nand U5318 (N_5318,N_3590,N_4469);
or U5319 (N_5319,N_3665,N_4466);
nor U5320 (N_5320,N_3339,N_3269);
or U5321 (N_5321,N_3917,N_4468);
nand U5322 (N_5322,N_4446,N_3345);
and U5323 (N_5323,N_3054,N_4107);
or U5324 (N_5324,N_3580,N_3667);
nor U5325 (N_5325,N_3234,N_3302);
and U5326 (N_5326,N_3025,N_4123);
nor U5327 (N_5327,N_3402,N_4176);
and U5328 (N_5328,N_3425,N_3279);
nand U5329 (N_5329,N_4319,N_4402);
nor U5330 (N_5330,N_4230,N_4282);
and U5331 (N_5331,N_3685,N_3403);
nor U5332 (N_5332,N_3433,N_4038);
nand U5333 (N_5333,N_3022,N_3543);
or U5334 (N_5334,N_4367,N_3961);
nor U5335 (N_5335,N_3669,N_4112);
and U5336 (N_5336,N_3732,N_4101);
or U5337 (N_5337,N_3514,N_4022);
nand U5338 (N_5338,N_3275,N_3311);
and U5339 (N_5339,N_4196,N_3174);
nand U5340 (N_5340,N_3801,N_3277);
nor U5341 (N_5341,N_3466,N_3933);
or U5342 (N_5342,N_3335,N_3831);
xnor U5343 (N_5343,N_3797,N_3826);
and U5344 (N_5344,N_4083,N_3746);
and U5345 (N_5345,N_4304,N_4077);
nand U5346 (N_5346,N_3652,N_3477);
and U5347 (N_5347,N_3557,N_3908);
nand U5348 (N_5348,N_4406,N_3228);
xor U5349 (N_5349,N_3918,N_4305);
or U5350 (N_5350,N_3774,N_3604);
and U5351 (N_5351,N_3279,N_3992);
xor U5352 (N_5352,N_3590,N_3779);
and U5353 (N_5353,N_3918,N_4172);
and U5354 (N_5354,N_3014,N_3939);
or U5355 (N_5355,N_3253,N_3652);
nor U5356 (N_5356,N_3223,N_3777);
and U5357 (N_5357,N_3036,N_3765);
nand U5358 (N_5358,N_4074,N_3042);
nand U5359 (N_5359,N_4452,N_3467);
xor U5360 (N_5360,N_4339,N_3293);
and U5361 (N_5361,N_3489,N_3343);
or U5362 (N_5362,N_3112,N_4487);
nand U5363 (N_5363,N_4393,N_3748);
and U5364 (N_5364,N_3322,N_3207);
and U5365 (N_5365,N_4245,N_3668);
nand U5366 (N_5366,N_4259,N_3416);
nand U5367 (N_5367,N_3882,N_3948);
or U5368 (N_5368,N_3679,N_3364);
nand U5369 (N_5369,N_4125,N_3190);
or U5370 (N_5370,N_3562,N_3199);
xor U5371 (N_5371,N_3643,N_4188);
and U5372 (N_5372,N_3456,N_4331);
or U5373 (N_5373,N_3859,N_3762);
nor U5374 (N_5374,N_4329,N_3109);
nor U5375 (N_5375,N_3405,N_4234);
nand U5376 (N_5376,N_3347,N_4196);
xnor U5377 (N_5377,N_4251,N_3752);
and U5378 (N_5378,N_3968,N_4221);
xor U5379 (N_5379,N_4403,N_4106);
nand U5380 (N_5380,N_3392,N_4454);
nand U5381 (N_5381,N_4032,N_4390);
nand U5382 (N_5382,N_3620,N_4130);
nor U5383 (N_5383,N_3763,N_3040);
or U5384 (N_5384,N_3627,N_3796);
nand U5385 (N_5385,N_3146,N_3019);
and U5386 (N_5386,N_3401,N_4101);
or U5387 (N_5387,N_4027,N_3322);
nor U5388 (N_5388,N_3117,N_4246);
nand U5389 (N_5389,N_3008,N_4131);
nor U5390 (N_5390,N_4013,N_3627);
or U5391 (N_5391,N_3381,N_3552);
and U5392 (N_5392,N_3210,N_4397);
nor U5393 (N_5393,N_3949,N_3655);
nor U5394 (N_5394,N_4482,N_3590);
or U5395 (N_5395,N_3791,N_3700);
and U5396 (N_5396,N_3589,N_3442);
nor U5397 (N_5397,N_3819,N_3553);
nand U5398 (N_5398,N_4317,N_3541);
xor U5399 (N_5399,N_3274,N_3978);
nor U5400 (N_5400,N_3290,N_3220);
nand U5401 (N_5401,N_3925,N_4228);
and U5402 (N_5402,N_3941,N_3461);
and U5403 (N_5403,N_3888,N_3350);
nor U5404 (N_5404,N_3087,N_3803);
nor U5405 (N_5405,N_4066,N_3152);
nor U5406 (N_5406,N_4348,N_3315);
and U5407 (N_5407,N_3033,N_3957);
nand U5408 (N_5408,N_4088,N_3208);
nand U5409 (N_5409,N_3243,N_3092);
and U5410 (N_5410,N_3702,N_4183);
or U5411 (N_5411,N_3546,N_3739);
nor U5412 (N_5412,N_3428,N_3679);
nand U5413 (N_5413,N_3637,N_3082);
xnor U5414 (N_5414,N_3600,N_3403);
nand U5415 (N_5415,N_4006,N_3537);
nor U5416 (N_5416,N_3852,N_3596);
nor U5417 (N_5417,N_3307,N_4095);
nand U5418 (N_5418,N_3539,N_3957);
or U5419 (N_5419,N_3923,N_3451);
and U5420 (N_5420,N_3311,N_3458);
and U5421 (N_5421,N_4422,N_3080);
xnor U5422 (N_5422,N_4458,N_3814);
nor U5423 (N_5423,N_3149,N_4468);
nor U5424 (N_5424,N_4439,N_3963);
and U5425 (N_5425,N_4295,N_3622);
or U5426 (N_5426,N_3417,N_4302);
or U5427 (N_5427,N_3129,N_4489);
or U5428 (N_5428,N_3606,N_3263);
nand U5429 (N_5429,N_4333,N_3171);
and U5430 (N_5430,N_4369,N_4441);
and U5431 (N_5431,N_3240,N_4103);
and U5432 (N_5432,N_3202,N_4284);
xnor U5433 (N_5433,N_3499,N_4140);
nand U5434 (N_5434,N_3514,N_4396);
and U5435 (N_5435,N_3115,N_4189);
nand U5436 (N_5436,N_3124,N_4436);
nor U5437 (N_5437,N_3460,N_3179);
nor U5438 (N_5438,N_3789,N_4028);
and U5439 (N_5439,N_4077,N_3035);
nor U5440 (N_5440,N_3028,N_4456);
nand U5441 (N_5441,N_3310,N_3977);
and U5442 (N_5442,N_3560,N_3874);
or U5443 (N_5443,N_3721,N_3746);
or U5444 (N_5444,N_4142,N_4350);
xnor U5445 (N_5445,N_4423,N_3861);
or U5446 (N_5446,N_4055,N_3324);
nor U5447 (N_5447,N_4453,N_4160);
nor U5448 (N_5448,N_3189,N_4291);
xor U5449 (N_5449,N_3511,N_3994);
or U5450 (N_5450,N_3449,N_4486);
and U5451 (N_5451,N_4319,N_4409);
and U5452 (N_5452,N_3276,N_3135);
or U5453 (N_5453,N_3301,N_4403);
and U5454 (N_5454,N_3044,N_3300);
nand U5455 (N_5455,N_4371,N_3551);
nor U5456 (N_5456,N_4417,N_3912);
nand U5457 (N_5457,N_4394,N_3836);
nand U5458 (N_5458,N_4233,N_4084);
and U5459 (N_5459,N_3716,N_4481);
nor U5460 (N_5460,N_3266,N_3115);
and U5461 (N_5461,N_4358,N_4262);
or U5462 (N_5462,N_3581,N_3717);
nor U5463 (N_5463,N_4055,N_3409);
and U5464 (N_5464,N_3675,N_4430);
nor U5465 (N_5465,N_4257,N_3939);
and U5466 (N_5466,N_3213,N_3121);
and U5467 (N_5467,N_3598,N_3157);
nand U5468 (N_5468,N_3639,N_4466);
nor U5469 (N_5469,N_4499,N_4473);
nand U5470 (N_5470,N_4392,N_4379);
nand U5471 (N_5471,N_3856,N_3786);
xnor U5472 (N_5472,N_3284,N_3829);
or U5473 (N_5473,N_4389,N_3992);
or U5474 (N_5474,N_3970,N_4070);
and U5475 (N_5475,N_3101,N_3162);
or U5476 (N_5476,N_3397,N_4312);
nand U5477 (N_5477,N_4331,N_3656);
or U5478 (N_5478,N_3255,N_3893);
nand U5479 (N_5479,N_3020,N_3178);
nand U5480 (N_5480,N_3593,N_4275);
nor U5481 (N_5481,N_4308,N_4142);
nand U5482 (N_5482,N_4357,N_3974);
nor U5483 (N_5483,N_4454,N_3368);
and U5484 (N_5484,N_4253,N_4430);
nand U5485 (N_5485,N_3739,N_3399);
and U5486 (N_5486,N_3598,N_4198);
or U5487 (N_5487,N_3623,N_3943);
and U5488 (N_5488,N_4071,N_3562);
nor U5489 (N_5489,N_3789,N_3654);
and U5490 (N_5490,N_4165,N_3816);
xnor U5491 (N_5491,N_3702,N_3239);
xor U5492 (N_5492,N_3825,N_3358);
and U5493 (N_5493,N_3335,N_3669);
or U5494 (N_5494,N_3107,N_3328);
and U5495 (N_5495,N_3285,N_4465);
or U5496 (N_5496,N_3536,N_3921);
nand U5497 (N_5497,N_4350,N_3493);
nor U5498 (N_5498,N_3010,N_3193);
or U5499 (N_5499,N_3546,N_3157);
or U5500 (N_5500,N_4438,N_3789);
or U5501 (N_5501,N_4275,N_3519);
nor U5502 (N_5502,N_3164,N_4008);
or U5503 (N_5503,N_3802,N_3554);
nand U5504 (N_5504,N_3833,N_4066);
and U5505 (N_5505,N_3774,N_4026);
xnor U5506 (N_5506,N_3481,N_3532);
nor U5507 (N_5507,N_3244,N_3012);
nor U5508 (N_5508,N_3682,N_3756);
or U5509 (N_5509,N_4407,N_4464);
xnor U5510 (N_5510,N_3698,N_4250);
xor U5511 (N_5511,N_3796,N_3868);
and U5512 (N_5512,N_3524,N_3067);
nand U5513 (N_5513,N_4234,N_4031);
and U5514 (N_5514,N_3926,N_3621);
nor U5515 (N_5515,N_3222,N_3800);
or U5516 (N_5516,N_4466,N_3758);
or U5517 (N_5517,N_3288,N_4070);
nand U5518 (N_5518,N_3485,N_3773);
or U5519 (N_5519,N_4436,N_3129);
nand U5520 (N_5520,N_4188,N_3707);
or U5521 (N_5521,N_3380,N_3606);
nor U5522 (N_5522,N_3532,N_3674);
nand U5523 (N_5523,N_3650,N_4403);
or U5524 (N_5524,N_4105,N_4051);
and U5525 (N_5525,N_4489,N_3037);
and U5526 (N_5526,N_4481,N_3506);
nor U5527 (N_5527,N_3440,N_4106);
xnor U5528 (N_5528,N_3856,N_4027);
xnor U5529 (N_5529,N_4238,N_4026);
or U5530 (N_5530,N_4011,N_4322);
nor U5531 (N_5531,N_3329,N_3476);
xnor U5532 (N_5532,N_3011,N_3086);
and U5533 (N_5533,N_3282,N_4158);
and U5534 (N_5534,N_3541,N_3292);
or U5535 (N_5535,N_4169,N_4476);
nor U5536 (N_5536,N_3726,N_3664);
or U5537 (N_5537,N_3860,N_4018);
xnor U5538 (N_5538,N_3722,N_4396);
xor U5539 (N_5539,N_3022,N_4077);
or U5540 (N_5540,N_3524,N_3867);
or U5541 (N_5541,N_3028,N_4086);
nor U5542 (N_5542,N_3440,N_4451);
xnor U5543 (N_5543,N_3605,N_3085);
nor U5544 (N_5544,N_3487,N_4188);
xor U5545 (N_5545,N_3089,N_3140);
nor U5546 (N_5546,N_4187,N_4465);
or U5547 (N_5547,N_4402,N_3649);
or U5548 (N_5548,N_3306,N_3970);
or U5549 (N_5549,N_4386,N_4433);
or U5550 (N_5550,N_3089,N_3670);
xnor U5551 (N_5551,N_3373,N_3177);
or U5552 (N_5552,N_3593,N_4303);
and U5553 (N_5553,N_3772,N_3960);
and U5554 (N_5554,N_3002,N_3118);
and U5555 (N_5555,N_3800,N_4215);
or U5556 (N_5556,N_3039,N_4231);
or U5557 (N_5557,N_3416,N_3035);
nor U5558 (N_5558,N_3626,N_3817);
nor U5559 (N_5559,N_3980,N_3692);
nor U5560 (N_5560,N_3311,N_3066);
nand U5561 (N_5561,N_3343,N_3346);
or U5562 (N_5562,N_3710,N_3637);
nor U5563 (N_5563,N_4150,N_3866);
nor U5564 (N_5564,N_4417,N_4023);
or U5565 (N_5565,N_3535,N_3391);
nand U5566 (N_5566,N_4226,N_4006);
and U5567 (N_5567,N_3552,N_3558);
xor U5568 (N_5568,N_4352,N_4439);
and U5569 (N_5569,N_3080,N_3032);
nand U5570 (N_5570,N_4293,N_3265);
or U5571 (N_5571,N_3343,N_3280);
xor U5572 (N_5572,N_4469,N_4436);
nor U5573 (N_5573,N_3945,N_4422);
or U5574 (N_5574,N_3737,N_3775);
xnor U5575 (N_5575,N_3473,N_4363);
nand U5576 (N_5576,N_4390,N_4295);
and U5577 (N_5577,N_4116,N_3455);
nand U5578 (N_5578,N_3136,N_3944);
or U5579 (N_5579,N_4123,N_4172);
and U5580 (N_5580,N_3874,N_3508);
nand U5581 (N_5581,N_4189,N_3941);
nand U5582 (N_5582,N_3412,N_3208);
or U5583 (N_5583,N_4021,N_4027);
nand U5584 (N_5584,N_4118,N_3881);
and U5585 (N_5585,N_3887,N_3004);
nand U5586 (N_5586,N_4262,N_3622);
xnor U5587 (N_5587,N_3463,N_4436);
and U5588 (N_5588,N_3159,N_3002);
nor U5589 (N_5589,N_3637,N_3859);
or U5590 (N_5590,N_3034,N_3180);
xnor U5591 (N_5591,N_3395,N_3497);
or U5592 (N_5592,N_3174,N_3009);
nand U5593 (N_5593,N_3973,N_3226);
nand U5594 (N_5594,N_4493,N_4461);
and U5595 (N_5595,N_3193,N_3371);
and U5596 (N_5596,N_4177,N_3088);
nand U5597 (N_5597,N_4483,N_3809);
nand U5598 (N_5598,N_3548,N_4216);
nor U5599 (N_5599,N_4122,N_4362);
xnor U5600 (N_5600,N_4188,N_3151);
nand U5601 (N_5601,N_3728,N_3144);
nor U5602 (N_5602,N_3603,N_3744);
nor U5603 (N_5603,N_3237,N_4432);
or U5604 (N_5604,N_4080,N_4209);
nand U5605 (N_5605,N_3619,N_4487);
and U5606 (N_5606,N_4134,N_4467);
nand U5607 (N_5607,N_3725,N_3963);
and U5608 (N_5608,N_4300,N_3278);
nand U5609 (N_5609,N_4275,N_4003);
and U5610 (N_5610,N_4327,N_3952);
and U5611 (N_5611,N_4497,N_3112);
nand U5612 (N_5612,N_3760,N_4469);
or U5613 (N_5613,N_3195,N_4474);
nor U5614 (N_5614,N_3676,N_3820);
nand U5615 (N_5615,N_4122,N_3587);
and U5616 (N_5616,N_3566,N_4238);
nand U5617 (N_5617,N_3040,N_3116);
and U5618 (N_5618,N_3876,N_3498);
nand U5619 (N_5619,N_3670,N_4451);
or U5620 (N_5620,N_3497,N_3454);
and U5621 (N_5621,N_4155,N_4419);
xor U5622 (N_5622,N_4095,N_4179);
nand U5623 (N_5623,N_4314,N_4081);
nand U5624 (N_5624,N_4369,N_4481);
or U5625 (N_5625,N_4105,N_3810);
nand U5626 (N_5626,N_4468,N_4050);
nand U5627 (N_5627,N_3665,N_4074);
or U5628 (N_5628,N_3918,N_3941);
nor U5629 (N_5629,N_4272,N_4447);
or U5630 (N_5630,N_3160,N_4249);
and U5631 (N_5631,N_4351,N_4041);
nor U5632 (N_5632,N_4296,N_4429);
xnor U5633 (N_5633,N_4040,N_4141);
and U5634 (N_5634,N_3939,N_3121);
or U5635 (N_5635,N_4184,N_4191);
nor U5636 (N_5636,N_3397,N_3138);
or U5637 (N_5637,N_3368,N_3631);
or U5638 (N_5638,N_4051,N_3772);
nor U5639 (N_5639,N_3089,N_3194);
nand U5640 (N_5640,N_3574,N_3428);
or U5641 (N_5641,N_3403,N_3236);
and U5642 (N_5642,N_3630,N_3930);
and U5643 (N_5643,N_3939,N_4313);
nor U5644 (N_5644,N_3246,N_3984);
nand U5645 (N_5645,N_4473,N_4049);
nand U5646 (N_5646,N_4369,N_3627);
nand U5647 (N_5647,N_3917,N_3694);
and U5648 (N_5648,N_3527,N_4022);
nor U5649 (N_5649,N_3545,N_3220);
or U5650 (N_5650,N_4262,N_3253);
nor U5651 (N_5651,N_4019,N_3258);
nor U5652 (N_5652,N_3224,N_3149);
and U5653 (N_5653,N_4241,N_3258);
nor U5654 (N_5654,N_3299,N_3191);
nand U5655 (N_5655,N_3968,N_3879);
nand U5656 (N_5656,N_4138,N_4474);
or U5657 (N_5657,N_3327,N_3545);
or U5658 (N_5658,N_3485,N_4232);
nor U5659 (N_5659,N_3821,N_3678);
nor U5660 (N_5660,N_3865,N_4207);
nand U5661 (N_5661,N_3146,N_4082);
and U5662 (N_5662,N_4462,N_3632);
or U5663 (N_5663,N_3389,N_4033);
and U5664 (N_5664,N_3194,N_3525);
nand U5665 (N_5665,N_3168,N_3856);
nor U5666 (N_5666,N_3027,N_3419);
and U5667 (N_5667,N_3164,N_3044);
or U5668 (N_5668,N_3617,N_3908);
nand U5669 (N_5669,N_3600,N_3591);
nor U5670 (N_5670,N_4429,N_3695);
nor U5671 (N_5671,N_4496,N_3158);
nor U5672 (N_5672,N_4368,N_4079);
or U5673 (N_5673,N_3812,N_4168);
or U5674 (N_5674,N_3695,N_4446);
nand U5675 (N_5675,N_3976,N_4310);
and U5676 (N_5676,N_3521,N_3058);
or U5677 (N_5677,N_4381,N_3026);
nand U5678 (N_5678,N_3901,N_4023);
xor U5679 (N_5679,N_3957,N_3826);
nand U5680 (N_5680,N_4262,N_3426);
nand U5681 (N_5681,N_3098,N_3884);
or U5682 (N_5682,N_4200,N_3908);
and U5683 (N_5683,N_4331,N_3634);
xor U5684 (N_5684,N_4359,N_3951);
or U5685 (N_5685,N_3961,N_4328);
nor U5686 (N_5686,N_4378,N_3076);
nor U5687 (N_5687,N_4122,N_3301);
nand U5688 (N_5688,N_3451,N_4051);
nor U5689 (N_5689,N_3295,N_3008);
nand U5690 (N_5690,N_3577,N_3518);
xor U5691 (N_5691,N_4244,N_3330);
and U5692 (N_5692,N_4098,N_3677);
nor U5693 (N_5693,N_4460,N_3657);
and U5694 (N_5694,N_3635,N_4214);
or U5695 (N_5695,N_3001,N_4485);
nor U5696 (N_5696,N_3102,N_3420);
and U5697 (N_5697,N_4187,N_3406);
or U5698 (N_5698,N_4081,N_3751);
nand U5699 (N_5699,N_3956,N_4495);
nor U5700 (N_5700,N_3736,N_4066);
and U5701 (N_5701,N_3448,N_4218);
xnor U5702 (N_5702,N_3196,N_4182);
nor U5703 (N_5703,N_4418,N_3695);
and U5704 (N_5704,N_3671,N_3550);
and U5705 (N_5705,N_3173,N_3114);
or U5706 (N_5706,N_4098,N_3806);
nand U5707 (N_5707,N_4346,N_4118);
nor U5708 (N_5708,N_3159,N_3282);
nor U5709 (N_5709,N_3089,N_3600);
nand U5710 (N_5710,N_3026,N_3170);
nor U5711 (N_5711,N_4064,N_3885);
nand U5712 (N_5712,N_4479,N_3629);
nand U5713 (N_5713,N_3206,N_3609);
and U5714 (N_5714,N_3995,N_3167);
nand U5715 (N_5715,N_4274,N_4071);
nor U5716 (N_5716,N_4072,N_3771);
or U5717 (N_5717,N_4164,N_3170);
or U5718 (N_5718,N_3785,N_3051);
nand U5719 (N_5719,N_3044,N_3879);
or U5720 (N_5720,N_3812,N_3643);
nand U5721 (N_5721,N_3226,N_4264);
and U5722 (N_5722,N_4147,N_3103);
or U5723 (N_5723,N_3728,N_4377);
nand U5724 (N_5724,N_4401,N_3260);
xnor U5725 (N_5725,N_4252,N_4224);
nor U5726 (N_5726,N_4165,N_4195);
nor U5727 (N_5727,N_3238,N_4073);
or U5728 (N_5728,N_3826,N_3523);
nand U5729 (N_5729,N_3538,N_3174);
and U5730 (N_5730,N_4213,N_3153);
or U5731 (N_5731,N_3371,N_3637);
and U5732 (N_5732,N_3251,N_3417);
or U5733 (N_5733,N_4377,N_4424);
and U5734 (N_5734,N_3341,N_4458);
nor U5735 (N_5735,N_3134,N_4416);
or U5736 (N_5736,N_4096,N_3123);
nor U5737 (N_5737,N_3268,N_3206);
nor U5738 (N_5738,N_3697,N_4143);
and U5739 (N_5739,N_3023,N_4191);
nor U5740 (N_5740,N_4166,N_3647);
nor U5741 (N_5741,N_3741,N_3191);
nand U5742 (N_5742,N_3296,N_4210);
or U5743 (N_5743,N_4277,N_3167);
xor U5744 (N_5744,N_4050,N_4287);
or U5745 (N_5745,N_3967,N_3139);
and U5746 (N_5746,N_3386,N_4019);
nand U5747 (N_5747,N_3798,N_3445);
and U5748 (N_5748,N_4316,N_4190);
and U5749 (N_5749,N_3838,N_3470);
nand U5750 (N_5750,N_3946,N_3855);
nand U5751 (N_5751,N_4369,N_4143);
xor U5752 (N_5752,N_3846,N_4356);
nor U5753 (N_5753,N_4205,N_3722);
nand U5754 (N_5754,N_3192,N_4286);
or U5755 (N_5755,N_4095,N_3692);
nor U5756 (N_5756,N_4193,N_3783);
and U5757 (N_5757,N_3965,N_4284);
nand U5758 (N_5758,N_3492,N_4452);
and U5759 (N_5759,N_3895,N_3281);
nor U5760 (N_5760,N_4172,N_3635);
or U5761 (N_5761,N_3065,N_4492);
and U5762 (N_5762,N_3788,N_3160);
nand U5763 (N_5763,N_3198,N_3533);
or U5764 (N_5764,N_4305,N_3528);
nor U5765 (N_5765,N_3132,N_3191);
nor U5766 (N_5766,N_3023,N_3021);
nand U5767 (N_5767,N_3731,N_3081);
and U5768 (N_5768,N_3649,N_4480);
xnor U5769 (N_5769,N_3290,N_4383);
nor U5770 (N_5770,N_4119,N_3219);
or U5771 (N_5771,N_4249,N_3367);
and U5772 (N_5772,N_4179,N_3457);
xnor U5773 (N_5773,N_3341,N_3988);
and U5774 (N_5774,N_4452,N_3577);
nand U5775 (N_5775,N_3070,N_4218);
nor U5776 (N_5776,N_4011,N_3214);
nand U5777 (N_5777,N_4032,N_4417);
nor U5778 (N_5778,N_4244,N_3709);
nor U5779 (N_5779,N_3292,N_3950);
nor U5780 (N_5780,N_4145,N_3041);
or U5781 (N_5781,N_4198,N_3699);
and U5782 (N_5782,N_4218,N_3695);
and U5783 (N_5783,N_3717,N_4417);
and U5784 (N_5784,N_3561,N_4472);
nor U5785 (N_5785,N_4361,N_4460);
nand U5786 (N_5786,N_4137,N_3199);
nand U5787 (N_5787,N_4454,N_4158);
nand U5788 (N_5788,N_4156,N_3174);
nand U5789 (N_5789,N_3195,N_3246);
nor U5790 (N_5790,N_4025,N_4200);
nand U5791 (N_5791,N_3799,N_3234);
nand U5792 (N_5792,N_3655,N_3045);
nand U5793 (N_5793,N_4453,N_3692);
and U5794 (N_5794,N_3821,N_3410);
or U5795 (N_5795,N_3153,N_4131);
nor U5796 (N_5796,N_3849,N_4187);
or U5797 (N_5797,N_3213,N_3644);
or U5798 (N_5798,N_3939,N_3947);
or U5799 (N_5799,N_3569,N_3016);
nand U5800 (N_5800,N_3454,N_3882);
nand U5801 (N_5801,N_4130,N_4201);
nor U5802 (N_5802,N_3451,N_3614);
nand U5803 (N_5803,N_4313,N_4448);
or U5804 (N_5804,N_3245,N_4097);
nor U5805 (N_5805,N_3329,N_3651);
and U5806 (N_5806,N_3048,N_3341);
nor U5807 (N_5807,N_4000,N_3824);
or U5808 (N_5808,N_4127,N_4474);
nand U5809 (N_5809,N_3696,N_3860);
nand U5810 (N_5810,N_3634,N_4125);
xnor U5811 (N_5811,N_4161,N_4273);
nand U5812 (N_5812,N_3933,N_3967);
nand U5813 (N_5813,N_3219,N_3763);
and U5814 (N_5814,N_3827,N_4139);
nand U5815 (N_5815,N_4163,N_3197);
nand U5816 (N_5816,N_4353,N_3365);
nor U5817 (N_5817,N_4377,N_4021);
nand U5818 (N_5818,N_3184,N_3099);
nand U5819 (N_5819,N_3406,N_3875);
xnor U5820 (N_5820,N_4078,N_3722);
nand U5821 (N_5821,N_3213,N_3606);
and U5822 (N_5822,N_3698,N_4478);
or U5823 (N_5823,N_4262,N_4241);
or U5824 (N_5824,N_3247,N_4278);
and U5825 (N_5825,N_4273,N_4129);
nor U5826 (N_5826,N_4326,N_4079);
nor U5827 (N_5827,N_3723,N_3472);
xor U5828 (N_5828,N_3021,N_3368);
and U5829 (N_5829,N_4319,N_3910);
nor U5830 (N_5830,N_3125,N_3102);
or U5831 (N_5831,N_3788,N_3046);
and U5832 (N_5832,N_3933,N_3009);
or U5833 (N_5833,N_3947,N_4198);
and U5834 (N_5834,N_4135,N_4153);
nor U5835 (N_5835,N_4133,N_3921);
and U5836 (N_5836,N_3243,N_4200);
nand U5837 (N_5837,N_3196,N_3247);
or U5838 (N_5838,N_3445,N_3982);
and U5839 (N_5839,N_3602,N_4088);
or U5840 (N_5840,N_3998,N_4249);
or U5841 (N_5841,N_3001,N_4111);
nand U5842 (N_5842,N_3956,N_3207);
nor U5843 (N_5843,N_3870,N_4409);
nand U5844 (N_5844,N_3555,N_3370);
nor U5845 (N_5845,N_4199,N_4418);
nor U5846 (N_5846,N_4127,N_4478);
and U5847 (N_5847,N_3481,N_3446);
and U5848 (N_5848,N_3158,N_4385);
nor U5849 (N_5849,N_4226,N_3249);
and U5850 (N_5850,N_3350,N_4177);
and U5851 (N_5851,N_3344,N_3812);
and U5852 (N_5852,N_4182,N_3617);
xnor U5853 (N_5853,N_4212,N_4274);
nand U5854 (N_5854,N_3955,N_3437);
and U5855 (N_5855,N_3215,N_3974);
and U5856 (N_5856,N_3431,N_4490);
or U5857 (N_5857,N_4414,N_3088);
and U5858 (N_5858,N_3660,N_4365);
nand U5859 (N_5859,N_3171,N_3247);
nor U5860 (N_5860,N_4426,N_3772);
nand U5861 (N_5861,N_3796,N_3902);
nor U5862 (N_5862,N_3417,N_4345);
or U5863 (N_5863,N_4441,N_3029);
nor U5864 (N_5864,N_4488,N_3582);
nand U5865 (N_5865,N_4365,N_4003);
nor U5866 (N_5866,N_4407,N_4253);
xor U5867 (N_5867,N_4298,N_3434);
nor U5868 (N_5868,N_3277,N_3180);
or U5869 (N_5869,N_3454,N_4175);
xor U5870 (N_5870,N_4490,N_4488);
and U5871 (N_5871,N_3130,N_4268);
nor U5872 (N_5872,N_3746,N_3366);
or U5873 (N_5873,N_3110,N_3852);
xnor U5874 (N_5874,N_3820,N_3912);
xor U5875 (N_5875,N_3762,N_3937);
nand U5876 (N_5876,N_3322,N_3637);
nand U5877 (N_5877,N_3844,N_3770);
xor U5878 (N_5878,N_4481,N_3424);
xor U5879 (N_5879,N_3828,N_3481);
and U5880 (N_5880,N_3573,N_3333);
and U5881 (N_5881,N_3764,N_4202);
or U5882 (N_5882,N_4025,N_3741);
and U5883 (N_5883,N_3454,N_3416);
nand U5884 (N_5884,N_4023,N_3600);
or U5885 (N_5885,N_3990,N_3267);
or U5886 (N_5886,N_3533,N_4393);
or U5887 (N_5887,N_3334,N_3387);
or U5888 (N_5888,N_3841,N_3511);
xnor U5889 (N_5889,N_3020,N_3132);
or U5890 (N_5890,N_4346,N_3571);
nand U5891 (N_5891,N_4103,N_3401);
nor U5892 (N_5892,N_3382,N_3348);
nand U5893 (N_5893,N_3050,N_3801);
nand U5894 (N_5894,N_4102,N_3351);
and U5895 (N_5895,N_3994,N_4034);
nor U5896 (N_5896,N_4428,N_3752);
and U5897 (N_5897,N_3704,N_4114);
xor U5898 (N_5898,N_4450,N_3576);
nand U5899 (N_5899,N_3376,N_3985);
and U5900 (N_5900,N_3753,N_3844);
and U5901 (N_5901,N_4418,N_4455);
or U5902 (N_5902,N_3404,N_3610);
and U5903 (N_5903,N_3655,N_3595);
nand U5904 (N_5904,N_3099,N_3113);
nor U5905 (N_5905,N_3101,N_3136);
nor U5906 (N_5906,N_3612,N_3355);
and U5907 (N_5907,N_3722,N_3019);
or U5908 (N_5908,N_3085,N_4486);
nand U5909 (N_5909,N_3231,N_4169);
and U5910 (N_5910,N_3109,N_3096);
and U5911 (N_5911,N_3795,N_3222);
and U5912 (N_5912,N_3333,N_3753);
nor U5913 (N_5913,N_4321,N_3608);
nand U5914 (N_5914,N_3090,N_3307);
or U5915 (N_5915,N_3538,N_3797);
and U5916 (N_5916,N_3531,N_4145);
xnor U5917 (N_5917,N_4441,N_3357);
nand U5918 (N_5918,N_3899,N_3891);
or U5919 (N_5919,N_4444,N_3692);
xor U5920 (N_5920,N_3236,N_3735);
or U5921 (N_5921,N_3810,N_4037);
nor U5922 (N_5922,N_4157,N_4016);
nand U5923 (N_5923,N_3765,N_4209);
or U5924 (N_5924,N_3562,N_3481);
nand U5925 (N_5925,N_4206,N_4245);
nand U5926 (N_5926,N_4183,N_3010);
nand U5927 (N_5927,N_4303,N_4291);
and U5928 (N_5928,N_3536,N_4039);
nand U5929 (N_5929,N_3122,N_4338);
and U5930 (N_5930,N_3622,N_4335);
nor U5931 (N_5931,N_4040,N_3522);
nor U5932 (N_5932,N_4450,N_4287);
or U5933 (N_5933,N_3465,N_4117);
nand U5934 (N_5934,N_4499,N_3261);
nand U5935 (N_5935,N_3048,N_3427);
and U5936 (N_5936,N_4132,N_4197);
nand U5937 (N_5937,N_3739,N_3326);
and U5938 (N_5938,N_3325,N_3937);
nor U5939 (N_5939,N_4388,N_3164);
or U5940 (N_5940,N_4064,N_4309);
xnor U5941 (N_5941,N_4255,N_3278);
xor U5942 (N_5942,N_4485,N_3005);
nor U5943 (N_5943,N_4236,N_3881);
nor U5944 (N_5944,N_4293,N_4283);
nand U5945 (N_5945,N_3950,N_3839);
nand U5946 (N_5946,N_3333,N_4144);
xnor U5947 (N_5947,N_3450,N_4330);
and U5948 (N_5948,N_3284,N_4263);
xnor U5949 (N_5949,N_4434,N_3818);
nor U5950 (N_5950,N_3590,N_3561);
nand U5951 (N_5951,N_4143,N_3068);
and U5952 (N_5952,N_4063,N_3848);
nor U5953 (N_5953,N_3330,N_4205);
xor U5954 (N_5954,N_4416,N_4247);
nand U5955 (N_5955,N_4323,N_3672);
nand U5956 (N_5956,N_4218,N_3050);
or U5957 (N_5957,N_4204,N_3703);
xor U5958 (N_5958,N_3996,N_3125);
nand U5959 (N_5959,N_4293,N_4353);
nand U5960 (N_5960,N_3464,N_3411);
or U5961 (N_5961,N_4091,N_3092);
and U5962 (N_5962,N_3383,N_4056);
xnor U5963 (N_5963,N_4420,N_3718);
or U5964 (N_5964,N_4327,N_4166);
nand U5965 (N_5965,N_4381,N_3945);
and U5966 (N_5966,N_3680,N_4284);
and U5967 (N_5967,N_4471,N_3177);
or U5968 (N_5968,N_4170,N_3837);
xnor U5969 (N_5969,N_3090,N_3453);
or U5970 (N_5970,N_3815,N_4297);
nor U5971 (N_5971,N_3271,N_3449);
nor U5972 (N_5972,N_3650,N_3536);
nand U5973 (N_5973,N_3155,N_4154);
nand U5974 (N_5974,N_4182,N_3621);
and U5975 (N_5975,N_3916,N_3760);
and U5976 (N_5976,N_3705,N_3976);
nor U5977 (N_5977,N_4357,N_3312);
nand U5978 (N_5978,N_3955,N_4099);
nand U5979 (N_5979,N_3984,N_4050);
nor U5980 (N_5980,N_4279,N_3255);
nand U5981 (N_5981,N_4280,N_3452);
and U5982 (N_5982,N_3308,N_4060);
nand U5983 (N_5983,N_4030,N_3988);
or U5984 (N_5984,N_4467,N_3506);
xor U5985 (N_5985,N_3032,N_4004);
or U5986 (N_5986,N_4391,N_3068);
nor U5987 (N_5987,N_4143,N_3167);
nand U5988 (N_5988,N_4467,N_3630);
and U5989 (N_5989,N_3280,N_3749);
and U5990 (N_5990,N_3821,N_3852);
or U5991 (N_5991,N_4359,N_3073);
nand U5992 (N_5992,N_4491,N_3064);
xnor U5993 (N_5993,N_3000,N_4201);
nor U5994 (N_5994,N_3086,N_3954);
and U5995 (N_5995,N_4219,N_4320);
or U5996 (N_5996,N_3634,N_3420);
nand U5997 (N_5997,N_3177,N_3018);
and U5998 (N_5998,N_4402,N_4091);
and U5999 (N_5999,N_4483,N_3219);
nand U6000 (N_6000,N_5763,N_5967);
and U6001 (N_6001,N_4676,N_5304);
or U6002 (N_6002,N_5698,N_4631);
xnor U6003 (N_6003,N_4638,N_5003);
nand U6004 (N_6004,N_5059,N_4980);
nor U6005 (N_6005,N_5801,N_4523);
or U6006 (N_6006,N_4788,N_4572);
or U6007 (N_6007,N_4987,N_4569);
nand U6008 (N_6008,N_5639,N_4560);
nor U6009 (N_6009,N_5173,N_4928);
or U6010 (N_6010,N_5308,N_5833);
nor U6011 (N_6011,N_4802,N_5566);
nor U6012 (N_6012,N_5167,N_5151);
xnor U6013 (N_6013,N_5751,N_5197);
xnor U6014 (N_6014,N_4862,N_5628);
nor U6015 (N_6015,N_4571,N_4827);
nor U6016 (N_6016,N_5079,N_5553);
or U6017 (N_6017,N_5839,N_5853);
and U6018 (N_6018,N_5903,N_5380);
or U6019 (N_6019,N_5448,N_5298);
nand U6020 (N_6020,N_5051,N_5679);
nor U6021 (N_6021,N_4771,N_5005);
nand U6022 (N_6022,N_5065,N_4597);
xor U6023 (N_6023,N_5602,N_4509);
and U6024 (N_6024,N_5860,N_5800);
nand U6025 (N_6025,N_5155,N_4901);
nand U6026 (N_6026,N_5940,N_4915);
nand U6027 (N_6027,N_4796,N_4990);
nor U6028 (N_6028,N_4511,N_5475);
and U6029 (N_6029,N_5507,N_4803);
and U6030 (N_6030,N_4902,N_4582);
and U6031 (N_6031,N_5343,N_4893);
nand U6032 (N_6032,N_5033,N_5152);
nand U6033 (N_6033,N_5489,N_5444);
xnor U6034 (N_6034,N_5458,N_5738);
xor U6035 (N_6035,N_5588,N_5206);
and U6036 (N_6036,N_4622,N_5867);
and U6037 (N_6037,N_5222,N_4800);
nand U6038 (N_6038,N_5815,N_5132);
nand U6039 (N_6039,N_4872,N_5876);
and U6040 (N_6040,N_5293,N_5412);
and U6041 (N_6041,N_4769,N_4508);
or U6042 (N_6042,N_5500,N_4999);
nor U6043 (N_6043,N_5965,N_5892);
or U6044 (N_6044,N_4846,N_5777);
nand U6045 (N_6045,N_4970,N_5520);
nand U6046 (N_6046,N_5269,N_5360);
or U6047 (N_6047,N_4659,N_5695);
nand U6048 (N_6048,N_5768,N_4557);
xnor U6049 (N_6049,N_4942,N_4691);
and U6050 (N_6050,N_4787,N_5970);
nor U6051 (N_6051,N_4592,N_5418);
or U6052 (N_6052,N_5002,N_5675);
nand U6053 (N_6053,N_4743,N_5527);
and U6054 (N_6054,N_5322,N_5341);
and U6055 (N_6055,N_5030,N_4965);
nand U6056 (N_6056,N_5519,N_5499);
nor U6057 (N_6057,N_5568,N_4640);
or U6058 (N_6058,N_4635,N_5376);
nand U6059 (N_6059,N_5202,N_4705);
xor U6060 (N_6060,N_5603,N_5462);
nor U6061 (N_6061,N_5313,N_5323);
nor U6062 (N_6062,N_4917,N_5516);
nor U6063 (N_6063,N_5439,N_5200);
nand U6064 (N_6064,N_5625,N_5311);
and U6065 (N_6065,N_5061,N_5897);
and U6066 (N_6066,N_5119,N_4782);
and U6067 (N_6067,N_5142,N_4945);
nor U6068 (N_6068,N_4543,N_5554);
nor U6069 (N_6069,N_5708,N_4766);
and U6070 (N_6070,N_5716,N_5433);
xor U6071 (N_6071,N_4794,N_5579);
and U6072 (N_6072,N_5630,N_5710);
xnor U6073 (N_6073,N_5348,N_4784);
nor U6074 (N_6074,N_4986,N_5547);
or U6075 (N_6075,N_5604,N_5232);
and U6076 (N_6076,N_4843,N_4645);
nor U6077 (N_6077,N_5596,N_5599);
nand U6078 (N_6078,N_5294,N_4927);
or U6079 (N_6079,N_5430,N_5368);
nand U6080 (N_6080,N_4727,N_4662);
and U6081 (N_6081,N_4867,N_5691);
nand U6082 (N_6082,N_5069,N_4922);
and U6083 (N_6083,N_4791,N_5153);
or U6084 (N_6084,N_4593,N_5822);
and U6085 (N_6085,N_4657,N_5624);
or U6086 (N_6086,N_5253,N_5001);
and U6087 (N_6087,N_5037,N_4778);
or U6088 (N_6088,N_5283,N_5621);
or U6089 (N_6089,N_5199,N_5943);
nand U6090 (N_6090,N_5674,N_5730);
and U6091 (N_6091,N_5884,N_4517);
or U6092 (N_6092,N_5830,N_5445);
or U6093 (N_6093,N_5807,N_5832);
nor U6094 (N_6094,N_5837,N_4684);
and U6095 (N_6095,N_5661,N_5670);
or U6096 (N_6096,N_5533,N_4751);
nor U6097 (N_6097,N_5141,N_5804);
nor U6098 (N_6098,N_5515,N_4541);
and U6099 (N_6099,N_5135,N_5618);
nor U6100 (N_6100,N_5175,N_4648);
or U6101 (N_6101,N_5045,N_5186);
xor U6102 (N_6102,N_4813,N_5361);
nor U6103 (N_6103,N_5413,N_4546);
nand U6104 (N_6104,N_5386,N_5461);
xnor U6105 (N_6105,N_4911,N_4905);
nor U6106 (N_6106,N_5310,N_5218);
xnor U6107 (N_6107,N_4768,N_5842);
nand U6108 (N_6108,N_5209,N_4786);
and U6109 (N_6109,N_5028,N_4644);
xnor U6110 (N_6110,N_4816,N_5177);
or U6111 (N_6111,N_4763,N_5834);
nor U6112 (N_6112,N_4741,N_5084);
and U6113 (N_6113,N_5782,N_5755);
nor U6114 (N_6114,N_5271,N_4797);
xor U6115 (N_6115,N_5983,N_5201);
nor U6116 (N_6116,N_5961,N_5287);
nand U6117 (N_6117,N_5063,N_5861);
or U6118 (N_6118,N_5565,N_4839);
nand U6119 (N_6119,N_5094,N_4701);
or U6120 (N_6120,N_5901,N_5594);
nor U6121 (N_6121,N_5849,N_4694);
or U6122 (N_6122,N_5728,N_5859);
nor U6123 (N_6123,N_4847,N_4716);
nand U6124 (N_6124,N_5948,N_5074);
nand U6125 (N_6125,N_4977,N_5297);
xor U6126 (N_6126,N_5761,N_5332);
and U6127 (N_6127,N_5279,N_5483);
and U6128 (N_6128,N_5052,N_5868);
xnor U6129 (N_6129,N_5981,N_5871);
xor U6130 (N_6130,N_5597,N_5355);
or U6131 (N_6131,N_4735,N_4721);
and U6132 (N_6132,N_5581,N_4835);
or U6133 (N_6133,N_5090,N_5934);
or U6134 (N_6134,N_5104,N_4682);
or U6135 (N_6135,N_5692,N_5466);
nor U6136 (N_6136,N_4711,N_4729);
or U6137 (N_6137,N_4836,N_5027);
nand U6138 (N_6138,N_5904,N_5543);
and U6139 (N_6139,N_5862,N_5518);
nand U6140 (N_6140,N_4929,N_5786);
and U6141 (N_6141,N_5685,N_5626);
and U6142 (N_6142,N_5473,N_4594);
or U6143 (N_6143,N_5858,N_5571);
and U6144 (N_6144,N_5098,N_5452);
and U6145 (N_6145,N_5771,N_4575);
and U6146 (N_6146,N_4725,N_5096);
xnor U6147 (N_6147,N_4527,N_4633);
or U6148 (N_6148,N_5337,N_5573);
or U6149 (N_6149,N_5422,N_5382);
nand U6150 (N_6150,N_4831,N_5406);
nand U6151 (N_6151,N_5133,N_4637);
nand U6152 (N_6152,N_4754,N_5787);
or U6153 (N_6153,N_4565,N_5798);
and U6154 (N_6154,N_4550,N_4742);
nand U6155 (N_6155,N_5923,N_4596);
or U6156 (N_6156,N_5657,N_5307);
and U6157 (N_6157,N_4628,N_4739);
and U6158 (N_6158,N_4530,N_5143);
nor U6159 (N_6159,N_5707,N_5012);
and U6160 (N_6160,N_5836,N_5379);
nor U6161 (N_6161,N_5536,N_5318);
nand U6162 (N_6162,N_5818,N_5600);
nor U6163 (N_6163,N_5668,N_4918);
nand U6164 (N_6164,N_4874,N_4608);
xor U6165 (N_6165,N_5211,N_4621);
nor U6166 (N_6166,N_5081,N_5844);
nor U6167 (N_6167,N_4762,N_4814);
nor U6168 (N_6168,N_4896,N_5053);
and U6169 (N_6169,N_5949,N_5721);
nand U6170 (N_6170,N_4781,N_5277);
or U6171 (N_6171,N_4719,N_4745);
nand U6172 (N_6172,N_5020,N_5673);
xor U6173 (N_6173,N_5963,N_5477);
nand U6174 (N_6174,N_4921,N_5369);
or U6175 (N_6175,N_5578,N_4825);
or U6176 (N_6176,N_4941,N_5300);
or U6177 (N_6177,N_4675,N_5916);
nor U6178 (N_6178,N_5829,N_5895);
or U6179 (N_6179,N_5956,N_4957);
or U6180 (N_6180,N_5817,N_5797);
nor U6181 (N_6181,N_5502,N_5306);
nor U6182 (N_6182,N_4618,N_5276);
nand U6183 (N_6183,N_5282,N_4907);
or U6184 (N_6184,N_5354,N_5016);
nor U6185 (N_6185,N_4764,N_5593);
or U6186 (N_6186,N_5711,N_5031);
nand U6187 (N_6187,N_5226,N_5749);
nor U6188 (N_6188,N_5678,N_4758);
nand U6189 (N_6189,N_4666,N_4604);
nor U6190 (N_6190,N_4544,N_5748);
xnor U6191 (N_6191,N_5291,N_5521);
nand U6192 (N_6192,N_5725,N_5776);
and U6193 (N_6193,N_5245,N_5442);
nor U6194 (N_6194,N_5023,N_5646);
and U6195 (N_6195,N_5150,N_4853);
or U6196 (N_6196,N_5178,N_5145);
nor U6197 (N_6197,N_5220,N_4536);
nand U6198 (N_6198,N_5945,N_5952);
and U6199 (N_6199,N_4677,N_5303);
or U6200 (N_6200,N_5043,N_4700);
xnor U6201 (N_6201,N_4547,N_5764);
xor U6202 (N_6202,N_4845,N_5899);
and U6203 (N_6203,N_5667,N_5498);
or U6204 (N_6204,N_5929,N_5056);
or U6205 (N_6205,N_5931,N_5476);
and U6206 (N_6206,N_4899,N_5078);
or U6207 (N_6207,N_5772,N_4548);
and U6208 (N_6208,N_5928,N_4903);
and U6209 (N_6209,N_5501,N_5780);
nor U6210 (N_6210,N_5456,N_4611);
nor U6211 (N_6211,N_5381,N_5932);
and U6212 (N_6212,N_5174,N_5130);
and U6213 (N_6213,N_5774,N_4649);
nand U6214 (N_6214,N_5877,N_5958);
nand U6215 (N_6215,N_5326,N_5508);
and U6216 (N_6216,N_4539,N_5008);
nor U6217 (N_6217,N_4968,N_4588);
xor U6218 (N_6218,N_5275,N_5947);
xnor U6219 (N_6219,N_5330,N_5658);
or U6220 (N_6220,N_5364,N_5273);
nand U6221 (N_6221,N_4605,N_4795);
nand U6222 (N_6222,N_4793,N_5762);
and U6223 (N_6223,N_5672,N_5723);
and U6224 (N_6224,N_5254,N_4576);
or U6225 (N_6225,N_5423,N_5257);
xnor U6226 (N_6226,N_4749,N_5587);
or U6227 (N_6227,N_4568,N_4889);
nor U6228 (N_6228,N_5816,N_4616);
nor U6229 (N_6229,N_5137,N_4856);
nor U6230 (N_6230,N_4993,N_4951);
or U6231 (N_6231,N_5560,N_5996);
nor U6232 (N_6232,N_4973,N_5214);
or U6233 (N_6233,N_5926,N_4686);
or U6234 (N_6234,N_4955,N_5927);
and U6235 (N_6235,N_5709,N_4943);
nor U6236 (N_6236,N_5154,N_4979);
nand U6237 (N_6237,N_5459,N_5266);
or U6238 (N_6238,N_5029,N_5985);
and U6239 (N_6239,N_5373,N_5595);
nand U6240 (N_6240,N_4533,N_4861);
and U6241 (N_6241,N_5921,N_5821);
nand U6242 (N_6242,N_5652,N_4776);
nor U6243 (N_6243,N_5605,N_5550);
nand U6244 (N_6244,N_4615,N_5457);
and U6245 (N_6245,N_5195,N_5083);
nand U6246 (N_6246,N_5555,N_5325);
xnor U6247 (N_6247,N_4809,N_4998);
xor U6248 (N_6248,N_4888,N_4953);
xor U6249 (N_6249,N_5460,N_5352);
nor U6250 (N_6250,N_5250,N_4949);
nor U6251 (N_6251,N_4702,N_5974);
nor U6252 (N_6252,N_5572,N_4878);
nor U6253 (N_6253,N_5158,N_4665);
nand U6254 (N_6254,N_5785,N_5885);
nor U6255 (N_6255,N_5471,N_5118);
or U6256 (N_6256,N_4906,N_5731);
nand U6257 (N_6257,N_5688,N_4822);
nand U6258 (N_6258,N_5788,N_5160);
or U6259 (N_6259,N_5169,N_5532);
nand U6260 (N_6260,N_5147,N_4969);
and U6261 (N_6261,N_5241,N_4512);
nand U6262 (N_6262,N_5035,N_4910);
or U6263 (N_6263,N_4894,N_4598);
xnor U6264 (N_6264,N_5700,N_5073);
nand U6265 (N_6265,N_5263,N_4866);
and U6266 (N_6266,N_5066,N_5334);
or U6267 (N_6267,N_5060,N_4963);
xor U6268 (N_6268,N_5993,N_5826);
and U6269 (N_6269,N_5845,N_5062);
nor U6270 (N_6270,N_5999,N_5436);
xnor U6271 (N_6271,N_5095,N_4559);
or U6272 (N_6272,N_4558,N_5126);
and U6273 (N_6273,N_4690,N_5631);
or U6274 (N_6274,N_4646,N_4890);
and U6275 (N_6275,N_5998,N_4678);
and U6276 (N_6276,N_4996,N_5684);
or U6277 (N_6277,N_4670,N_5643);
or U6278 (N_6278,N_5331,N_5907);
xnor U6279 (N_6279,N_5900,N_5584);
or U6280 (N_6280,N_5823,N_5429);
or U6281 (N_6281,N_5875,N_5942);
and U6282 (N_6282,N_5264,N_5258);
and U6283 (N_6283,N_4937,N_4715);
nand U6284 (N_6284,N_4868,N_5619);
nand U6285 (N_6285,N_5613,N_5997);
and U6286 (N_6286,N_5906,N_5280);
and U6287 (N_6287,N_5737,N_4783);
nand U6288 (N_6288,N_5038,N_5562);
xnor U6289 (N_6289,N_5611,N_5980);
nor U6290 (N_6290,N_5085,N_4962);
and U6291 (N_6291,N_5662,N_5064);
nand U6292 (N_6292,N_5159,N_4514);
or U6293 (N_6293,N_5795,N_5835);
or U6294 (N_6294,N_4760,N_5493);
nand U6295 (N_6295,N_4857,N_5262);
nor U6296 (N_6296,N_5274,N_4526);
xnor U6297 (N_6297,N_5359,N_5941);
and U6298 (N_6298,N_5704,N_4602);
and U6299 (N_6299,N_4551,N_5370);
nor U6300 (N_6300,N_5752,N_5401);
and U6301 (N_6301,N_4699,N_5874);
xnor U6302 (N_6302,N_4817,N_5347);
and U6303 (N_6303,N_4900,N_5960);
nand U6304 (N_6304,N_5358,N_5905);
and U6305 (N_6305,N_4829,N_4587);
or U6306 (N_6306,N_5210,N_4601);
nand U6307 (N_6307,N_4556,N_5015);
nand U6308 (N_6308,N_4661,N_4887);
and U6309 (N_6309,N_5641,N_5295);
xor U6310 (N_6310,N_4698,N_5225);
and U6311 (N_6311,N_5349,N_5841);
or U6312 (N_6312,N_5100,N_4688);
or U6313 (N_6313,N_5720,N_5191);
nor U6314 (N_6314,N_4734,N_5486);
or U6315 (N_6315,N_5338,N_5181);
or U6316 (N_6316,N_5248,N_5231);
nand U6317 (N_6317,N_4832,N_4767);
and U6318 (N_6318,N_4983,N_5117);
or U6319 (N_6319,N_4938,N_4780);
and U6320 (N_6320,N_5627,N_5070);
nor U6321 (N_6321,N_5350,N_4529);
xor U6322 (N_6322,N_5371,N_5789);
and U6323 (N_6323,N_4920,N_4561);
or U6324 (N_6324,N_5950,N_4830);
and U6325 (N_6325,N_4620,N_5729);
and U6326 (N_6326,N_4507,N_4750);
and U6327 (N_6327,N_4570,N_4641);
xor U6328 (N_6328,N_5478,N_5328);
nand U6329 (N_6329,N_5650,N_4926);
nand U6330 (N_6330,N_5067,N_5089);
or U6331 (N_6331,N_4583,N_5831);
or U6332 (N_6332,N_5959,N_4720);
xnor U6333 (N_6333,N_5592,N_5660);
and U6334 (N_6334,N_4824,N_4730);
and U6335 (N_6335,N_5116,N_5474);
nor U6336 (N_6336,N_5243,N_5055);
nand U6337 (N_6337,N_5425,N_4540);
nand U6338 (N_6338,N_5114,N_4685);
nand U6339 (N_6339,N_5221,N_5353);
nor U6340 (N_6340,N_5977,N_5395);
nor U6341 (N_6341,N_4988,N_4908);
nor U6342 (N_6342,N_4854,N_5865);
or U6343 (N_6343,N_5915,N_5889);
and U6344 (N_6344,N_5124,N_5071);
nor U6345 (N_6345,N_5170,N_5414);
xor U6346 (N_6346,N_5681,N_5086);
xnor U6347 (N_6347,N_5428,N_5744);
nand U6348 (N_6348,N_5718,N_5793);
nand U6349 (N_6349,N_5740,N_5006);
nor U6350 (N_6350,N_4756,N_4643);
and U6351 (N_6351,N_4673,N_5356);
or U6352 (N_6352,N_4870,N_5449);
or U6353 (N_6353,N_4947,N_4710);
nor U6354 (N_6354,N_5447,N_4834);
or U6355 (N_6355,N_4519,N_5470);
xnor U6356 (N_6356,N_5690,N_5107);
xor U6357 (N_6357,N_5261,N_5431);
nor U6358 (N_6358,N_4744,N_5256);
or U6359 (N_6359,N_5575,N_5995);
and U6360 (N_6360,N_5072,N_5882);
or U6361 (N_6361,N_5769,N_5446);
nand U6362 (N_6362,N_5405,N_5854);
nor U6363 (N_6363,N_4757,N_5714);
and U6364 (N_6364,N_5054,N_5409);
and U6365 (N_6365,N_5184,N_5205);
and U6366 (N_6366,N_5228,N_4554);
and U6367 (N_6367,N_5068,N_5548);
nor U6368 (N_6368,N_5391,N_5659);
nor U6369 (N_6369,N_4808,N_4833);
and U6370 (N_6370,N_5676,N_5187);
nor U6371 (N_6371,N_5601,N_4939);
nor U6372 (N_6372,N_5863,N_5286);
nor U6373 (N_6373,N_5962,N_5305);
nor U6374 (N_6374,N_5973,N_5230);
and U6375 (N_6375,N_5203,N_5252);
and U6376 (N_6376,N_5524,N_5810);
and U6377 (N_6377,N_4772,N_4599);
and U6378 (N_6378,N_4978,N_5635);
or U6379 (N_6379,N_4549,N_5978);
nand U6380 (N_6380,N_4703,N_5517);
nor U6381 (N_6381,N_5757,N_5157);
or U6382 (N_6382,N_4610,N_5563);
or U6383 (N_6383,N_5847,N_5649);
or U6384 (N_6384,N_5229,N_4828);
nor U6385 (N_6385,N_5827,N_5435);
xor U6386 (N_6386,N_5792,N_5050);
or U6387 (N_6387,N_4667,N_5247);
nand U6388 (N_6388,N_4934,N_4591);
and U6389 (N_6389,N_5496,N_4502);
nand U6390 (N_6390,N_5309,N_5136);
nand U6391 (N_6391,N_5781,N_5144);
or U6392 (N_6392,N_5267,N_5614);
nor U6393 (N_6393,N_5421,N_4818);
or U6394 (N_6394,N_5383,N_4707);
xor U6395 (N_6395,N_4736,N_5411);
nor U6396 (N_6396,N_5146,N_5869);
nor U6397 (N_6397,N_5735,N_4859);
nand U6398 (N_6398,N_5281,N_4562);
and U6399 (N_6399,N_4789,N_5042);
or U6400 (N_6400,N_5879,N_5481);
and U6401 (N_6401,N_4731,N_4737);
nand U6402 (N_6402,N_4869,N_5416);
nand U6403 (N_6403,N_5522,N_5290);
or U6404 (N_6404,N_4580,N_5864);
nand U6405 (N_6405,N_4848,N_4566);
or U6406 (N_6406,N_5622,N_5213);
or U6407 (N_6407,N_4586,N_4932);
and U6408 (N_6408,N_5128,N_5758);
nand U6409 (N_6409,N_4724,N_5888);
nand U6410 (N_6410,N_4679,N_5558);
nor U6411 (N_6411,N_5388,N_5122);
xor U6412 (N_6412,N_5873,N_5883);
nand U6413 (N_6413,N_4520,N_4653);
and U6414 (N_6414,N_4722,N_4807);
and U6415 (N_6415,N_4801,N_5149);
or U6416 (N_6416,N_5389,N_5312);
nor U6417 (N_6417,N_4681,N_4634);
nor U6418 (N_6418,N_5492,N_4972);
or U6419 (N_6419,N_5467,N_5936);
and U6420 (N_6420,N_4753,N_4775);
nand U6421 (N_6421,N_4812,N_5426);
nor U6422 (N_6422,N_4627,N_5766);
and U6423 (N_6423,N_4785,N_5022);
xor U6424 (N_6424,N_5753,N_4858);
or U6425 (N_6425,N_5301,N_4819);
nor U6426 (N_6426,N_4642,N_5687);
and U6427 (N_6427,N_5537,N_5384);
nand U6428 (N_6428,N_5469,N_5011);
or U6429 (N_6429,N_5724,N_5227);
or U6430 (N_6430,N_5574,N_5912);
or U6431 (N_6431,N_5494,N_4689);
or U6432 (N_6432,N_5443,N_4933);
nand U6433 (N_6433,N_5234,N_4579);
and U6434 (N_6434,N_4585,N_4823);
nor U6435 (N_6435,N_5398,N_5196);
nand U6436 (N_6436,N_5607,N_4936);
or U6437 (N_6437,N_4733,N_5803);
or U6438 (N_6438,N_4991,N_5726);
and U6439 (N_6439,N_5866,N_5420);
and U6440 (N_6440,N_5819,N_4738);
and U6441 (N_6441,N_5924,N_5212);
and U6442 (N_6442,N_5825,N_4884);
and U6443 (N_6443,N_5026,N_4518);
or U6444 (N_6444,N_5327,N_4864);
or U6445 (N_6445,N_5397,N_5561);
nand U6446 (N_6446,N_5288,N_4697);
and U6447 (N_6447,N_4948,N_5182);
nand U6448 (N_6448,N_5925,N_5390);
or U6449 (N_6449,N_5168,N_4909);
nor U6450 (N_6450,N_5018,N_5972);
and U6451 (N_6451,N_5034,N_5633);
or U6452 (N_6452,N_5259,N_5106);
nor U6453 (N_6453,N_5556,N_5669);
xor U6454 (N_6454,N_4704,N_5392);
or U6455 (N_6455,N_4882,N_5189);
and U6456 (N_6456,N_4981,N_5138);
and U6457 (N_6457,N_5653,N_5655);
nand U6458 (N_6458,N_4984,N_5260);
nor U6459 (N_6459,N_5609,N_5108);
or U6460 (N_6460,N_4912,N_5166);
and U6461 (N_6461,N_5564,N_4654);
xnor U6462 (N_6462,N_5233,N_4687);
and U6463 (N_6463,N_5796,N_5506);
nand U6464 (N_6464,N_4871,N_5249);
or U6465 (N_6465,N_5497,N_4924);
or U6466 (N_6466,N_4625,N_5680);
and U6467 (N_6467,N_4564,N_5616);
nor U6468 (N_6468,N_5188,N_5741);
or U6469 (N_6469,N_5677,N_5238);
nand U6470 (N_6470,N_5994,N_4728);
nand U6471 (N_6471,N_5165,N_4895);
and U6472 (N_6472,N_5407,N_4614);
or U6473 (N_6473,N_5617,N_5989);
nand U6474 (N_6474,N_5346,N_4537);
nor U6475 (N_6475,N_4726,N_4804);
or U6476 (N_6476,N_5846,N_5468);
and U6477 (N_6477,N_5415,N_5246);
nand U6478 (N_6478,N_5190,N_5434);
nor U6479 (N_6479,N_5036,N_5127);
or U6480 (N_6480,N_5747,N_5756);
xnor U6481 (N_6481,N_5185,N_5419);
and U6482 (N_6482,N_4723,N_5482);
nand U6483 (N_6483,N_4680,N_5966);
nand U6484 (N_6484,N_5240,N_5585);
nand U6485 (N_6485,N_5284,N_4574);
and U6486 (N_6486,N_4841,N_5180);
nand U6487 (N_6487,N_5582,N_5664);
nor U6488 (N_6488,N_4779,N_5530);
xor U6489 (N_6489,N_5134,N_5316);
and U6490 (N_6490,N_5779,N_5441);
and U6491 (N_6491,N_5850,N_5340);
or U6492 (N_6492,N_5239,N_4950);
or U6493 (N_6493,N_5976,N_4747);
and U6494 (N_6494,N_5911,N_5285);
nor U6495 (N_6495,N_5544,N_5784);
or U6496 (N_6496,N_5387,N_5080);
nor U6497 (N_6497,N_4664,N_5656);
and U6498 (N_6498,N_5612,N_5296);
and U6499 (N_6499,N_5852,N_5606);
and U6500 (N_6500,N_4590,N_4504);
or U6501 (N_6501,N_4852,N_5366);
nor U6502 (N_6502,N_4531,N_5615);
xnor U6503 (N_6503,N_4595,N_4521);
xor U6504 (N_6504,N_5463,N_5374);
nand U6505 (N_6505,N_5894,N_5986);
or U6506 (N_6506,N_5265,N_5552);
or U6507 (N_6507,N_5908,N_5717);
xor U6508 (N_6508,N_4844,N_4515);
nor U6509 (N_6509,N_5317,N_5534);
and U6510 (N_6510,N_5523,N_5887);
and U6511 (N_6511,N_5372,N_4904);
nand U6512 (N_6512,N_5339,N_5870);
nand U6513 (N_6513,N_5820,N_5909);
nand U6514 (N_6514,N_4600,N_5007);
nor U6515 (N_6515,N_4660,N_5828);
nor U6516 (N_6516,N_5629,N_5465);
and U6517 (N_6517,N_5025,N_5964);
nor U6518 (N_6518,N_5968,N_4522);
and U6519 (N_6519,N_5598,N_5734);
nand U6520 (N_6520,N_5451,N_5333);
and U6521 (N_6521,N_5770,N_4994);
nor U6522 (N_6522,N_5937,N_5076);
nand U6523 (N_6523,N_5855,N_5988);
and U6524 (N_6524,N_5946,N_5851);
nor U6525 (N_6525,N_5693,N_4880);
or U6526 (N_6526,N_4506,N_4940);
nand U6527 (N_6527,N_4573,N_5215);
or U6528 (N_6528,N_5363,N_5933);
xnor U6529 (N_6529,N_5378,N_4877);
nand U6530 (N_6530,N_5099,N_5408);
nor U6531 (N_6531,N_5299,N_5204);
xnor U6532 (N_6532,N_4958,N_5048);
nor U6533 (N_6533,N_4706,N_5019);
or U6534 (N_6534,N_5918,N_4647);
nor U6535 (N_6535,N_5583,N_4840);
nor U6536 (N_6536,N_5024,N_5512);
nor U6537 (N_6537,N_4913,N_5739);
and U6538 (N_6538,N_5857,N_4919);
nor U6539 (N_6539,N_5638,N_5697);
or U6540 (N_6540,N_5944,N_4525);
xor U6541 (N_6541,N_5917,N_4790);
xnor U6542 (N_6542,N_5375,N_4740);
and U6543 (N_6543,N_4708,N_4589);
nor U6544 (N_6544,N_5955,N_5041);
or U6545 (N_6545,N_5637,N_5345);
nor U6546 (N_6546,N_4626,N_5087);
or U6547 (N_6547,N_5896,N_4837);
xor U6548 (N_6548,N_5694,N_4851);
nand U6549 (N_6549,N_5910,N_4607);
nand U6550 (N_6550,N_4876,N_4553);
nor U6551 (N_6551,N_4538,N_5654);
or U6552 (N_6552,N_5393,N_4606);
or U6553 (N_6553,N_5808,N_5632);
or U6554 (N_6554,N_5647,N_5577);
xnor U6555 (N_6555,N_5013,N_5957);
nor U6556 (N_6556,N_5791,N_5236);
and U6557 (N_6557,N_5886,N_4931);
and U6558 (N_6558,N_5403,N_5163);
or U6559 (N_6559,N_5890,N_5112);
or U6560 (N_6560,N_4759,N_4952);
nand U6561 (N_6561,N_4985,N_4632);
nand U6562 (N_6562,N_5775,N_5715);
and U6563 (N_6563,N_5148,N_5365);
nand U6564 (N_6564,N_5032,N_4891);
nand U6565 (N_6565,N_5545,N_5251);
nor U6566 (N_6566,N_5809,N_4528);
nor U6567 (N_6567,N_5156,N_5759);
xnor U6568 (N_6568,N_5139,N_5125);
xor U6569 (N_6569,N_5039,N_5878);
and U6570 (N_6570,N_5289,N_5951);
nand U6571 (N_6571,N_5671,N_5838);
nand U6572 (N_6572,N_5495,N_5546);
or U6573 (N_6573,N_5736,N_5472);
and U6574 (N_6574,N_5417,N_4672);
nand U6575 (N_6575,N_4752,N_4693);
and U6576 (N_6576,N_5046,N_5292);
nor U6577 (N_6577,N_5696,N_5400);
or U6578 (N_6578,N_5712,N_4656);
or U6579 (N_6579,N_5705,N_4805);
nor U6580 (N_6580,N_4695,N_4923);
and U6581 (N_6581,N_5319,N_4992);
or U6582 (N_6582,N_4567,N_5610);
nand U6583 (N_6583,N_4658,N_5329);
nor U6584 (N_6584,N_4886,N_5802);
nand U6585 (N_6585,N_4503,N_4714);
nor U6586 (N_6586,N_5713,N_5984);
nor U6587 (N_6587,N_5531,N_4946);
or U6588 (N_6588,N_4624,N_4885);
nor U6589 (N_6589,N_5424,N_4930);
nand U6590 (N_6590,N_5235,N_5767);
nand U6591 (N_6591,N_5314,N_5953);
and U6592 (N_6592,N_4961,N_4944);
and U6593 (N_6593,N_5490,N_5902);
or U6594 (N_6594,N_5919,N_5743);
and U6595 (N_6595,N_4956,N_5569);
nand U6596 (N_6596,N_4532,N_5432);
xnor U6597 (N_6597,N_5485,N_5224);
and U6598 (N_6598,N_5898,N_4732);
xnor U6599 (N_6599,N_5453,N_5848);
nor U6600 (N_6600,N_4954,N_5636);
and U6601 (N_6601,N_4577,N_5437);
and U6602 (N_6602,N_5320,N_4774);
or U6603 (N_6603,N_5105,N_4668);
or U6604 (N_6604,N_5014,N_5193);
and U6605 (N_6605,N_4964,N_4612);
nand U6606 (N_6606,N_5454,N_5856);
or U6607 (N_6607,N_4630,N_5207);
and U6608 (N_6608,N_5754,N_5047);
nand U6609 (N_6609,N_5806,N_5487);
nand U6610 (N_6610,N_4623,N_5402);
xor U6611 (N_6611,N_5514,N_5396);
nor U6612 (N_6612,N_4770,N_5399);
xnor U6613 (N_6613,N_4935,N_5101);
nand U6614 (N_6614,N_4975,N_5760);
or U6615 (N_6615,N_5140,N_5255);
and U6616 (N_6616,N_5336,N_4545);
nand U6617 (N_6617,N_4842,N_4516);
or U6618 (N_6618,N_5733,N_5131);
and U6619 (N_6619,N_5161,N_5703);
nand U6620 (N_6620,N_5666,N_5969);
or U6621 (N_6621,N_5686,N_5103);
xnor U6622 (N_6622,N_5732,N_5044);
nand U6623 (N_6623,N_4892,N_4603);
nor U6624 (N_6624,N_5077,N_5367);
xor U6625 (N_6625,N_5750,N_5479);
nand U6626 (N_6626,N_4960,N_4976);
nand U6627 (N_6627,N_5746,N_5183);
nor U6628 (N_6628,N_5324,N_4692);
or U6629 (N_6629,N_4717,N_5745);
and U6630 (N_6630,N_4820,N_5427);
nand U6631 (N_6631,N_5542,N_5216);
nor U6632 (N_6632,N_5362,N_4925);
nand U6633 (N_6633,N_5377,N_5129);
or U6634 (N_6634,N_5491,N_5171);
or U6635 (N_6635,N_5110,N_5794);
nor U6636 (N_6636,N_5773,N_5464);
and U6637 (N_6637,N_4683,N_4578);
or U6638 (N_6638,N_4709,N_4655);
or U6639 (N_6639,N_5765,N_4959);
xnor U6640 (N_6640,N_5088,N_5509);
nor U6641 (N_6641,N_5891,N_5778);
xor U6642 (N_6642,N_5805,N_5164);
and U6643 (N_6643,N_5410,N_4815);
nand U6644 (N_6644,N_5590,N_4513);
nand U6645 (N_6645,N_5505,N_5799);
and U6646 (N_6646,N_5930,N_4617);
and U6647 (N_6647,N_4806,N_5811);
xor U6648 (N_6648,N_5455,N_5082);
or U6649 (N_6649,N_5814,N_5321);
xor U6650 (N_6650,N_5484,N_5513);
and U6651 (N_6651,N_5576,N_5840);
nor U6652 (N_6652,N_5651,N_5990);
nor U6653 (N_6653,N_5529,N_5111);
nand U6654 (N_6654,N_4652,N_5722);
and U6655 (N_6655,N_4897,N_5872);
or U6656 (N_6656,N_4639,N_5109);
nand U6657 (N_6657,N_4581,N_5608);
or U6658 (N_6658,N_4777,N_4997);
nor U6659 (N_6659,N_4712,N_5992);
nor U6660 (N_6660,N_5057,N_5438);
and U6661 (N_6661,N_4792,N_4881);
and U6662 (N_6662,N_5115,N_5683);
nor U6663 (N_6663,N_5935,N_5640);
xnor U6664 (N_6664,N_5557,N_4883);
and U6665 (N_6665,N_4860,N_5979);
and U6666 (N_6666,N_5278,N_5812);
nand U6667 (N_6667,N_4838,N_5701);
nor U6668 (N_6668,N_5634,N_5162);
nand U6669 (N_6669,N_5342,N_5268);
nor U6670 (N_6670,N_5938,N_5010);
and U6671 (N_6671,N_5075,N_4995);
or U6672 (N_6672,N_5121,N_5102);
or U6673 (N_6673,N_5824,N_5893);
nand U6674 (N_6674,N_5315,N_4609);
nor U6675 (N_6675,N_5488,N_5480);
nor U6676 (N_6676,N_5120,N_4748);
nand U6677 (N_6677,N_4865,N_5682);
or U6678 (N_6678,N_5541,N_5913);
or U6679 (N_6679,N_4773,N_5058);
nor U6680 (N_6680,N_5237,N_4916);
nand U6681 (N_6681,N_5539,N_5702);
or U6682 (N_6682,N_5727,N_4798);
nand U6683 (N_6683,N_4799,N_5663);
nor U6684 (N_6684,N_5176,N_5567);
nand U6685 (N_6685,N_4713,N_5244);
xor U6686 (N_6686,N_4761,N_5219);
or U6687 (N_6687,N_5549,N_4524);
or U6688 (N_6688,N_4636,N_5385);
xnor U6689 (N_6689,N_4534,N_5991);
nand U6690 (N_6690,N_5242,N_5922);
or U6691 (N_6691,N_5987,N_5302);
xnor U6692 (N_6692,N_4879,N_5049);
xnor U6693 (N_6693,N_4875,N_5881);
nor U6694 (N_6694,N_5017,N_4619);
nand U6695 (N_6695,N_4914,N_4849);
or U6696 (N_6696,N_4718,N_5689);
nor U6697 (N_6697,N_5351,N_5645);
and U6698 (N_6698,N_4555,N_4826);
and U6699 (N_6699,N_5009,N_4535);
and U6700 (N_6700,N_5503,N_5644);
nor U6701 (N_6701,N_5440,N_4584);
nand U6702 (N_6702,N_5208,N_5172);
nand U6703 (N_6703,N_5344,N_4669);
xor U6704 (N_6704,N_5004,N_5192);
nor U6705 (N_6705,N_5021,N_5123);
and U6706 (N_6706,N_4811,N_4873);
xnor U6707 (N_6707,N_5699,N_5843);
and U6708 (N_6708,N_5113,N_4650);
nor U6709 (N_6709,N_5620,N_4974);
and U6710 (N_6710,N_5357,N_4971);
nor U6711 (N_6711,N_5813,N_5528);
xor U6712 (N_6712,N_4629,N_5270);
nor U6713 (N_6713,N_5591,N_5975);
and U6714 (N_6714,N_4663,N_5880);
nand U6715 (N_6715,N_4651,N_5217);
nand U6716 (N_6716,N_5510,N_5538);
and U6717 (N_6717,N_5706,N_5790);
and U6718 (N_6718,N_5093,N_5097);
nor U6719 (N_6719,N_5540,N_5920);
nor U6720 (N_6720,N_5580,N_5194);
or U6721 (N_6721,N_5450,N_4855);
nand U6722 (N_6722,N_5198,N_5394);
nand U6723 (N_6723,N_4671,N_4810);
nor U6724 (N_6724,N_5525,N_5642);
nand U6725 (N_6725,N_5742,N_5648);
nand U6726 (N_6726,N_5223,N_5589);
and U6727 (N_6727,N_4500,N_4967);
nor U6728 (N_6728,N_4505,N_5551);
nor U6729 (N_6729,N_4898,N_5000);
or U6730 (N_6730,N_4510,N_5526);
nand U6731 (N_6731,N_4982,N_5665);
nor U6732 (N_6732,N_5783,N_5272);
and U6733 (N_6733,N_5040,N_4765);
or U6734 (N_6734,N_5511,N_5179);
nor U6735 (N_6735,N_5535,N_5623);
nor U6736 (N_6736,N_4746,N_4542);
and U6737 (N_6737,N_5504,N_4863);
or U6738 (N_6738,N_5335,N_5092);
nand U6739 (N_6739,N_4989,N_4563);
nand U6740 (N_6740,N_4552,N_5559);
nand U6741 (N_6741,N_5954,N_4755);
and U6742 (N_6742,N_4613,N_5570);
nand U6743 (N_6743,N_4821,N_4674);
nand U6744 (N_6744,N_5091,N_5404);
or U6745 (N_6745,N_5982,N_5914);
nand U6746 (N_6746,N_4696,N_5719);
nor U6747 (N_6747,N_5939,N_5586);
nor U6748 (N_6748,N_4850,N_4966);
xnor U6749 (N_6749,N_4501,N_5971);
and U6750 (N_6750,N_5532,N_5044);
xnor U6751 (N_6751,N_4624,N_4892);
nand U6752 (N_6752,N_5882,N_5279);
and U6753 (N_6753,N_5082,N_4633);
and U6754 (N_6754,N_5187,N_4928);
and U6755 (N_6755,N_4546,N_4813);
nand U6756 (N_6756,N_5195,N_5645);
nor U6757 (N_6757,N_4732,N_5967);
or U6758 (N_6758,N_5840,N_4610);
and U6759 (N_6759,N_5298,N_5806);
nand U6760 (N_6760,N_4969,N_5809);
nand U6761 (N_6761,N_5015,N_4754);
and U6762 (N_6762,N_5839,N_5796);
nor U6763 (N_6763,N_5429,N_5476);
or U6764 (N_6764,N_4638,N_4707);
nor U6765 (N_6765,N_4784,N_4726);
and U6766 (N_6766,N_4501,N_5094);
and U6767 (N_6767,N_5932,N_4647);
or U6768 (N_6768,N_4605,N_5199);
and U6769 (N_6769,N_5993,N_5157);
nor U6770 (N_6770,N_4592,N_5327);
nor U6771 (N_6771,N_5173,N_4529);
and U6772 (N_6772,N_5484,N_4812);
nand U6773 (N_6773,N_5684,N_5247);
and U6774 (N_6774,N_4897,N_5543);
or U6775 (N_6775,N_5231,N_5677);
nand U6776 (N_6776,N_5334,N_5597);
and U6777 (N_6777,N_5562,N_5906);
nor U6778 (N_6778,N_5740,N_5870);
nor U6779 (N_6779,N_5473,N_5253);
nor U6780 (N_6780,N_5329,N_5705);
nand U6781 (N_6781,N_5330,N_4883);
and U6782 (N_6782,N_5730,N_5948);
nor U6783 (N_6783,N_5148,N_4975);
or U6784 (N_6784,N_5767,N_5748);
and U6785 (N_6785,N_5753,N_4550);
or U6786 (N_6786,N_5356,N_5474);
and U6787 (N_6787,N_5140,N_5597);
nand U6788 (N_6788,N_5397,N_5904);
nor U6789 (N_6789,N_5525,N_5038);
nand U6790 (N_6790,N_5239,N_5991);
nor U6791 (N_6791,N_5597,N_4905);
or U6792 (N_6792,N_5070,N_5587);
or U6793 (N_6793,N_5512,N_5808);
and U6794 (N_6794,N_5150,N_4747);
and U6795 (N_6795,N_5613,N_4959);
xnor U6796 (N_6796,N_4508,N_5789);
and U6797 (N_6797,N_4875,N_4791);
nor U6798 (N_6798,N_5238,N_5920);
xnor U6799 (N_6799,N_4796,N_4886);
or U6800 (N_6800,N_4561,N_5575);
nand U6801 (N_6801,N_4638,N_5962);
xnor U6802 (N_6802,N_4623,N_5105);
and U6803 (N_6803,N_5954,N_4818);
nor U6804 (N_6804,N_5124,N_4862);
nand U6805 (N_6805,N_5709,N_4996);
xor U6806 (N_6806,N_5330,N_5471);
nand U6807 (N_6807,N_5932,N_5711);
nor U6808 (N_6808,N_4913,N_5524);
or U6809 (N_6809,N_5666,N_5726);
nand U6810 (N_6810,N_5758,N_5870);
nor U6811 (N_6811,N_4725,N_4672);
xor U6812 (N_6812,N_4741,N_4621);
or U6813 (N_6813,N_4733,N_5146);
nand U6814 (N_6814,N_4895,N_5115);
nand U6815 (N_6815,N_5078,N_5109);
nor U6816 (N_6816,N_5120,N_4679);
nor U6817 (N_6817,N_4948,N_4570);
and U6818 (N_6818,N_5958,N_5085);
nor U6819 (N_6819,N_5537,N_5318);
and U6820 (N_6820,N_5254,N_4897);
or U6821 (N_6821,N_5958,N_4786);
nand U6822 (N_6822,N_5435,N_4809);
nor U6823 (N_6823,N_5747,N_4859);
nand U6824 (N_6824,N_5758,N_5643);
and U6825 (N_6825,N_5269,N_4744);
nor U6826 (N_6826,N_4657,N_5352);
nand U6827 (N_6827,N_5101,N_5163);
and U6828 (N_6828,N_5134,N_5861);
nor U6829 (N_6829,N_4747,N_5454);
or U6830 (N_6830,N_5447,N_5445);
nand U6831 (N_6831,N_5237,N_5213);
and U6832 (N_6832,N_5198,N_4969);
nand U6833 (N_6833,N_4516,N_5580);
nand U6834 (N_6834,N_4623,N_5959);
xor U6835 (N_6835,N_5925,N_5127);
xnor U6836 (N_6836,N_4529,N_5139);
nand U6837 (N_6837,N_5084,N_5416);
nor U6838 (N_6838,N_5955,N_5242);
nand U6839 (N_6839,N_5837,N_4613);
or U6840 (N_6840,N_5236,N_5669);
nand U6841 (N_6841,N_4920,N_5607);
nor U6842 (N_6842,N_5697,N_5257);
nand U6843 (N_6843,N_4550,N_4674);
nor U6844 (N_6844,N_5356,N_4548);
and U6845 (N_6845,N_4741,N_4577);
nor U6846 (N_6846,N_5943,N_5523);
nor U6847 (N_6847,N_5495,N_4923);
or U6848 (N_6848,N_4998,N_5646);
nor U6849 (N_6849,N_5964,N_5324);
and U6850 (N_6850,N_5238,N_4899);
or U6851 (N_6851,N_5189,N_5377);
and U6852 (N_6852,N_4978,N_4976);
and U6853 (N_6853,N_5011,N_4812);
or U6854 (N_6854,N_5973,N_5368);
and U6855 (N_6855,N_5390,N_4561);
or U6856 (N_6856,N_5777,N_5354);
or U6857 (N_6857,N_5982,N_5559);
nor U6858 (N_6858,N_5621,N_5851);
or U6859 (N_6859,N_4766,N_5329);
or U6860 (N_6860,N_4787,N_5962);
and U6861 (N_6861,N_5103,N_5934);
and U6862 (N_6862,N_5311,N_5937);
or U6863 (N_6863,N_4735,N_5903);
nor U6864 (N_6864,N_5774,N_4622);
or U6865 (N_6865,N_5691,N_5234);
and U6866 (N_6866,N_5653,N_5976);
and U6867 (N_6867,N_5514,N_5411);
nor U6868 (N_6868,N_5865,N_5649);
nor U6869 (N_6869,N_4503,N_4988);
nor U6870 (N_6870,N_5215,N_4841);
nand U6871 (N_6871,N_5891,N_5915);
or U6872 (N_6872,N_4682,N_5211);
nor U6873 (N_6873,N_5092,N_5190);
xnor U6874 (N_6874,N_5485,N_4748);
and U6875 (N_6875,N_5394,N_5546);
nand U6876 (N_6876,N_5246,N_5493);
and U6877 (N_6877,N_5075,N_5977);
and U6878 (N_6878,N_5151,N_5572);
or U6879 (N_6879,N_4549,N_5544);
or U6880 (N_6880,N_5304,N_5860);
nand U6881 (N_6881,N_4544,N_5622);
or U6882 (N_6882,N_4672,N_5639);
nor U6883 (N_6883,N_5476,N_5529);
nor U6884 (N_6884,N_4677,N_5496);
xnor U6885 (N_6885,N_5233,N_5249);
or U6886 (N_6886,N_5053,N_5122);
nand U6887 (N_6887,N_5544,N_5812);
nor U6888 (N_6888,N_5865,N_4650);
and U6889 (N_6889,N_5203,N_5668);
nand U6890 (N_6890,N_4911,N_4949);
nand U6891 (N_6891,N_4851,N_4911);
xor U6892 (N_6892,N_5917,N_4958);
nand U6893 (N_6893,N_5377,N_5572);
or U6894 (N_6894,N_5216,N_5785);
xor U6895 (N_6895,N_5886,N_5490);
xnor U6896 (N_6896,N_5476,N_5716);
and U6897 (N_6897,N_5509,N_5460);
and U6898 (N_6898,N_5128,N_5896);
or U6899 (N_6899,N_5930,N_5437);
nor U6900 (N_6900,N_4864,N_5801);
nand U6901 (N_6901,N_5800,N_4716);
and U6902 (N_6902,N_5909,N_5142);
nand U6903 (N_6903,N_4592,N_5140);
and U6904 (N_6904,N_4631,N_5584);
nor U6905 (N_6905,N_5940,N_4865);
and U6906 (N_6906,N_5984,N_4993);
or U6907 (N_6907,N_5808,N_4925);
or U6908 (N_6908,N_4960,N_5068);
nor U6909 (N_6909,N_4637,N_4808);
nor U6910 (N_6910,N_5635,N_5595);
and U6911 (N_6911,N_5541,N_5786);
and U6912 (N_6912,N_5227,N_4889);
or U6913 (N_6913,N_4854,N_4975);
nor U6914 (N_6914,N_5121,N_5009);
nand U6915 (N_6915,N_4750,N_4607);
and U6916 (N_6916,N_5620,N_5872);
nor U6917 (N_6917,N_5650,N_4974);
or U6918 (N_6918,N_4898,N_5724);
or U6919 (N_6919,N_4654,N_5696);
xor U6920 (N_6920,N_5177,N_4664);
nor U6921 (N_6921,N_5630,N_5616);
nor U6922 (N_6922,N_5748,N_4825);
or U6923 (N_6923,N_5654,N_5780);
nor U6924 (N_6924,N_4729,N_4887);
or U6925 (N_6925,N_4679,N_4526);
xor U6926 (N_6926,N_5803,N_4761);
and U6927 (N_6927,N_5854,N_5092);
nor U6928 (N_6928,N_4534,N_5195);
nand U6929 (N_6929,N_5622,N_5379);
xnor U6930 (N_6930,N_5484,N_5755);
nor U6931 (N_6931,N_5501,N_5971);
or U6932 (N_6932,N_5647,N_4976);
nor U6933 (N_6933,N_5922,N_5836);
or U6934 (N_6934,N_5888,N_4762);
nand U6935 (N_6935,N_5870,N_4544);
nand U6936 (N_6936,N_5432,N_4613);
nand U6937 (N_6937,N_4719,N_4611);
or U6938 (N_6938,N_4771,N_4567);
and U6939 (N_6939,N_5844,N_5479);
nand U6940 (N_6940,N_5642,N_4646);
xor U6941 (N_6941,N_4882,N_5319);
and U6942 (N_6942,N_4946,N_5334);
and U6943 (N_6943,N_5151,N_5040);
xor U6944 (N_6944,N_4860,N_5711);
and U6945 (N_6945,N_4796,N_5471);
or U6946 (N_6946,N_4607,N_5874);
nand U6947 (N_6947,N_4500,N_5816);
and U6948 (N_6948,N_4821,N_4862);
nor U6949 (N_6949,N_5508,N_5374);
and U6950 (N_6950,N_5028,N_5765);
xor U6951 (N_6951,N_4883,N_4870);
nand U6952 (N_6952,N_4883,N_5181);
nor U6953 (N_6953,N_5862,N_5767);
nand U6954 (N_6954,N_4525,N_4500);
nand U6955 (N_6955,N_4694,N_4978);
nand U6956 (N_6956,N_5593,N_4911);
nand U6957 (N_6957,N_5864,N_5133);
nand U6958 (N_6958,N_5754,N_4684);
or U6959 (N_6959,N_4869,N_5972);
or U6960 (N_6960,N_5979,N_5364);
and U6961 (N_6961,N_5547,N_5261);
or U6962 (N_6962,N_5533,N_4725);
nor U6963 (N_6963,N_5554,N_5476);
nor U6964 (N_6964,N_5842,N_5214);
nand U6965 (N_6965,N_5111,N_5558);
or U6966 (N_6966,N_5944,N_5063);
nor U6967 (N_6967,N_5064,N_4584);
or U6968 (N_6968,N_5907,N_4867);
or U6969 (N_6969,N_4975,N_5772);
or U6970 (N_6970,N_5666,N_4928);
nand U6971 (N_6971,N_4578,N_4697);
nor U6972 (N_6972,N_5021,N_5871);
or U6973 (N_6973,N_5923,N_5733);
or U6974 (N_6974,N_5364,N_5405);
and U6975 (N_6975,N_4805,N_5737);
nor U6976 (N_6976,N_4974,N_5474);
nand U6977 (N_6977,N_5744,N_5857);
xnor U6978 (N_6978,N_5353,N_5807);
nand U6979 (N_6979,N_5503,N_5468);
or U6980 (N_6980,N_4820,N_5057);
or U6981 (N_6981,N_5578,N_5773);
xnor U6982 (N_6982,N_5300,N_5209);
nand U6983 (N_6983,N_4966,N_5810);
or U6984 (N_6984,N_4988,N_5803);
and U6985 (N_6985,N_5521,N_4934);
or U6986 (N_6986,N_4705,N_5815);
xor U6987 (N_6987,N_4683,N_5941);
and U6988 (N_6988,N_4979,N_5397);
and U6989 (N_6989,N_5014,N_4983);
nor U6990 (N_6990,N_5232,N_5855);
and U6991 (N_6991,N_5935,N_4996);
nand U6992 (N_6992,N_4856,N_5839);
nor U6993 (N_6993,N_5727,N_4966);
and U6994 (N_6994,N_5261,N_5862);
and U6995 (N_6995,N_5319,N_5429);
and U6996 (N_6996,N_5977,N_4500);
or U6997 (N_6997,N_5219,N_4636);
nand U6998 (N_6998,N_4551,N_5123);
xor U6999 (N_6999,N_5916,N_5593);
and U7000 (N_7000,N_5235,N_4925);
or U7001 (N_7001,N_5075,N_4716);
and U7002 (N_7002,N_5484,N_5815);
nand U7003 (N_7003,N_5313,N_5610);
nand U7004 (N_7004,N_4939,N_5342);
and U7005 (N_7005,N_4674,N_5184);
and U7006 (N_7006,N_5039,N_5445);
or U7007 (N_7007,N_4659,N_4639);
nor U7008 (N_7008,N_5501,N_5918);
nand U7009 (N_7009,N_5271,N_4974);
or U7010 (N_7010,N_5347,N_5733);
or U7011 (N_7011,N_5979,N_4672);
nor U7012 (N_7012,N_5881,N_5972);
nand U7013 (N_7013,N_5364,N_5599);
or U7014 (N_7014,N_4982,N_5290);
nand U7015 (N_7015,N_4768,N_5093);
nor U7016 (N_7016,N_5594,N_4595);
or U7017 (N_7017,N_4742,N_5830);
nand U7018 (N_7018,N_4924,N_4869);
xor U7019 (N_7019,N_5753,N_4556);
nand U7020 (N_7020,N_5658,N_4616);
or U7021 (N_7021,N_5222,N_4771);
and U7022 (N_7022,N_4907,N_5352);
and U7023 (N_7023,N_5575,N_5412);
nand U7024 (N_7024,N_5041,N_5080);
nand U7025 (N_7025,N_4730,N_5667);
nor U7026 (N_7026,N_4781,N_5290);
or U7027 (N_7027,N_5466,N_5766);
and U7028 (N_7028,N_5412,N_5125);
or U7029 (N_7029,N_5638,N_4924);
nand U7030 (N_7030,N_5596,N_5940);
and U7031 (N_7031,N_4850,N_5463);
or U7032 (N_7032,N_4683,N_5081);
or U7033 (N_7033,N_4766,N_5538);
nand U7034 (N_7034,N_4945,N_4796);
nor U7035 (N_7035,N_5929,N_5605);
or U7036 (N_7036,N_4646,N_5913);
nor U7037 (N_7037,N_4798,N_4667);
or U7038 (N_7038,N_4726,N_5390);
or U7039 (N_7039,N_5352,N_4778);
or U7040 (N_7040,N_5188,N_5943);
xnor U7041 (N_7041,N_5571,N_4896);
nor U7042 (N_7042,N_5891,N_5101);
or U7043 (N_7043,N_4954,N_5433);
xor U7044 (N_7044,N_5708,N_5545);
and U7045 (N_7045,N_5171,N_5706);
nor U7046 (N_7046,N_4522,N_5397);
nand U7047 (N_7047,N_5326,N_5123);
nor U7048 (N_7048,N_5323,N_4803);
nand U7049 (N_7049,N_4795,N_4914);
nand U7050 (N_7050,N_5537,N_5362);
and U7051 (N_7051,N_4925,N_5219);
nor U7052 (N_7052,N_4563,N_5099);
nor U7053 (N_7053,N_5725,N_4627);
or U7054 (N_7054,N_5024,N_5553);
or U7055 (N_7055,N_4811,N_5322);
and U7056 (N_7056,N_5064,N_5556);
xor U7057 (N_7057,N_5473,N_4783);
nand U7058 (N_7058,N_5187,N_5561);
nor U7059 (N_7059,N_4889,N_4718);
or U7060 (N_7060,N_5589,N_5232);
nand U7061 (N_7061,N_5303,N_5613);
nor U7062 (N_7062,N_5436,N_4620);
nand U7063 (N_7063,N_5791,N_5518);
or U7064 (N_7064,N_5392,N_4505);
and U7065 (N_7065,N_5025,N_5271);
and U7066 (N_7066,N_4857,N_5413);
or U7067 (N_7067,N_5168,N_5091);
xor U7068 (N_7068,N_4632,N_5011);
nor U7069 (N_7069,N_5428,N_5179);
xor U7070 (N_7070,N_5542,N_4880);
nand U7071 (N_7071,N_4573,N_4664);
and U7072 (N_7072,N_5220,N_4916);
or U7073 (N_7073,N_5279,N_4584);
or U7074 (N_7074,N_4584,N_5491);
nand U7075 (N_7075,N_4976,N_5667);
nor U7076 (N_7076,N_4801,N_5094);
nor U7077 (N_7077,N_5714,N_5098);
or U7078 (N_7078,N_4974,N_5884);
and U7079 (N_7079,N_4557,N_5133);
nor U7080 (N_7080,N_5738,N_4734);
or U7081 (N_7081,N_5865,N_4681);
and U7082 (N_7082,N_5797,N_5825);
nand U7083 (N_7083,N_5332,N_4949);
nor U7084 (N_7084,N_5345,N_5227);
and U7085 (N_7085,N_5723,N_4691);
and U7086 (N_7086,N_5679,N_5027);
nand U7087 (N_7087,N_4623,N_5448);
and U7088 (N_7088,N_4992,N_4711);
and U7089 (N_7089,N_5924,N_4673);
and U7090 (N_7090,N_4641,N_5141);
nor U7091 (N_7091,N_5031,N_5451);
and U7092 (N_7092,N_5609,N_5094);
and U7093 (N_7093,N_5349,N_4682);
or U7094 (N_7094,N_4644,N_5077);
nand U7095 (N_7095,N_5941,N_5892);
or U7096 (N_7096,N_5099,N_5538);
nand U7097 (N_7097,N_5423,N_4789);
nand U7098 (N_7098,N_5720,N_4922);
nand U7099 (N_7099,N_5424,N_4582);
or U7100 (N_7100,N_5546,N_5381);
nor U7101 (N_7101,N_4728,N_5999);
or U7102 (N_7102,N_5469,N_5918);
nand U7103 (N_7103,N_4586,N_5525);
nor U7104 (N_7104,N_5805,N_4737);
nand U7105 (N_7105,N_4510,N_4974);
or U7106 (N_7106,N_5780,N_5744);
or U7107 (N_7107,N_4829,N_5809);
nand U7108 (N_7108,N_5737,N_5163);
or U7109 (N_7109,N_5503,N_5965);
and U7110 (N_7110,N_4721,N_5506);
xor U7111 (N_7111,N_5647,N_4706);
and U7112 (N_7112,N_4923,N_5170);
nor U7113 (N_7113,N_4768,N_5607);
and U7114 (N_7114,N_4870,N_5634);
and U7115 (N_7115,N_5369,N_4830);
nand U7116 (N_7116,N_4777,N_5463);
and U7117 (N_7117,N_4740,N_4625);
nor U7118 (N_7118,N_5190,N_4895);
and U7119 (N_7119,N_5247,N_5525);
nand U7120 (N_7120,N_5471,N_4519);
nor U7121 (N_7121,N_4906,N_5598);
xnor U7122 (N_7122,N_5728,N_5693);
nor U7123 (N_7123,N_5790,N_4656);
nor U7124 (N_7124,N_4877,N_5000);
and U7125 (N_7125,N_5385,N_5788);
nand U7126 (N_7126,N_4716,N_5509);
nor U7127 (N_7127,N_4919,N_4657);
and U7128 (N_7128,N_5112,N_5121);
nand U7129 (N_7129,N_5788,N_5093);
nand U7130 (N_7130,N_5739,N_5550);
nand U7131 (N_7131,N_5514,N_4676);
nor U7132 (N_7132,N_5094,N_5830);
and U7133 (N_7133,N_5065,N_5536);
nor U7134 (N_7134,N_5556,N_4732);
nand U7135 (N_7135,N_5619,N_5757);
nand U7136 (N_7136,N_4826,N_5567);
or U7137 (N_7137,N_5317,N_5054);
or U7138 (N_7138,N_5259,N_5246);
or U7139 (N_7139,N_4734,N_4813);
or U7140 (N_7140,N_5448,N_4928);
nor U7141 (N_7141,N_5293,N_4727);
and U7142 (N_7142,N_5149,N_5176);
nor U7143 (N_7143,N_4728,N_5479);
nand U7144 (N_7144,N_5133,N_4564);
nand U7145 (N_7145,N_5232,N_4666);
xnor U7146 (N_7146,N_5941,N_5637);
and U7147 (N_7147,N_5365,N_5292);
or U7148 (N_7148,N_4907,N_5117);
nand U7149 (N_7149,N_5907,N_5259);
nand U7150 (N_7150,N_5746,N_4998);
nand U7151 (N_7151,N_5105,N_4591);
nor U7152 (N_7152,N_5710,N_4613);
or U7153 (N_7153,N_5356,N_4648);
nor U7154 (N_7154,N_5197,N_4563);
nor U7155 (N_7155,N_5956,N_5369);
or U7156 (N_7156,N_4669,N_4550);
or U7157 (N_7157,N_5372,N_5597);
xor U7158 (N_7158,N_5198,N_5381);
nor U7159 (N_7159,N_5564,N_4598);
nand U7160 (N_7160,N_5767,N_5283);
and U7161 (N_7161,N_4506,N_5297);
or U7162 (N_7162,N_4570,N_4836);
xor U7163 (N_7163,N_5379,N_4880);
nor U7164 (N_7164,N_4811,N_5362);
and U7165 (N_7165,N_5030,N_5791);
nand U7166 (N_7166,N_5621,N_4589);
or U7167 (N_7167,N_5802,N_5022);
xnor U7168 (N_7168,N_5197,N_4938);
and U7169 (N_7169,N_4845,N_4762);
xor U7170 (N_7170,N_4575,N_5802);
or U7171 (N_7171,N_5031,N_5685);
and U7172 (N_7172,N_4801,N_4802);
or U7173 (N_7173,N_5077,N_5566);
nand U7174 (N_7174,N_5224,N_4847);
nor U7175 (N_7175,N_5715,N_5420);
or U7176 (N_7176,N_5988,N_5269);
nand U7177 (N_7177,N_4844,N_5866);
or U7178 (N_7178,N_4629,N_5223);
nand U7179 (N_7179,N_4853,N_5131);
and U7180 (N_7180,N_5094,N_5275);
xor U7181 (N_7181,N_5646,N_4966);
and U7182 (N_7182,N_5733,N_5917);
nand U7183 (N_7183,N_5573,N_5060);
nand U7184 (N_7184,N_5646,N_4712);
nor U7185 (N_7185,N_4688,N_5971);
and U7186 (N_7186,N_5826,N_5639);
or U7187 (N_7187,N_4932,N_4862);
nor U7188 (N_7188,N_4890,N_4819);
nand U7189 (N_7189,N_5231,N_4813);
and U7190 (N_7190,N_5880,N_5245);
xor U7191 (N_7191,N_5103,N_5819);
and U7192 (N_7192,N_5703,N_5915);
and U7193 (N_7193,N_5655,N_4783);
nor U7194 (N_7194,N_5397,N_5199);
and U7195 (N_7195,N_5804,N_4992);
or U7196 (N_7196,N_4589,N_4994);
and U7197 (N_7197,N_4985,N_5878);
and U7198 (N_7198,N_5164,N_5135);
or U7199 (N_7199,N_5581,N_5859);
nor U7200 (N_7200,N_4539,N_5514);
or U7201 (N_7201,N_5602,N_5015);
or U7202 (N_7202,N_4839,N_5067);
nor U7203 (N_7203,N_4882,N_5390);
nand U7204 (N_7204,N_4553,N_4751);
or U7205 (N_7205,N_5525,N_5982);
nor U7206 (N_7206,N_4806,N_4830);
and U7207 (N_7207,N_5910,N_5890);
and U7208 (N_7208,N_4677,N_4842);
nand U7209 (N_7209,N_5692,N_4945);
nor U7210 (N_7210,N_5164,N_4629);
nor U7211 (N_7211,N_5568,N_5295);
and U7212 (N_7212,N_4610,N_4549);
and U7213 (N_7213,N_5186,N_4919);
or U7214 (N_7214,N_4512,N_5795);
nand U7215 (N_7215,N_4627,N_4634);
nand U7216 (N_7216,N_4927,N_5575);
and U7217 (N_7217,N_5883,N_4790);
nand U7218 (N_7218,N_5237,N_4694);
nand U7219 (N_7219,N_5633,N_5086);
nand U7220 (N_7220,N_5813,N_5769);
nand U7221 (N_7221,N_5219,N_4896);
or U7222 (N_7222,N_4513,N_5773);
and U7223 (N_7223,N_5830,N_5138);
nand U7224 (N_7224,N_5626,N_4537);
nor U7225 (N_7225,N_5117,N_5276);
nand U7226 (N_7226,N_4600,N_5230);
or U7227 (N_7227,N_5448,N_5918);
xor U7228 (N_7228,N_5376,N_4559);
nand U7229 (N_7229,N_5968,N_5226);
or U7230 (N_7230,N_5074,N_5209);
and U7231 (N_7231,N_5070,N_5025);
nor U7232 (N_7232,N_5812,N_4934);
and U7233 (N_7233,N_5118,N_5245);
nor U7234 (N_7234,N_5778,N_5559);
and U7235 (N_7235,N_5512,N_4954);
and U7236 (N_7236,N_4552,N_5755);
nand U7237 (N_7237,N_5685,N_5402);
or U7238 (N_7238,N_5817,N_5620);
and U7239 (N_7239,N_4701,N_4697);
or U7240 (N_7240,N_5405,N_4904);
nor U7241 (N_7241,N_5243,N_4699);
nand U7242 (N_7242,N_5021,N_5342);
and U7243 (N_7243,N_5247,N_4672);
xor U7244 (N_7244,N_5173,N_4952);
nand U7245 (N_7245,N_5020,N_5405);
or U7246 (N_7246,N_5149,N_5623);
and U7247 (N_7247,N_5029,N_5129);
and U7248 (N_7248,N_5875,N_5814);
nor U7249 (N_7249,N_5576,N_5018);
and U7250 (N_7250,N_5979,N_5633);
nand U7251 (N_7251,N_5040,N_5028);
nor U7252 (N_7252,N_5906,N_5210);
nor U7253 (N_7253,N_5200,N_4922);
xnor U7254 (N_7254,N_5495,N_4969);
nor U7255 (N_7255,N_5785,N_4737);
nand U7256 (N_7256,N_4704,N_5690);
and U7257 (N_7257,N_5926,N_5377);
and U7258 (N_7258,N_5229,N_5578);
or U7259 (N_7259,N_5995,N_5837);
nor U7260 (N_7260,N_5342,N_5520);
and U7261 (N_7261,N_5202,N_4983);
and U7262 (N_7262,N_4779,N_5323);
and U7263 (N_7263,N_5628,N_4985);
and U7264 (N_7264,N_4782,N_4968);
nor U7265 (N_7265,N_4670,N_4737);
nand U7266 (N_7266,N_4804,N_4535);
and U7267 (N_7267,N_4747,N_5174);
or U7268 (N_7268,N_4866,N_5990);
xor U7269 (N_7269,N_5862,N_5508);
nor U7270 (N_7270,N_5167,N_5282);
or U7271 (N_7271,N_5357,N_5398);
and U7272 (N_7272,N_5324,N_5167);
or U7273 (N_7273,N_4533,N_5980);
nand U7274 (N_7274,N_4726,N_5722);
and U7275 (N_7275,N_5849,N_4532);
nand U7276 (N_7276,N_5523,N_5050);
and U7277 (N_7277,N_5213,N_4763);
and U7278 (N_7278,N_5142,N_5079);
nor U7279 (N_7279,N_5347,N_4923);
and U7280 (N_7280,N_5380,N_5463);
or U7281 (N_7281,N_5248,N_4952);
and U7282 (N_7282,N_4992,N_5720);
nor U7283 (N_7283,N_5423,N_5163);
nand U7284 (N_7284,N_5362,N_5431);
or U7285 (N_7285,N_5991,N_5484);
nor U7286 (N_7286,N_4746,N_4761);
or U7287 (N_7287,N_4800,N_5680);
or U7288 (N_7288,N_5352,N_5042);
nor U7289 (N_7289,N_5358,N_5853);
xor U7290 (N_7290,N_4801,N_4948);
nand U7291 (N_7291,N_5239,N_5163);
nor U7292 (N_7292,N_4660,N_4987);
and U7293 (N_7293,N_5264,N_5041);
and U7294 (N_7294,N_5112,N_4599);
nand U7295 (N_7295,N_5832,N_5855);
or U7296 (N_7296,N_5586,N_5654);
xor U7297 (N_7297,N_5844,N_4657);
and U7298 (N_7298,N_5495,N_4895);
nor U7299 (N_7299,N_5034,N_5684);
nand U7300 (N_7300,N_5286,N_4579);
or U7301 (N_7301,N_4886,N_5661);
and U7302 (N_7302,N_5626,N_5326);
nand U7303 (N_7303,N_5566,N_5974);
or U7304 (N_7304,N_4501,N_4585);
xor U7305 (N_7305,N_4507,N_5513);
nor U7306 (N_7306,N_5042,N_5682);
or U7307 (N_7307,N_4866,N_5036);
xor U7308 (N_7308,N_4766,N_4655);
nand U7309 (N_7309,N_5020,N_5822);
nand U7310 (N_7310,N_5544,N_5905);
and U7311 (N_7311,N_5748,N_4528);
and U7312 (N_7312,N_4976,N_5257);
and U7313 (N_7313,N_5760,N_5324);
and U7314 (N_7314,N_5227,N_5077);
or U7315 (N_7315,N_4912,N_4955);
nand U7316 (N_7316,N_5207,N_5742);
nand U7317 (N_7317,N_4603,N_4762);
nor U7318 (N_7318,N_4681,N_5548);
nor U7319 (N_7319,N_5649,N_4598);
nand U7320 (N_7320,N_5903,N_5416);
nand U7321 (N_7321,N_5630,N_4675);
and U7322 (N_7322,N_5194,N_5490);
nand U7323 (N_7323,N_4989,N_5346);
nor U7324 (N_7324,N_5392,N_5995);
nand U7325 (N_7325,N_4694,N_5156);
nor U7326 (N_7326,N_5857,N_5537);
xnor U7327 (N_7327,N_4596,N_5690);
and U7328 (N_7328,N_4933,N_5463);
and U7329 (N_7329,N_4886,N_5852);
nand U7330 (N_7330,N_5950,N_5093);
xor U7331 (N_7331,N_5332,N_4588);
nor U7332 (N_7332,N_4554,N_4764);
nor U7333 (N_7333,N_4652,N_5021);
or U7334 (N_7334,N_5095,N_4611);
and U7335 (N_7335,N_4960,N_4646);
or U7336 (N_7336,N_5604,N_5158);
nand U7337 (N_7337,N_5700,N_4581);
xnor U7338 (N_7338,N_4950,N_5237);
nand U7339 (N_7339,N_4892,N_5593);
or U7340 (N_7340,N_5857,N_4523);
nor U7341 (N_7341,N_5331,N_5066);
nor U7342 (N_7342,N_5762,N_5131);
nand U7343 (N_7343,N_4940,N_5813);
or U7344 (N_7344,N_5150,N_5895);
nand U7345 (N_7345,N_5751,N_4745);
or U7346 (N_7346,N_5040,N_5102);
nand U7347 (N_7347,N_5820,N_5267);
or U7348 (N_7348,N_5912,N_5426);
and U7349 (N_7349,N_5615,N_5378);
nand U7350 (N_7350,N_5166,N_5136);
and U7351 (N_7351,N_5059,N_5272);
xnor U7352 (N_7352,N_5011,N_5882);
nand U7353 (N_7353,N_4833,N_5393);
nand U7354 (N_7354,N_5768,N_5744);
and U7355 (N_7355,N_5438,N_4577);
or U7356 (N_7356,N_5638,N_5750);
and U7357 (N_7357,N_5970,N_5213);
nor U7358 (N_7358,N_5242,N_5344);
or U7359 (N_7359,N_5640,N_5167);
and U7360 (N_7360,N_4818,N_4682);
xor U7361 (N_7361,N_5858,N_5721);
nor U7362 (N_7362,N_4710,N_5994);
and U7363 (N_7363,N_5625,N_5837);
nor U7364 (N_7364,N_4754,N_4951);
xor U7365 (N_7365,N_4995,N_5796);
nand U7366 (N_7366,N_5917,N_4563);
or U7367 (N_7367,N_5718,N_5517);
and U7368 (N_7368,N_5242,N_5554);
or U7369 (N_7369,N_5953,N_4521);
xnor U7370 (N_7370,N_4920,N_4531);
and U7371 (N_7371,N_5515,N_4561);
and U7372 (N_7372,N_5183,N_5903);
nor U7373 (N_7373,N_5479,N_5991);
nor U7374 (N_7374,N_5744,N_4947);
and U7375 (N_7375,N_5636,N_5319);
nor U7376 (N_7376,N_5240,N_5218);
nand U7377 (N_7377,N_5397,N_4716);
and U7378 (N_7378,N_5207,N_5584);
nor U7379 (N_7379,N_5639,N_4941);
and U7380 (N_7380,N_5112,N_5299);
or U7381 (N_7381,N_4742,N_5332);
nor U7382 (N_7382,N_4517,N_4805);
and U7383 (N_7383,N_4502,N_5335);
nor U7384 (N_7384,N_5368,N_4663);
xnor U7385 (N_7385,N_4823,N_5965);
nand U7386 (N_7386,N_5023,N_5405);
nand U7387 (N_7387,N_5619,N_5211);
nor U7388 (N_7388,N_5483,N_5070);
nand U7389 (N_7389,N_5447,N_4727);
nand U7390 (N_7390,N_5332,N_4994);
or U7391 (N_7391,N_5059,N_5973);
nand U7392 (N_7392,N_5575,N_4828);
nand U7393 (N_7393,N_5412,N_5901);
and U7394 (N_7394,N_4607,N_5958);
or U7395 (N_7395,N_5919,N_5991);
and U7396 (N_7396,N_5528,N_4642);
nor U7397 (N_7397,N_4856,N_5108);
and U7398 (N_7398,N_4930,N_5768);
and U7399 (N_7399,N_4636,N_5233);
nand U7400 (N_7400,N_5540,N_4748);
nand U7401 (N_7401,N_5401,N_5247);
nor U7402 (N_7402,N_4550,N_4610);
nor U7403 (N_7403,N_5620,N_4752);
nor U7404 (N_7404,N_5829,N_4773);
and U7405 (N_7405,N_5076,N_4552);
and U7406 (N_7406,N_5106,N_4999);
nor U7407 (N_7407,N_5874,N_5309);
nand U7408 (N_7408,N_4742,N_5933);
or U7409 (N_7409,N_5005,N_5881);
or U7410 (N_7410,N_4512,N_5193);
nand U7411 (N_7411,N_4992,N_4984);
and U7412 (N_7412,N_4821,N_5986);
or U7413 (N_7413,N_5461,N_5656);
xnor U7414 (N_7414,N_5221,N_4669);
and U7415 (N_7415,N_5464,N_4990);
and U7416 (N_7416,N_4833,N_4830);
or U7417 (N_7417,N_5709,N_4884);
nand U7418 (N_7418,N_4991,N_5134);
or U7419 (N_7419,N_5469,N_5612);
and U7420 (N_7420,N_5549,N_5289);
nand U7421 (N_7421,N_4803,N_5396);
nand U7422 (N_7422,N_5174,N_5125);
or U7423 (N_7423,N_5610,N_4690);
nand U7424 (N_7424,N_5835,N_5769);
and U7425 (N_7425,N_4569,N_5467);
or U7426 (N_7426,N_5337,N_5208);
or U7427 (N_7427,N_5802,N_5797);
and U7428 (N_7428,N_5698,N_5905);
xor U7429 (N_7429,N_5475,N_4809);
nor U7430 (N_7430,N_5485,N_5751);
or U7431 (N_7431,N_4838,N_5612);
nor U7432 (N_7432,N_4973,N_5499);
nand U7433 (N_7433,N_4683,N_5645);
or U7434 (N_7434,N_5169,N_4588);
or U7435 (N_7435,N_5143,N_5098);
nor U7436 (N_7436,N_4957,N_5490);
nor U7437 (N_7437,N_4544,N_4901);
and U7438 (N_7438,N_5139,N_4805);
or U7439 (N_7439,N_5304,N_5774);
nand U7440 (N_7440,N_5199,N_5860);
nand U7441 (N_7441,N_5793,N_5318);
or U7442 (N_7442,N_5263,N_4590);
or U7443 (N_7443,N_4635,N_4894);
and U7444 (N_7444,N_5989,N_4632);
and U7445 (N_7445,N_4502,N_5379);
nor U7446 (N_7446,N_5447,N_4641);
nand U7447 (N_7447,N_5020,N_5881);
nand U7448 (N_7448,N_5219,N_5419);
xnor U7449 (N_7449,N_4948,N_5876);
or U7450 (N_7450,N_5984,N_4780);
nor U7451 (N_7451,N_5386,N_4948);
or U7452 (N_7452,N_5635,N_4811);
and U7453 (N_7453,N_5776,N_5087);
xnor U7454 (N_7454,N_5440,N_4927);
nand U7455 (N_7455,N_5254,N_5729);
nor U7456 (N_7456,N_5778,N_4568);
and U7457 (N_7457,N_4810,N_5840);
nand U7458 (N_7458,N_5769,N_4890);
nor U7459 (N_7459,N_5845,N_5745);
xor U7460 (N_7460,N_5047,N_4611);
and U7461 (N_7461,N_5599,N_5186);
nand U7462 (N_7462,N_4795,N_5435);
and U7463 (N_7463,N_5282,N_5871);
and U7464 (N_7464,N_4558,N_4657);
or U7465 (N_7465,N_5647,N_4623);
nor U7466 (N_7466,N_5196,N_5872);
and U7467 (N_7467,N_4550,N_4799);
and U7468 (N_7468,N_5277,N_5729);
or U7469 (N_7469,N_5963,N_5351);
or U7470 (N_7470,N_5060,N_5727);
nand U7471 (N_7471,N_5549,N_5704);
nor U7472 (N_7472,N_5912,N_5046);
or U7473 (N_7473,N_5059,N_4930);
nand U7474 (N_7474,N_4939,N_4636);
nor U7475 (N_7475,N_4623,N_4601);
nand U7476 (N_7476,N_5980,N_4683);
and U7477 (N_7477,N_4820,N_4754);
and U7478 (N_7478,N_5909,N_4517);
nand U7479 (N_7479,N_5368,N_5790);
and U7480 (N_7480,N_4505,N_5200);
nor U7481 (N_7481,N_4727,N_4561);
or U7482 (N_7482,N_4767,N_4635);
nor U7483 (N_7483,N_5283,N_5468);
nor U7484 (N_7484,N_5043,N_5766);
and U7485 (N_7485,N_4767,N_5672);
xor U7486 (N_7486,N_4714,N_5343);
or U7487 (N_7487,N_5380,N_4632);
and U7488 (N_7488,N_4989,N_5199);
and U7489 (N_7489,N_5060,N_5629);
and U7490 (N_7490,N_4856,N_4772);
nand U7491 (N_7491,N_5394,N_4680);
and U7492 (N_7492,N_5192,N_5208);
or U7493 (N_7493,N_5850,N_5797);
and U7494 (N_7494,N_5555,N_5864);
nor U7495 (N_7495,N_5218,N_5430);
nor U7496 (N_7496,N_5592,N_4676);
or U7497 (N_7497,N_4711,N_5515);
or U7498 (N_7498,N_5913,N_5355);
and U7499 (N_7499,N_5426,N_5487);
and U7500 (N_7500,N_6065,N_6274);
and U7501 (N_7501,N_7443,N_6938);
or U7502 (N_7502,N_7089,N_6594);
nand U7503 (N_7503,N_6596,N_7447);
and U7504 (N_7504,N_6214,N_6651);
nand U7505 (N_7505,N_6371,N_6471);
nand U7506 (N_7506,N_6438,N_6018);
nand U7507 (N_7507,N_6201,N_6983);
nand U7508 (N_7508,N_6708,N_6827);
nand U7509 (N_7509,N_7318,N_7245);
and U7510 (N_7510,N_6969,N_7000);
nor U7511 (N_7511,N_7257,N_6432);
and U7512 (N_7512,N_7441,N_7128);
and U7513 (N_7513,N_6888,N_6057);
or U7514 (N_7514,N_6038,N_6473);
nor U7515 (N_7515,N_6877,N_6653);
and U7516 (N_7516,N_7383,N_6446);
xnor U7517 (N_7517,N_6093,N_6039);
nand U7518 (N_7518,N_6304,N_6073);
nor U7519 (N_7519,N_7234,N_6428);
nand U7520 (N_7520,N_7141,N_7213);
nand U7521 (N_7521,N_6222,N_7157);
and U7522 (N_7522,N_7220,N_6010);
nand U7523 (N_7523,N_7153,N_7290);
and U7524 (N_7524,N_6531,N_6683);
and U7525 (N_7525,N_6436,N_7082);
nand U7526 (N_7526,N_6617,N_6379);
nor U7527 (N_7527,N_6020,N_6665);
nand U7528 (N_7528,N_6536,N_7097);
and U7529 (N_7529,N_7123,N_6066);
xor U7530 (N_7530,N_6507,N_6814);
and U7531 (N_7531,N_7091,N_7103);
nor U7532 (N_7532,N_6732,N_6560);
nand U7533 (N_7533,N_6481,N_7379);
nand U7534 (N_7534,N_6024,N_7288);
xor U7535 (N_7535,N_6159,N_7171);
nor U7536 (N_7536,N_6794,N_6074);
and U7537 (N_7537,N_6184,N_7325);
nand U7538 (N_7538,N_6144,N_7084);
xor U7539 (N_7539,N_7183,N_6944);
nand U7540 (N_7540,N_6289,N_7155);
or U7541 (N_7541,N_6285,N_6445);
xor U7542 (N_7542,N_7203,N_6994);
nor U7543 (N_7543,N_6405,N_7007);
or U7544 (N_7544,N_6959,N_6303);
xor U7545 (N_7545,N_7148,N_6311);
nand U7546 (N_7546,N_7285,N_7139);
nor U7547 (N_7547,N_6966,N_6764);
or U7548 (N_7548,N_7174,N_6402);
and U7549 (N_7549,N_7254,N_6450);
nor U7550 (N_7550,N_6845,N_6253);
xnor U7551 (N_7551,N_6096,N_6978);
nor U7552 (N_7552,N_7231,N_6566);
and U7553 (N_7553,N_6784,N_6676);
nand U7554 (N_7554,N_6607,N_7436);
or U7555 (N_7555,N_6085,N_7010);
and U7556 (N_7556,N_7466,N_6687);
and U7557 (N_7557,N_7238,N_6633);
or U7558 (N_7558,N_7137,N_7068);
nor U7559 (N_7559,N_6684,N_6142);
nor U7560 (N_7560,N_6156,N_6401);
and U7561 (N_7561,N_7262,N_6133);
xnor U7562 (N_7562,N_6650,N_6023);
and U7563 (N_7563,N_6368,N_6005);
or U7564 (N_7564,N_6451,N_6908);
or U7565 (N_7565,N_7016,N_6170);
or U7566 (N_7566,N_6280,N_7134);
and U7567 (N_7567,N_6858,N_7445);
nor U7568 (N_7568,N_6951,N_7126);
xnor U7569 (N_7569,N_7005,N_6957);
or U7570 (N_7570,N_6677,N_6776);
or U7571 (N_7571,N_6278,N_7277);
nand U7572 (N_7572,N_6734,N_6928);
nor U7573 (N_7573,N_7395,N_7361);
nor U7574 (N_7574,N_6111,N_7145);
and U7575 (N_7575,N_6674,N_6275);
and U7576 (N_7576,N_7184,N_6881);
nor U7577 (N_7577,N_7461,N_6592);
nand U7578 (N_7578,N_6316,N_6931);
and U7579 (N_7579,N_6558,N_6455);
xnor U7580 (N_7580,N_6958,N_6070);
or U7581 (N_7581,N_6069,N_6027);
or U7582 (N_7582,N_7278,N_6487);
nand U7583 (N_7583,N_6341,N_6816);
or U7584 (N_7584,N_7070,N_7198);
or U7585 (N_7585,N_6168,N_7357);
xnor U7586 (N_7586,N_6935,N_6780);
and U7587 (N_7587,N_6079,N_6756);
and U7588 (N_7588,N_6921,N_6661);
or U7589 (N_7589,N_6087,N_7384);
nor U7590 (N_7590,N_6964,N_6392);
and U7591 (N_7591,N_6891,N_7226);
or U7592 (N_7592,N_6916,N_7087);
nor U7593 (N_7593,N_7259,N_7107);
nand U7594 (N_7594,N_7050,N_6895);
nand U7595 (N_7595,N_7022,N_6099);
xnor U7596 (N_7596,N_6228,N_7235);
and U7597 (N_7597,N_6823,N_7094);
or U7598 (N_7598,N_6887,N_6279);
and U7599 (N_7599,N_6801,N_6318);
nand U7600 (N_7600,N_6642,N_7421);
or U7601 (N_7601,N_7410,N_6512);
nor U7602 (N_7602,N_7472,N_6840);
and U7603 (N_7603,N_6656,N_6520);
and U7604 (N_7604,N_6902,N_6897);
and U7605 (N_7605,N_6103,N_6422);
nor U7606 (N_7606,N_6517,N_7402);
xnor U7607 (N_7607,N_6048,N_6768);
nand U7608 (N_7608,N_6165,N_6293);
nand U7609 (N_7609,N_6238,N_7047);
and U7610 (N_7610,N_7268,N_6765);
nor U7611 (N_7611,N_6798,N_6830);
nand U7612 (N_7612,N_6723,N_7434);
and U7613 (N_7613,N_6415,N_6062);
nor U7614 (N_7614,N_6207,N_6197);
or U7615 (N_7615,N_6047,N_6145);
and U7616 (N_7616,N_7215,N_6081);
or U7617 (N_7617,N_6855,N_7041);
and U7618 (N_7618,N_7356,N_6775);
and U7619 (N_7619,N_6488,N_6485);
xnor U7620 (N_7620,N_6680,N_6249);
xnor U7621 (N_7621,N_6766,N_6452);
and U7622 (N_7622,N_7380,N_7192);
and U7623 (N_7623,N_6985,N_6611);
and U7624 (N_7624,N_6094,N_6856);
nand U7625 (N_7625,N_6718,N_6227);
nor U7626 (N_7626,N_7182,N_6540);
and U7627 (N_7627,N_7476,N_6475);
nor U7628 (N_7628,N_7227,N_6792);
nor U7629 (N_7629,N_6970,N_7154);
nor U7630 (N_7630,N_6442,N_7300);
or U7631 (N_7631,N_7400,N_6610);
and U7632 (N_7632,N_7031,N_7081);
or U7633 (N_7633,N_6534,N_7195);
nor U7634 (N_7634,N_7104,N_6853);
nor U7635 (N_7635,N_6456,N_6403);
or U7636 (N_7636,N_6000,N_6230);
nor U7637 (N_7637,N_7149,N_7424);
or U7638 (N_7638,N_6091,N_6878);
and U7639 (N_7639,N_6256,N_7037);
nand U7640 (N_7640,N_6109,N_6625);
and U7641 (N_7641,N_6879,N_7427);
nor U7642 (N_7642,N_7314,N_6180);
or U7643 (N_7643,N_7429,N_6578);
nand U7644 (N_7644,N_7034,N_6905);
nor U7645 (N_7645,N_7164,N_6478);
xnor U7646 (N_7646,N_6444,N_7200);
and U7647 (N_7647,N_6904,N_6961);
xor U7648 (N_7648,N_6510,N_6712);
nand U7649 (N_7649,N_6562,N_6807);
and U7650 (N_7650,N_7111,N_6244);
or U7651 (N_7651,N_6729,N_7260);
or U7652 (N_7652,N_7072,N_7014);
nor U7653 (N_7653,N_6463,N_6051);
nand U7654 (N_7654,N_6396,N_7438);
and U7655 (N_7655,N_7396,N_6364);
nor U7656 (N_7656,N_6545,N_6312);
nand U7657 (N_7657,N_6971,N_7333);
nand U7658 (N_7658,N_6575,N_7376);
and U7659 (N_7659,N_7020,N_7317);
and U7660 (N_7660,N_6567,N_6174);
and U7661 (N_7661,N_6603,N_7113);
or U7662 (N_7662,N_6128,N_6583);
and U7663 (N_7663,N_7054,N_6528);
nand U7664 (N_7664,N_6624,N_6692);
or U7665 (N_7665,N_7003,N_7046);
nand U7666 (N_7666,N_7437,N_6647);
nand U7667 (N_7667,N_6383,N_6299);
nand U7668 (N_7668,N_7147,N_7464);
xnor U7669 (N_7669,N_7100,N_6818);
xnor U7670 (N_7670,N_6115,N_7011);
nor U7671 (N_7671,N_6181,N_6309);
or U7672 (N_7672,N_7355,N_7292);
and U7673 (N_7673,N_7323,N_6516);
nor U7674 (N_7674,N_6532,N_6494);
or U7675 (N_7675,N_7143,N_6548);
or U7676 (N_7676,N_6929,N_6486);
and U7677 (N_7677,N_6581,N_6678);
nor U7678 (N_7678,N_6172,N_6050);
or U7679 (N_7679,N_6060,N_6009);
nor U7680 (N_7680,N_7120,N_6731);
or U7681 (N_7681,N_7482,N_7197);
or U7682 (N_7682,N_6307,N_6715);
nand U7683 (N_7683,N_7255,N_6542);
or U7684 (N_7684,N_6154,N_7144);
nor U7685 (N_7685,N_7353,N_6640);
or U7686 (N_7686,N_6773,N_6913);
xnor U7687 (N_7687,N_6914,N_7112);
and U7688 (N_7688,N_7075,N_7205);
nand U7689 (N_7689,N_7223,N_6835);
xnor U7690 (N_7690,N_6264,N_7276);
and U7691 (N_7691,N_7351,N_6602);
nand U7692 (N_7692,N_6762,N_7105);
nor U7693 (N_7693,N_7418,N_6590);
or U7694 (N_7694,N_6667,N_6454);
nand U7695 (N_7695,N_6740,N_7074);
nand U7696 (N_7696,N_6384,N_6308);
and U7697 (N_7697,N_6591,N_6056);
nand U7698 (N_7698,N_6219,N_7388);
nand U7699 (N_7699,N_6382,N_6441);
and U7700 (N_7700,N_6703,N_6979);
and U7701 (N_7701,N_6988,N_6329);
or U7702 (N_7702,N_6811,N_6063);
and U7703 (N_7703,N_7085,N_7432);
nor U7704 (N_7704,N_7480,N_6385);
nand U7705 (N_7705,N_7341,N_6272);
nand U7706 (N_7706,N_6618,N_7138);
or U7707 (N_7707,N_7258,N_6433);
xnor U7708 (N_7708,N_7252,N_6167);
and U7709 (N_7709,N_6636,N_7228);
nand U7710 (N_7710,N_6090,N_7015);
nand U7711 (N_7711,N_7499,N_7233);
nor U7712 (N_7712,N_6348,N_6470);
or U7713 (N_7713,N_7374,N_6614);
and U7714 (N_7714,N_6083,N_6286);
nor U7715 (N_7715,N_6831,N_6484);
xnor U7716 (N_7716,N_6515,N_6116);
and U7717 (N_7717,N_7495,N_7008);
xor U7718 (N_7718,N_6239,N_7332);
nor U7719 (N_7719,N_7168,N_6263);
and U7720 (N_7720,N_7417,N_7405);
nand U7721 (N_7721,N_6394,N_7090);
nor U7722 (N_7722,N_6287,N_7454);
or U7723 (N_7723,N_6380,N_6414);
nor U7724 (N_7724,N_7284,N_6419);
xnor U7725 (N_7725,N_6034,N_7193);
nor U7726 (N_7726,N_6098,N_6439);
nand U7727 (N_7727,N_6785,N_6637);
nor U7728 (N_7728,N_6924,N_6497);
or U7729 (N_7729,N_6015,N_7267);
and U7730 (N_7730,N_6721,N_7216);
nor U7731 (N_7731,N_6277,N_7142);
and U7732 (N_7732,N_6124,N_7286);
xor U7733 (N_7733,N_6210,N_6421);
nor U7734 (N_7734,N_6118,N_7253);
nand U7735 (N_7735,N_6714,N_6986);
nor U7736 (N_7736,N_6679,N_6948);
nand U7737 (N_7737,N_6499,N_6300);
and U7738 (N_7738,N_7492,N_6584);
or U7739 (N_7739,N_6993,N_6786);
or U7740 (N_7740,N_6072,N_6490);
and U7741 (N_7741,N_6330,N_7140);
or U7742 (N_7742,N_6086,N_6525);
nor U7743 (N_7743,N_6996,N_6870);
and U7744 (N_7744,N_7350,N_7033);
and U7745 (N_7745,N_6854,N_7196);
nor U7746 (N_7746,N_6460,N_6195);
nor U7747 (N_7747,N_7358,N_7251);
or U7748 (N_7748,N_6416,N_6701);
or U7749 (N_7749,N_6121,N_6342);
xnor U7750 (N_7750,N_6459,N_6572);
nor U7751 (N_7751,N_6457,N_6477);
nor U7752 (N_7752,N_6220,N_6291);
nor U7753 (N_7753,N_6612,N_7407);
or U7754 (N_7754,N_7188,N_6351);
nand U7755 (N_7755,N_6990,N_6193);
nand U7756 (N_7756,N_6243,N_6503);
nand U7757 (N_7757,N_6161,N_6643);
nor U7758 (N_7758,N_6907,N_6273);
and U7759 (N_7759,N_7321,N_7056);
nor U7760 (N_7760,N_7224,N_6896);
nor U7761 (N_7761,N_7179,N_7177);
nor U7762 (N_7762,N_6101,N_6231);
or U7763 (N_7763,N_6192,N_7219);
or U7764 (N_7764,N_6354,N_7281);
nor U7765 (N_7765,N_6621,N_7308);
or U7766 (N_7766,N_6114,N_7266);
or U7767 (N_7767,N_7346,N_7398);
nor U7768 (N_7768,N_6390,N_6537);
and U7769 (N_7769,N_6569,N_6530);
nand U7770 (N_7770,N_6875,N_6313);
xor U7771 (N_7771,N_6909,N_6660);
nor U7772 (N_7772,N_6869,N_7039);
nand U7773 (N_7773,N_6587,N_7108);
nand U7774 (N_7774,N_6999,N_7331);
nand U7775 (N_7775,N_6014,N_6725);
xnor U7776 (N_7776,N_6754,N_6557);
nand U7777 (N_7777,N_6003,N_7058);
nand U7778 (N_7778,N_6682,N_6952);
or U7779 (N_7779,N_6209,N_6926);
and U7780 (N_7780,N_6846,N_6864);
nand U7781 (N_7781,N_6568,N_7237);
nand U7782 (N_7782,N_6322,N_6589);
nand U7783 (N_7783,N_6704,N_6898);
nand U7784 (N_7784,N_7060,N_6758);
nor U7785 (N_7785,N_6155,N_6821);
nand U7786 (N_7786,N_6270,N_6779);
and U7787 (N_7787,N_7069,N_6733);
nor U7788 (N_7788,N_6182,N_6685);
or U7789 (N_7789,N_7449,N_7368);
xor U7790 (N_7790,N_6886,N_6406);
nor U7791 (N_7791,N_7294,N_6746);
nor U7792 (N_7792,N_7017,N_6054);
or U7793 (N_7793,N_6426,N_6315);
and U7794 (N_7794,N_6523,N_6737);
nor U7795 (N_7795,N_6186,N_6113);
or U7796 (N_7796,N_7389,N_6302);
or U7797 (N_7797,N_7280,N_6839);
nor U7798 (N_7798,N_7488,N_6500);
and U7799 (N_7799,N_7435,N_6011);
nand U7800 (N_7800,N_6213,N_6296);
xor U7801 (N_7801,N_6828,N_7404);
nand U7802 (N_7802,N_6799,N_6972);
nor U7803 (N_7803,N_6707,N_6218);
nor U7804 (N_7804,N_6565,N_7282);
and U7805 (N_7805,N_7204,N_6190);
nand U7806 (N_7806,N_6325,N_7027);
or U7807 (N_7807,N_6912,N_7159);
and U7808 (N_7808,N_6947,N_6026);
nor U7809 (N_7809,N_7324,N_7354);
and U7810 (N_7810,N_6435,N_7293);
nor U7811 (N_7811,N_7067,N_7044);
or U7812 (N_7812,N_7176,N_6346);
or U7813 (N_7813,N_6755,N_6321);
or U7814 (N_7814,N_7337,N_7130);
nand U7815 (N_7815,N_6409,N_6104);
nand U7816 (N_7816,N_7412,N_6025);
and U7817 (N_7817,N_6205,N_6388);
nand U7818 (N_7818,N_7116,N_7269);
nor U7819 (N_7819,N_6608,N_6769);
and U7820 (N_7820,N_6224,N_6783);
nor U7821 (N_7821,N_7287,N_6787);
or U7822 (N_7822,N_6634,N_6899);
or U7823 (N_7823,N_6453,N_6880);
nor U7824 (N_7824,N_6847,N_6395);
and U7825 (N_7825,N_6225,N_7403);
nor U7826 (N_7826,N_6489,N_6071);
and U7827 (N_7827,N_6204,N_7099);
and U7828 (N_7828,N_6082,N_6750);
nand U7829 (N_7829,N_6593,N_6366);
nand U7830 (N_7830,N_6804,N_7250);
or U7831 (N_7831,N_6652,N_7343);
or U7832 (N_7832,N_6177,N_6255);
nand U7833 (N_7833,N_6246,N_7001);
or U7834 (N_7834,N_6805,N_7040);
and U7835 (N_7835,N_6882,N_6049);
and U7836 (N_7836,N_6012,N_6981);
or U7837 (N_7837,N_7475,N_6851);
and U7838 (N_7838,N_7261,N_6915);
nor U7839 (N_7839,N_7018,N_7129);
and U7840 (N_7840,N_7484,N_7271);
and U7841 (N_7841,N_7092,N_6713);
nor U7842 (N_7842,N_7439,N_7497);
and U7843 (N_7843,N_7028,N_6262);
nor U7844 (N_7844,N_6092,N_6447);
nand U7845 (N_7845,N_6495,N_7401);
and U7846 (N_7846,N_6646,N_6501);
and U7847 (N_7847,N_7229,N_7273);
nand U7848 (N_7848,N_6857,N_7232);
or U7849 (N_7849,N_6088,N_6953);
and U7850 (N_7850,N_6350,N_6939);
xnor U7851 (N_7851,N_6788,N_7474);
or U7852 (N_7852,N_7121,N_7026);
and U7853 (N_7853,N_6781,N_6188);
nand U7854 (N_7854,N_6868,N_6389);
nand U7855 (N_7855,N_6859,N_6055);
or U7856 (N_7856,N_6221,N_6730);
xnor U7857 (N_7857,N_6976,N_7481);
nor U7858 (N_7858,N_6203,N_6173);
and U7859 (N_7859,N_7486,N_6185);
and U7860 (N_7860,N_6657,N_6339);
xor U7861 (N_7861,N_6918,N_6335);
xor U7862 (N_7862,N_6358,N_6900);
nand U7863 (N_7863,N_7132,N_6372);
nor U7864 (N_7864,N_6808,N_7408);
and U7865 (N_7865,N_6894,N_7265);
or U7866 (N_7866,N_7347,N_6668);
and U7867 (N_7867,N_6705,N_6251);
xor U7868 (N_7868,N_6605,N_7306);
nand U7869 (N_7869,N_7217,N_6240);
or U7870 (N_7870,N_6564,N_6910);
nand U7871 (N_7871,N_7342,N_6694);
and U7872 (N_7872,N_6053,N_7411);
and U7873 (N_7873,N_6247,N_6283);
or U7874 (N_7874,N_7024,N_6458);
nor U7875 (N_7875,N_7391,N_6550);
nand U7876 (N_7876,N_6982,N_7124);
and U7877 (N_7877,N_7275,N_6582);
and U7878 (N_7878,N_6361,N_6942);
or U7879 (N_7879,N_7369,N_6196);
and U7880 (N_7880,N_7473,N_7344);
nand U7881 (N_7881,N_6007,N_7460);
nand U7882 (N_7882,N_6355,N_6615);
nor U7883 (N_7883,N_7419,N_6386);
nor U7884 (N_7884,N_6340,N_6298);
and U7885 (N_7885,N_6949,N_6077);
xor U7886 (N_7886,N_6535,N_6100);
and U7887 (N_7887,N_7161,N_7249);
and U7888 (N_7888,N_7242,N_7088);
and U7889 (N_7889,N_7002,N_6613);
and U7890 (N_7890,N_6266,N_6043);
and U7891 (N_7891,N_7201,N_6029);
and U7892 (N_7892,N_6268,N_6987);
nor U7893 (N_7893,N_7185,N_6719);
nor U7894 (N_7894,N_7209,N_6427);
nand U7895 (N_7895,N_7352,N_7448);
or U7896 (N_7896,N_7025,N_7365);
nor U7897 (N_7897,N_7326,N_6008);
and U7898 (N_7898,N_6626,N_7079);
or U7899 (N_7899,N_6774,N_7319);
or U7900 (N_7900,N_7338,N_6136);
nor U7901 (N_7901,N_6521,N_7426);
nor U7902 (N_7902,N_7021,N_6362);
nand U7903 (N_7903,N_6089,N_6843);
nand U7904 (N_7904,N_6338,N_7189);
xnor U7905 (N_7905,N_6932,N_6373);
or U7906 (N_7906,N_7225,N_6940);
xor U7907 (N_7907,N_6695,N_6398);
or U7908 (N_7908,N_6261,N_7372);
xnor U7909 (N_7909,N_7119,N_6825);
and U7910 (N_7910,N_6127,N_7366);
or U7911 (N_7911,N_6215,N_7377);
nand U7912 (N_7912,N_6199,N_6374);
and U7913 (N_7913,N_6876,N_7106);
or U7914 (N_7914,N_6666,N_7178);
nand U7915 (N_7915,N_6138,N_7425);
nor U7916 (N_7916,N_7152,N_6276);
nand U7917 (N_7917,N_6933,N_6058);
nand U7918 (N_7918,N_7236,N_6620);
nor U7919 (N_7919,N_7243,N_6526);
or U7920 (N_7920,N_6601,N_6871);
and U7921 (N_7921,N_6954,N_7162);
nand U7922 (N_7922,N_6002,N_7078);
nor U7923 (N_7923,N_6748,N_7470);
or U7924 (N_7924,N_6693,N_6906);
or U7925 (N_7925,N_7452,N_6706);
xnor U7926 (N_7926,N_7221,N_7298);
and U7927 (N_7927,N_6559,N_6553);
nor U7928 (N_7928,N_6789,N_6194);
nand U7929 (N_7929,N_6377,N_6429);
and U7930 (N_7930,N_7468,N_6849);
nor U7931 (N_7931,N_7459,N_6519);
and U7932 (N_7932,N_6709,N_6102);
xnor U7933 (N_7933,N_6006,N_7030);
and U7934 (N_7934,N_6597,N_7309);
nand U7935 (N_7935,N_6033,N_6357);
and U7936 (N_7936,N_7127,N_6604);
nand U7937 (N_7937,N_6418,N_7210);
and U7938 (N_7938,N_6749,N_7165);
nand U7939 (N_7939,N_7042,N_6956);
nand U7940 (N_7940,N_7310,N_6742);
nand U7941 (N_7941,N_6367,N_6267);
nand U7942 (N_7942,N_7390,N_6580);
nand U7943 (N_7943,N_6042,N_6290);
nand U7944 (N_7944,N_7095,N_6105);
or U7945 (N_7945,N_6673,N_6645);
and U7946 (N_7946,N_7151,N_6412);
nor U7947 (N_7947,N_6206,N_6934);
nor U7948 (N_7948,N_6397,N_7433);
nor U7949 (N_7949,N_6378,N_6824);
xnor U7950 (N_7950,N_6122,N_6360);
or U7951 (N_7951,N_7212,N_6236);
and U7952 (N_7952,N_6962,N_6506);
and U7953 (N_7953,N_6728,N_6862);
nand U7954 (N_7954,N_7170,N_6662);
nor U7955 (N_7955,N_7431,N_7371);
nor U7956 (N_7956,N_6861,N_7399);
nor U7957 (N_7957,N_6903,N_6237);
and U7958 (N_7958,N_7296,N_6820);
xor U7959 (N_7959,N_6641,N_6152);
nand U7960 (N_7960,N_6717,N_6294);
and U7961 (N_7961,N_6735,N_6872);
nor U7962 (N_7962,N_6430,N_7320);
nor U7963 (N_7963,N_7387,N_6649);
or U7964 (N_7964,N_6356,N_6021);
xnor U7965 (N_7965,N_7264,N_7023);
nor U7966 (N_7966,N_7135,N_6040);
nand U7967 (N_7967,N_6297,N_6822);
nor U7968 (N_7968,N_6370,N_6802);
nor U7969 (N_7969,N_6208,N_6393);
and U7970 (N_7970,N_6157,N_7247);
nor U7971 (N_7971,N_6068,N_6420);
nor U7972 (N_7972,N_7214,N_6538);
xnor U7973 (N_7973,N_6771,N_6585);
nand U7974 (N_7974,N_6777,N_6967);
nand U7975 (N_7975,N_6084,N_6140);
or U7976 (N_7976,N_6920,N_7272);
or U7977 (N_7977,N_6837,N_6211);
or U7978 (N_7978,N_7362,N_7163);
nor U7979 (N_7979,N_7297,N_6977);
xor U7980 (N_7980,N_6245,N_6327);
nand U7981 (N_7981,N_6483,N_6505);
nor U7982 (N_7982,N_6997,N_7180);
nor U7983 (N_7983,N_6659,N_7167);
nand U7984 (N_7984,N_6829,N_7202);
or U7985 (N_7985,N_7334,N_6806);
nand U7986 (N_7986,N_6533,N_6809);
nor U7987 (N_7987,N_7289,N_7455);
and U7988 (N_7988,N_6400,N_7458);
and U7989 (N_7989,N_7175,N_6848);
nor U7990 (N_7990,N_7463,N_6125);
and U7991 (N_7991,N_7240,N_6782);
or U7992 (N_7992,N_6305,N_6844);
or U7993 (N_7993,N_7392,N_6834);
and U7994 (N_7994,N_7316,N_6793);
nor U7995 (N_7995,N_6080,N_7457);
nor U7996 (N_7996,N_6022,N_6555);
and U7997 (N_7997,N_6417,N_7125);
and U7998 (N_7998,N_6153,N_6271);
xnor U7999 (N_7999,N_6711,N_7160);
nand U8000 (N_8000,N_7446,N_7038);
nor U8001 (N_8001,N_6522,N_6466);
xnor U8002 (N_8002,N_6130,N_6045);
nand U8003 (N_8003,N_6097,N_7048);
xnor U8004 (N_8004,N_6465,N_7156);
xnor U8005 (N_8005,N_7146,N_7057);
and U8006 (N_8006,N_6328,N_7328);
or U8007 (N_8007,N_6689,N_7363);
and U8008 (N_8008,N_7440,N_6893);
or U8009 (N_8009,N_6107,N_6013);
nor U8010 (N_8010,N_7348,N_6151);
and U8011 (N_8011,N_7397,N_6509);
nand U8012 (N_8012,N_6376,N_6573);
nand U8013 (N_8013,N_7246,N_7494);
nor U8014 (N_8014,N_6233,N_6778);
and U8015 (N_8015,N_7222,N_7349);
and U8016 (N_8016,N_6627,N_6179);
or U8017 (N_8017,N_6937,N_6336);
or U8018 (N_8018,N_7239,N_7420);
or U8019 (N_8019,N_6075,N_6654);
or U8020 (N_8020,N_6320,N_6158);
nand U8021 (N_8021,N_6187,N_7327);
nand U8022 (N_8022,N_6556,N_6763);
and U8023 (N_8023,N_6235,N_6129);
nand U8024 (N_8024,N_6472,N_6681);
or U8025 (N_8025,N_6036,N_6968);
nor U8026 (N_8026,N_6698,N_7430);
or U8027 (N_8027,N_6301,N_6757);
or U8028 (N_8028,N_6600,N_6044);
and U8029 (N_8029,N_6984,N_6425);
nor U8030 (N_8030,N_6817,N_6663);
or U8031 (N_8031,N_6028,N_6198);
nor U8032 (N_8032,N_6539,N_6606);
or U8033 (N_8033,N_6306,N_6690);
xnor U8034 (N_8034,N_7409,N_6178);
and U8035 (N_8035,N_7471,N_6745);
xor U8036 (N_8036,N_6200,N_6797);
or U8037 (N_8037,N_6697,N_6016);
and U8038 (N_8038,N_7049,N_6365);
or U8039 (N_8039,N_6404,N_6992);
or U8040 (N_8040,N_7248,N_6874);
and U8041 (N_8041,N_6126,N_6106);
nor U8042 (N_8042,N_7364,N_6216);
nor U8043 (N_8043,N_6059,N_7115);
nor U8044 (N_8044,N_6212,N_6139);
nand U8045 (N_8045,N_7444,N_7322);
nand U8046 (N_8046,N_6443,N_6511);
nor U8047 (N_8047,N_6175,N_6078);
nand U8048 (N_8048,N_6284,N_6310);
and U8049 (N_8049,N_6541,N_6696);
and U8050 (N_8050,N_6836,N_7076);
and U8051 (N_8051,N_7462,N_6399);
nor U8052 (N_8052,N_7062,N_7263);
nor U8053 (N_8053,N_6479,N_6669);
nor U8054 (N_8054,N_6169,N_6448);
nand U8055 (N_8055,N_6759,N_6037);
nand U8056 (N_8056,N_6588,N_7393);
nor U8057 (N_8057,N_6727,N_6381);
or U8058 (N_8058,N_7491,N_7329);
xnor U8059 (N_8059,N_6469,N_6767);
nand U8060 (N_8060,N_6547,N_6543);
nand U8061 (N_8061,N_7206,N_6146);
nor U8062 (N_8062,N_6493,N_7406);
nand U8063 (N_8063,N_6137,N_6226);
and U8064 (N_8064,N_7498,N_6884);
xnor U8065 (N_8065,N_6349,N_6975);
or U8066 (N_8066,N_7299,N_6945);
nand U8067 (N_8067,N_6061,N_7181);
nand U8068 (N_8068,N_6946,N_6032);
or U8069 (N_8069,N_6770,N_7312);
nand U8070 (N_8070,N_7375,N_7065);
and U8071 (N_8071,N_6234,N_6440);
or U8072 (N_8072,N_6574,N_7133);
nand U8073 (N_8073,N_7093,N_6551);
and U8074 (N_8074,N_6973,N_6630);
nor U8075 (N_8075,N_6867,N_7493);
nor U8076 (N_8076,N_6260,N_6616);
nor U8077 (N_8077,N_7051,N_6282);
and U8078 (N_8078,N_7013,N_7467);
nor U8079 (N_8079,N_6960,N_7194);
nand U8080 (N_8080,N_6810,N_6549);
or U8081 (N_8081,N_6710,N_6826);
nand U8082 (N_8082,N_6554,N_7360);
nand U8083 (N_8083,N_6259,N_6747);
nand U8084 (N_8084,N_6004,N_6344);
nand U8085 (N_8085,N_6424,N_6974);
nor U8086 (N_8086,N_6726,N_6108);
nand U8087 (N_8087,N_6700,N_6552);
xor U8088 (N_8088,N_6191,N_6223);
and U8089 (N_8089,N_6019,N_6334);
nand U8090 (N_8090,N_7045,N_7098);
nand U8091 (N_8091,N_6150,N_6164);
nand U8092 (N_8092,N_6671,N_7102);
nand U8093 (N_8093,N_6434,N_6248);
nor U8094 (N_8094,N_7230,N_6563);
and U8095 (N_8095,N_6132,N_7279);
and U8096 (N_8096,N_7169,N_6595);
nor U8097 (N_8097,N_7428,N_6281);
nand U8098 (N_8098,N_6609,N_7118);
and U8099 (N_8099,N_7313,N_7301);
and U8100 (N_8100,N_6323,N_6866);
and U8101 (N_8101,N_7330,N_7077);
or U8102 (N_8102,N_6135,N_6675);
and U8103 (N_8103,N_6319,N_6850);
or U8104 (N_8104,N_6664,N_6119);
nand U8105 (N_8105,N_7053,N_6720);
and U8106 (N_8106,N_6265,N_6407);
xnor U8107 (N_8107,N_7373,N_6217);
or U8108 (N_8108,N_6258,N_7066);
nor U8109 (N_8109,N_7370,N_6250);
nor U8110 (N_8110,N_6885,N_6639);
and U8111 (N_8111,N_6148,N_6317);
or U8112 (N_8112,N_7186,N_6739);
or U8113 (N_8113,N_6923,N_6468);
and U8114 (N_8114,N_6041,N_6347);
nand U8115 (N_8115,N_6925,N_7256);
xnor U8116 (N_8116,N_7218,N_7442);
xnor U8117 (N_8117,N_6922,N_6324);
nor U8118 (N_8118,N_6352,N_6691);
nor U8119 (N_8119,N_6067,N_7414);
or U8120 (N_8120,N_6638,N_6699);
and U8121 (N_8121,N_7291,N_6513);
and U8122 (N_8122,N_6369,N_6702);
and U8123 (N_8123,N_6995,N_6752);
and U8124 (N_8124,N_7035,N_7304);
and U8125 (N_8125,N_7340,N_6670);
nand U8126 (N_8126,N_6819,N_7339);
or U8127 (N_8127,N_6269,N_6579);
nand U8128 (N_8128,N_7423,N_7422);
or U8129 (N_8129,N_6813,N_6524);
nor U8130 (N_8130,N_7083,N_6842);
and U8131 (N_8131,N_6431,N_7483);
nand U8132 (N_8132,N_6254,N_6387);
or U8133 (N_8133,N_6760,N_6860);
nor U8134 (N_8134,N_6901,N_6546);
xnor U8135 (N_8135,N_6648,N_7073);
nand U8136 (N_8136,N_7009,N_7019);
nand U8137 (N_8137,N_6252,N_6744);
nor U8138 (N_8138,N_6017,N_7208);
nand U8139 (N_8139,N_6833,N_6736);
and U8140 (N_8140,N_6686,N_6359);
and U8141 (N_8141,N_7190,N_6189);
nand U8142 (N_8142,N_7150,N_6927);
nand U8143 (N_8143,N_6658,N_6919);
nand U8144 (N_8144,N_6772,N_6232);
nor U8145 (N_8145,N_6391,N_6980);
nand U8146 (N_8146,N_7052,N_6076);
nand U8147 (N_8147,N_6331,N_7465);
nor U8148 (N_8148,N_7315,N_7345);
and U8149 (N_8149,N_6411,N_6716);
and U8150 (N_8150,N_7490,N_6134);
or U8151 (N_8151,N_7311,N_6464);
nor U8152 (N_8152,N_6800,N_6795);
nand U8153 (N_8153,N_6120,N_7451);
nor U8154 (N_8154,N_6889,N_6337);
nand U8155 (N_8155,N_6815,N_6117);
and U8156 (N_8156,N_7131,N_7036);
nor U8157 (N_8157,N_6644,N_6408);
or U8158 (N_8158,N_6461,N_6865);
or U8159 (N_8159,N_6753,N_6035);
and U8160 (N_8160,N_6936,N_6295);
or U8161 (N_8161,N_6527,N_6143);
nand U8162 (N_8162,N_7158,N_7136);
and U8163 (N_8163,N_6635,N_7477);
nor U8164 (N_8164,N_7335,N_6176);
or U8165 (N_8165,N_6599,N_6110);
or U8166 (N_8166,N_6561,N_6672);
nand U8167 (N_8167,N_7478,N_6046);
and U8168 (N_8168,N_6943,N_6229);
nor U8169 (N_8169,N_6803,N_6571);
nor U8170 (N_8170,N_6911,N_7378);
and U8171 (N_8171,N_7485,N_7096);
nand U8172 (N_8172,N_6498,N_6941);
or U8173 (N_8173,N_7063,N_7110);
or U8174 (N_8174,N_6375,N_6480);
nor U8175 (N_8175,N_6838,N_7367);
nor U8176 (N_8176,N_6363,N_6462);
nor U8177 (N_8177,N_7117,N_6655);
nor U8178 (N_8178,N_6123,N_6183);
or U8179 (N_8179,N_6332,N_7244);
nand U8180 (N_8180,N_6241,N_6989);
nor U8181 (N_8181,N_6492,N_7270);
or U8182 (N_8182,N_6623,N_6504);
or U8183 (N_8183,N_7453,N_6288);
nand U8184 (N_8184,N_7385,N_6141);
or U8185 (N_8185,N_6688,N_6345);
and U8186 (N_8186,N_6622,N_6529);
or U8187 (N_8187,N_6991,N_6171);
xor U8188 (N_8188,N_7307,N_6852);
or U8189 (N_8189,N_7283,N_6883);
nor U8190 (N_8190,N_7064,N_7416);
nand U8191 (N_8191,N_7114,N_6724);
nand U8192 (N_8192,N_6491,N_6518);
nand U8193 (N_8193,N_6950,N_6052);
nand U8194 (N_8194,N_6413,N_6095);
nor U8195 (N_8195,N_7302,N_6314);
nor U8196 (N_8196,N_6064,N_6632);
xnor U8197 (N_8197,N_6570,N_6812);
nor U8198 (N_8198,N_6131,N_6410);
and U8199 (N_8199,N_6514,N_6292);
or U8200 (N_8200,N_6343,N_6163);
nor U8201 (N_8201,N_6738,N_7241);
or U8202 (N_8202,N_6147,N_6963);
nor U8203 (N_8203,N_6791,N_6751);
nor U8204 (N_8204,N_7191,N_6202);
nor U8205 (N_8205,N_7211,N_7456);
nor U8206 (N_8206,N_6722,N_6326);
nor U8207 (N_8207,N_6955,N_7469);
nor U8208 (N_8208,N_7295,N_7055);
nand U8209 (N_8209,N_7336,N_6333);
xnor U8210 (N_8210,N_6631,N_6892);
and U8211 (N_8211,N_7303,N_7274);
xnor U8212 (N_8212,N_7382,N_6628);
nor U8213 (N_8213,N_6743,N_7059);
nand U8214 (N_8214,N_6476,N_6965);
and U8215 (N_8215,N_6160,N_7043);
nor U8216 (N_8216,N_7415,N_6437);
and U8217 (N_8217,N_6930,N_7487);
nand U8218 (N_8218,N_6741,N_6619);
nand U8219 (N_8219,N_7012,N_6761);
nor U8220 (N_8220,N_7032,N_6031);
nand U8221 (N_8221,N_6482,N_7101);
nor U8222 (N_8222,N_6449,N_6577);
nand U8223 (N_8223,N_6576,N_6502);
xor U8224 (N_8224,N_6586,N_6508);
and U8225 (N_8225,N_7381,N_6790);
nand U8226 (N_8226,N_6841,N_6873);
and U8227 (N_8227,N_6353,N_7173);
or U8228 (N_8228,N_7496,N_7109);
and U8229 (N_8229,N_6998,N_6863);
and U8230 (N_8230,N_7450,N_6166);
nor U8231 (N_8231,N_7413,N_7029);
nor U8232 (N_8232,N_7479,N_6917);
and U8233 (N_8233,N_6112,N_6598);
nand U8234 (N_8234,N_6001,N_6890);
and U8235 (N_8235,N_7086,N_6474);
nor U8236 (N_8236,N_7305,N_6030);
nor U8237 (N_8237,N_6162,N_7187);
and U8238 (N_8238,N_6149,N_6467);
nand U8239 (N_8239,N_7489,N_7359);
and U8240 (N_8240,N_7071,N_7004);
nand U8241 (N_8241,N_6242,N_6629);
nor U8242 (N_8242,N_7006,N_6257);
nand U8243 (N_8243,N_7207,N_6423);
or U8244 (N_8244,N_6832,N_6796);
nor U8245 (N_8245,N_7394,N_6496);
nand U8246 (N_8246,N_7386,N_6544);
or U8247 (N_8247,N_7172,N_7080);
and U8248 (N_8248,N_7166,N_7199);
nor U8249 (N_8249,N_7061,N_7122);
nor U8250 (N_8250,N_7431,N_6383);
and U8251 (N_8251,N_6135,N_6790);
or U8252 (N_8252,N_6754,N_7013);
or U8253 (N_8253,N_6204,N_7401);
or U8254 (N_8254,N_6567,N_6173);
nor U8255 (N_8255,N_6254,N_6933);
or U8256 (N_8256,N_6959,N_6413);
or U8257 (N_8257,N_7244,N_6080);
nand U8258 (N_8258,N_7136,N_7321);
nor U8259 (N_8259,N_6151,N_7321);
or U8260 (N_8260,N_6889,N_6845);
and U8261 (N_8261,N_7065,N_6767);
or U8262 (N_8262,N_6918,N_6059);
xnor U8263 (N_8263,N_7086,N_6713);
or U8264 (N_8264,N_6996,N_7212);
or U8265 (N_8265,N_7076,N_6854);
xor U8266 (N_8266,N_6433,N_6929);
xor U8267 (N_8267,N_7491,N_6042);
or U8268 (N_8268,N_7008,N_7012);
nor U8269 (N_8269,N_6729,N_7108);
nand U8270 (N_8270,N_7333,N_7334);
nor U8271 (N_8271,N_6510,N_7461);
or U8272 (N_8272,N_7262,N_6004);
nand U8273 (N_8273,N_6455,N_6672);
and U8274 (N_8274,N_6458,N_6877);
nor U8275 (N_8275,N_6561,N_7183);
nor U8276 (N_8276,N_6826,N_6913);
and U8277 (N_8277,N_6534,N_6336);
nor U8278 (N_8278,N_7171,N_7220);
nor U8279 (N_8279,N_6275,N_6423);
nor U8280 (N_8280,N_6964,N_7318);
and U8281 (N_8281,N_6875,N_7183);
and U8282 (N_8282,N_6356,N_6694);
xnor U8283 (N_8283,N_6744,N_7364);
or U8284 (N_8284,N_6439,N_7318);
xor U8285 (N_8285,N_6564,N_6312);
nor U8286 (N_8286,N_6792,N_7068);
and U8287 (N_8287,N_7221,N_6966);
and U8288 (N_8288,N_6435,N_6598);
nor U8289 (N_8289,N_7151,N_7309);
and U8290 (N_8290,N_6192,N_6010);
nor U8291 (N_8291,N_6918,N_7145);
nor U8292 (N_8292,N_7381,N_7108);
xor U8293 (N_8293,N_7321,N_6141);
nand U8294 (N_8294,N_7381,N_7291);
nor U8295 (N_8295,N_6439,N_7149);
and U8296 (N_8296,N_7193,N_6304);
and U8297 (N_8297,N_7019,N_6343);
nor U8298 (N_8298,N_6183,N_6868);
or U8299 (N_8299,N_6074,N_6320);
nor U8300 (N_8300,N_6102,N_6442);
and U8301 (N_8301,N_7231,N_6724);
nor U8302 (N_8302,N_6843,N_6264);
or U8303 (N_8303,N_6757,N_6755);
and U8304 (N_8304,N_7404,N_7057);
nand U8305 (N_8305,N_7356,N_7400);
and U8306 (N_8306,N_6409,N_6469);
or U8307 (N_8307,N_6667,N_6760);
nor U8308 (N_8308,N_6856,N_7165);
or U8309 (N_8309,N_6490,N_6999);
nor U8310 (N_8310,N_6751,N_6748);
nor U8311 (N_8311,N_6333,N_6004);
nand U8312 (N_8312,N_6694,N_7330);
nor U8313 (N_8313,N_6082,N_6955);
nor U8314 (N_8314,N_6511,N_6082);
nand U8315 (N_8315,N_6252,N_6153);
or U8316 (N_8316,N_6821,N_6124);
or U8317 (N_8317,N_7108,N_6475);
and U8318 (N_8318,N_7311,N_6637);
or U8319 (N_8319,N_6682,N_6323);
and U8320 (N_8320,N_6743,N_7454);
and U8321 (N_8321,N_7479,N_6658);
and U8322 (N_8322,N_6535,N_6025);
xnor U8323 (N_8323,N_7062,N_7125);
nor U8324 (N_8324,N_7436,N_6418);
or U8325 (N_8325,N_7018,N_6910);
nor U8326 (N_8326,N_6793,N_6710);
or U8327 (N_8327,N_6495,N_6600);
nand U8328 (N_8328,N_6421,N_6366);
nor U8329 (N_8329,N_6459,N_7119);
nor U8330 (N_8330,N_6818,N_7356);
or U8331 (N_8331,N_6033,N_6017);
nand U8332 (N_8332,N_7220,N_7221);
nor U8333 (N_8333,N_6855,N_6967);
and U8334 (N_8334,N_6024,N_6979);
nand U8335 (N_8335,N_7373,N_6878);
or U8336 (N_8336,N_6509,N_6870);
and U8337 (N_8337,N_6820,N_7308);
or U8338 (N_8338,N_6342,N_7158);
nand U8339 (N_8339,N_6748,N_6238);
nor U8340 (N_8340,N_6335,N_6352);
nor U8341 (N_8341,N_6602,N_7470);
nor U8342 (N_8342,N_6071,N_7411);
nand U8343 (N_8343,N_6682,N_7323);
nor U8344 (N_8344,N_7043,N_7175);
xnor U8345 (N_8345,N_6776,N_6162);
nand U8346 (N_8346,N_7028,N_7330);
nand U8347 (N_8347,N_7303,N_6938);
nand U8348 (N_8348,N_7035,N_7488);
xor U8349 (N_8349,N_7153,N_7171);
nand U8350 (N_8350,N_6703,N_6715);
or U8351 (N_8351,N_6847,N_7259);
or U8352 (N_8352,N_7261,N_6912);
xor U8353 (N_8353,N_7125,N_7106);
nand U8354 (N_8354,N_7343,N_7103);
and U8355 (N_8355,N_7046,N_6681);
and U8356 (N_8356,N_7404,N_6907);
nand U8357 (N_8357,N_6224,N_7499);
nor U8358 (N_8358,N_6486,N_6166);
or U8359 (N_8359,N_6671,N_6485);
and U8360 (N_8360,N_7290,N_6122);
or U8361 (N_8361,N_6249,N_7278);
or U8362 (N_8362,N_6891,N_6354);
nand U8363 (N_8363,N_7065,N_6554);
and U8364 (N_8364,N_6604,N_6938);
or U8365 (N_8365,N_6537,N_6018);
nand U8366 (N_8366,N_6038,N_6880);
nand U8367 (N_8367,N_7227,N_7136);
or U8368 (N_8368,N_7108,N_6569);
nand U8369 (N_8369,N_6939,N_6666);
or U8370 (N_8370,N_6810,N_7167);
and U8371 (N_8371,N_6893,N_6566);
or U8372 (N_8372,N_7470,N_6459);
xor U8373 (N_8373,N_6550,N_7075);
nand U8374 (N_8374,N_6767,N_7091);
or U8375 (N_8375,N_6299,N_7336);
and U8376 (N_8376,N_6203,N_6308);
nor U8377 (N_8377,N_6556,N_7316);
xor U8378 (N_8378,N_7020,N_6489);
nand U8379 (N_8379,N_6393,N_6888);
nand U8380 (N_8380,N_6048,N_7396);
nor U8381 (N_8381,N_6452,N_6883);
or U8382 (N_8382,N_7031,N_7383);
nand U8383 (N_8383,N_6673,N_6727);
and U8384 (N_8384,N_6981,N_7431);
or U8385 (N_8385,N_7120,N_7239);
nor U8386 (N_8386,N_7472,N_6542);
or U8387 (N_8387,N_7053,N_7100);
nand U8388 (N_8388,N_6684,N_6779);
and U8389 (N_8389,N_6792,N_7226);
and U8390 (N_8390,N_6342,N_7480);
and U8391 (N_8391,N_6787,N_6213);
nor U8392 (N_8392,N_6047,N_7254);
or U8393 (N_8393,N_6065,N_7302);
and U8394 (N_8394,N_6733,N_7208);
and U8395 (N_8395,N_6993,N_7408);
or U8396 (N_8396,N_6330,N_6140);
nand U8397 (N_8397,N_7052,N_7296);
or U8398 (N_8398,N_6476,N_7486);
or U8399 (N_8399,N_6575,N_6184);
or U8400 (N_8400,N_6100,N_7221);
nor U8401 (N_8401,N_7430,N_6862);
nor U8402 (N_8402,N_6838,N_7461);
or U8403 (N_8403,N_6708,N_7265);
nor U8404 (N_8404,N_6702,N_6139);
or U8405 (N_8405,N_7488,N_7107);
and U8406 (N_8406,N_7264,N_6882);
and U8407 (N_8407,N_6559,N_7083);
and U8408 (N_8408,N_7244,N_7103);
xnor U8409 (N_8409,N_6249,N_7126);
nor U8410 (N_8410,N_6660,N_6049);
or U8411 (N_8411,N_7386,N_6254);
nand U8412 (N_8412,N_6318,N_6268);
nor U8413 (N_8413,N_6618,N_7223);
or U8414 (N_8414,N_7194,N_7115);
and U8415 (N_8415,N_6402,N_6451);
or U8416 (N_8416,N_6068,N_6748);
or U8417 (N_8417,N_6320,N_6708);
nand U8418 (N_8418,N_6242,N_6187);
nor U8419 (N_8419,N_7377,N_6895);
or U8420 (N_8420,N_6230,N_6685);
or U8421 (N_8421,N_6055,N_6846);
or U8422 (N_8422,N_6636,N_7430);
and U8423 (N_8423,N_7229,N_7005);
nor U8424 (N_8424,N_7220,N_7148);
and U8425 (N_8425,N_6082,N_6245);
nor U8426 (N_8426,N_7407,N_6258);
or U8427 (N_8427,N_7429,N_6642);
or U8428 (N_8428,N_7303,N_7430);
nor U8429 (N_8429,N_7368,N_6301);
nand U8430 (N_8430,N_6827,N_6865);
and U8431 (N_8431,N_7273,N_7323);
nand U8432 (N_8432,N_6414,N_6861);
xnor U8433 (N_8433,N_6843,N_6119);
nor U8434 (N_8434,N_7435,N_6676);
nand U8435 (N_8435,N_6606,N_6511);
and U8436 (N_8436,N_7108,N_6921);
or U8437 (N_8437,N_7066,N_6244);
xnor U8438 (N_8438,N_7468,N_6493);
and U8439 (N_8439,N_6605,N_7037);
nor U8440 (N_8440,N_6401,N_6086);
and U8441 (N_8441,N_7082,N_6244);
or U8442 (N_8442,N_7058,N_6594);
xnor U8443 (N_8443,N_6178,N_6456);
or U8444 (N_8444,N_7352,N_6320);
nor U8445 (N_8445,N_6830,N_7157);
xor U8446 (N_8446,N_6721,N_6636);
and U8447 (N_8447,N_7225,N_6427);
nand U8448 (N_8448,N_6002,N_7469);
nor U8449 (N_8449,N_6452,N_6084);
nand U8450 (N_8450,N_6606,N_6601);
or U8451 (N_8451,N_6676,N_6768);
and U8452 (N_8452,N_6052,N_6742);
nand U8453 (N_8453,N_6404,N_7468);
xor U8454 (N_8454,N_7002,N_6328);
and U8455 (N_8455,N_7447,N_7167);
and U8456 (N_8456,N_6357,N_6244);
xnor U8457 (N_8457,N_6999,N_7373);
nand U8458 (N_8458,N_6143,N_7402);
or U8459 (N_8459,N_6000,N_6914);
nor U8460 (N_8460,N_6715,N_6508);
nor U8461 (N_8461,N_6590,N_6903);
nand U8462 (N_8462,N_6139,N_6394);
and U8463 (N_8463,N_6205,N_6586);
nand U8464 (N_8464,N_6419,N_6839);
xnor U8465 (N_8465,N_6708,N_7290);
nor U8466 (N_8466,N_6127,N_7377);
or U8467 (N_8467,N_6338,N_6691);
nor U8468 (N_8468,N_6662,N_6722);
or U8469 (N_8469,N_6643,N_7238);
and U8470 (N_8470,N_7098,N_6457);
nor U8471 (N_8471,N_6090,N_7221);
nor U8472 (N_8472,N_6516,N_6058);
xor U8473 (N_8473,N_7424,N_7458);
and U8474 (N_8474,N_6735,N_7299);
xor U8475 (N_8475,N_6283,N_7462);
and U8476 (N_8476,N_6304,N_6613);
and U8477 (N_8477,N_7132,N_7417);
or U8478 (N_8478,N_6294,N_6827);
xor U8479 (N_8479,N_7461,N_6835);
xnor U8480 (N_8480,N_6386,N_6160);
xnor U8481 (N_8481,N_6182,N_7269);
and U8482 (N_8482,N_7418,N_7314);
nor U8483 (N_8483,N_6888,N_6222);
xnor U8484 (N_8484,N_7377,N_6051);
or U8485 (N_8485,N_7107,N_6760);
nand U8486 (N_8486,N_7028,N_7093);
xnor U8487 (N_8487,N_6608,N_7055);
nor U8488 (N_8488,N_6067,N_6525);
nor U8489 (N_8489,N_7357,N_6844);
nand U8490 (N_8490,N_6882,N_6212);
and U8491 (N_8491,N_7445,N_6438);
and U8492 (N_8492,N_6319,N_7325);
nand U8493 (N_8493,N_7131,N_6888);
nor U8494 (N_8494,N_7498,N_7152);
nand U8495 (N_8495,N_6582,N_6384);
xnor U8496 (N_8496,N_6828,N_6311);
xnor U8497 (N_8497,N_6367,N_6086);
or U8498 (N_8498,N_7008,N_6227);
and U8499 (N_8499,N_6707,N_6099);
xnor U8500 (N_8500,N_6046,N_6949);
and U8501 (N_8501,N_7331,N_6119);
nand U8502 (N_8502,N_6212,N_6539);
and U8503 (N_8503,N_6043,N_7326);
or U8504 (N_8504,N_6968,N_7374);
or U8505 (N_8505,N_6463,N_7115);
or U8506 (N_8506,N_7076,N_6630);
nand U8507 (N_8507,N_6433,N_7495);
or U8508 (N_8508,N_6595,N_7491);
or U8509 (N_8509,N_6314,N_6861);
or U8510 (N_8510,N_6649,N_6536);
nor U8511 (N_8511,N_6747,N_6107);
nand U8512 (N_8512,N_6739,N_6632);
or U8513 (N_8513,N_6660,N_7089);
or U8514 (N_8514,N_6945,N_6650);
nand U8515 (N_8515,N_6946,N_6233);
nand U8516 (N_8516,N_6319,N_6363);
nor U8517 (N_8517,N_7225,N_6699);
and U8518 (N_8518,N_6711,N_6159);
and U8519 (N_8519,N_6350,N_6286);
or U8520 (N_8520,N_6982,N_7328);
nand U8521 (N_8521,N_6462,N_7353);
nor U8522 (N_8522,N_6839,N_7023);
nor U8523 (N_8523,N_6220,N_6232);
and U8524 (N_8524,N_7068,N_6353);
nand U8525 (N_8525,N_7347,N_7385);
xor U8526 (N_8526,N_7326,N_6595);
xor U8527 (N_8527,N_7162,N_7045);
nor U8528 (N_8528,N_7409,N_6202);
and U8529 (N_8529,N_7239,N_6505);
nor U8530 (N_8530,N_6673,N_6803);
or U8531 (N_8531,N_6902,N_6683);
or U8532 (N_8532,N_7486,N_6451);
xnor U8533 (N_8533,N_6468,N_6099);
and U8534 (N_8534,N_6580,N_7076);
nor U8535 (N_8535,N_7490,N_7270);
nand U8536 (N_8536,N_6084,N_6713);
or U8537 (N_8537,N_6012,N_7144);
nand U8538 (N_8538,N_6849,N_6779);
xor U8539 (N_8539,N_7359,N_7131);
nand U8540 (N_8540,N_6276,N_6832);
and U8541 (N_8541,N_6358,N_6065);
and U8542 (N_8542,N_7473,N_7443);
or U8543 (N_8543,N_6199,N_7320);
or U8544 (N_8544,N_6931,N_6661);
nor U8545 (N_8545,N_7040,N_6586);
nor U8546 (N_8546,N_6614,N_6492);
nor U8547 (N_8547,N_7150,N_6003);
nand U8548 (N_8548,N_7175,N_6855);
and U8549 (N_8549,N_6081,N_6485);
nor U8550 (N_8550,N_6966,N_6658);
and U8551 (N_8551,N_7396,N_6459);
and U8552 (N_8552,N_6724,N_6497);
nand U8553 (N_8553,N_6857,N_6494);
nand U8554 (N_8554,N_7498,N_6999);
or U8555 (N_8555,N_6122,N_7151);
nand U8556 (N_8556,N_7145,N_6882);
nor U8557 (N_8557,N_7204,N_6429);
and U8558 (N_8558,N_7467,N_7214);
and U8559 (N_8559,N_6578,N_6346);
and U8560 (N_8560,N_6463,N_6959);
nor U8561 (N_8561,N_6841,N_6352);
nor U8562 (N_8562,N_6399,N_7155);
and U8563 (N_8563,N_7046,N_7081);
nor U8564 (N_8564,N_6923,N_6748);
xor U8565 (N_8565,N_7223,N_7450);
nor U8566 (N_8566,N_6661,N_6157);
nor U8567 (N_8567,N_6655,N_6795);
nor U8568 (N_8568,N_6376,N_6808);
and U8569 (N_8569,N_6610,N_6491);
or U8570 (N_8570,N_6152,N_6742);
nand U8571 (N_8571,N_6579,N_7240);
nor U8572 (N_8572,N_6733,N_6575);
and U8573 (N_8573,N_6032,N_7386);
nand U8574 (N_8574,N_6840,N_6650);
nand U8575 (N_8575,N_6991,N_6347);
nor U8576 (N_8576,N_7091,N_7282);
and U8577 (N_8577,N_7144,N_6441);
and U8578 (N_8578,N_7071,N_7070);
and U8579 (N_8579,N_7284,N_6689);
nor U8580 (N_8580,N_6994,N_7052);
nand U8581 (N_8581,N_6749,N_6271);
and U8582 (N_8582,N_6372,N_6040);
nor U8583 (N_8583,N_7266,N_7452);
and U8584 (N_8584,N_7366,N_6951);
and U8585 (N_8585,N_6496,N_7431);
nor U8586 (N_8586,N_6394,N_6578);
nor U8587 (N_8587,N_6313,N_6523);
and U8588 (N_8588,N_6088,N_6125);
nand U8589 (N_8589,N_7130,N_6400);
and U8590 (N_8590,N_7380,N_6449);
or U8591 (N_8591,N_6058,N_6453);
or U8592 (N_8592,N_6417,N_6936);
or U8593 (N_8593,N_7156,N_6078);
nor U8594 (N_8594,N_7323,N_7259);
nor U8595 (N_8595,N_6873,N_6134);
nor U8596 (N_8596,N_6613,N_6280);
and U8597 (N_8597,N_6830,N_6158);
and U8598 (N_8598,N_6435,N_6332);
xnor U8599 (N_8599,N_6517,N_6738);
and U8600 (N_8600,N_6541,N_6495);
or U8601 (N_8601,N_6748,N_6735);
and U8602 (N_8602,N_6191,N_6204);
or U8603 (N_8603,N_6316,N_6424);
nor U8604 (N_8604,N_6833,N_6312);
nand U8605 (N_8605,N_6024,N_6033);
xnor U8606 (N_8606,N_6672,N_6241);
and U8607 (N_8607,N_7429,N_6429);
xor U8608 (N_8608,N_6676,N_7081);
and U8609 (N_8609,N_6258,N_6757);
or U8610 (N_8610,N_7097,N_7455);
and U8611 (N_8611,N_6573,N_6593);
and U8612 (N_8612,N_6483,N_7020);
or U8613 (N_8613,N_7062,N_6657);
nor U8614 (N_8614,N_6784,N_6460);
or U8615 (N_8615,N_6944,N_6097);
nor U8616 (N_8616,N_7379,N_6321);
nor U8617 (N_8617,N_6802,N_6708);
or U8618 (N_8618,N_6306,N_6547);
and U8619 (N_8619,N_6012,N_7042);
xnor U8620 (N_8620,N_7197,N_6883);
nand U8621 (N_8621,N_6203,N_7218);
nor U8622 (N_8622,N_6762,N_6446);
nand U8623 (N_8623,N_6900,N_7007);
or U8624 (N_8624,N_6872,N_6517);
and U8625 (N_8625,N_7054,N_6326);
or U8626 (N_8626,N_7192,N_6363);
and U8627 (N_8627,N_7383,N_7308);
and U8628 (N_8628,N_7217,N_6152);
or U8629 (N_8629,N_7280,N_6568);
or U8630 (N_8630,N_6534,N_6928);
nor U8631 (N_8631,N_6280,N_6098);
nor U8632 (N_8632,N_6462,N_6263);
nor U8633 (N_8633,N_6634,N_7473);
nor U8634 (N_8634,N_6135,N_6978);
nand U8635 (N_8635,N_7458,N_6828);
nor U8636 (N_8636,N_6429,N_7292);
and U8637 (N_8637,N_6853,N_7127);
nor U8638 (N_8638,N_6197,N_6691);
nor U8639 (N_8639,N_6519,N_7436);
nand U8640 (N_8640,N_6423,N_6408);
xnor U8641 (N_8641,N_6593,N_6921);
and U8642 (N_8642,N_6202,N_6562);
or U8643 (N_8643,N_6925,N_6739);
nor U8644 (N_8644,N_7045,N_6954);
xor U8645 (N_8645,N_7258,N_6242);
xnor U8646 (N_8646,N_7389,N_6756);
nor U8647 (N_8647,N_7258,N_7096);
xnor U8648 (N_8648,N_6108,N_6207);
and U8649 (N_8649,N_7212,N_6361);
or U8650 (N_8650,N_6221,N_7345);
nor U8651 (N_8651,N_7233,N_7257);
nand U8652 (N_8652,N_7456,N_7495);
or U8653 (N_8653,N_6349,N_7393);
or U8654 (N_8654,N_6331,N_6371);
and U8655 (N_8655,N_6971,N_6547);
or U8656 (N_8656,N_6908,N_6914);
and U8657 (N_8657,N_7235,N_7060);
nor U8658 (N_8658,N_7413,N_7175);
and U8659 (N_8659,N_6054,N_7265);
nor U8660 (N_8660,N_6433,N_6624);
nor U8661 (N_8661,N_6428,N_6395);
nor U8662 (N_8662,N_6180,N_7469);
nand U8663 (N_8663,N_6418,N_7468);
nor U8664 (N_8664,N_6020,N_7318);
nand U8665 (N_8665,N_6169,N_6153);
xnor U8666 (N_8666,N_7327,N_6447);
nand U8667 (N_8667,N_6386,N_6518);
nor U8668 (N_8668,N_7076,N_6967);
nor U8669 (N_8669,N_6930,N_7472);
and U8670 (N_8670,N_7027,N_6716);
and U8671 (N_8671,N_6843,N_6733);
nor U8672 (N_8672,N_7459,N_7382);
and U8673 (N_8673,N_6133,N_6586);
nand U8674 (N_8674,N_7162,N_6005);
nand U8675 (N_8675,N_6506,N_7241);
and U8676 (N_8676,N_7301,N_6663);
or U8677 (N_8677,N_7447,N_7495);
xnor U8678 (N_8678,N_6162,N_7017);
or U8679 (N_8679,N_6255,N_6463);
nor U8680 (N_8680,N_6852,N_6118);
nand U8681 (N_8681,N_6900,N_6512);
nor U8682 (N_8682,N_6860,N_6336);
or U8683 (N_8683,N_6822,N_7341);
and U8684 (N_8684,N_6064,N_6090);
nor U8685 (N_8685,N_6258,N_7137);
nor U8686 (N_8686,N_6058,N_7079);
nand U8687 (N_8687,N_7017,N_7483);
nand U8688 (N_8688,N_6995,N_6282);
or U8689 (N_8689,N_7018,N_6076);
nor U8690 (N_8690,N_6438,N_6230);
or U8691 (N_8691,N_7463,N_7338);
nand U8692 (N_8692,N_6584,N_6398);
or U8693 (N_8693,N_6496,N_6701);
xnor U8694 (N_8694,N_6231,N_6453);
nand U8695 (N_8695,N_6730,N_7066);
or U8696 (N_8696,N_7129,N_6902);
and U8697 (N_8697,N_7173,N_7169);
or U8698 (N_8698,N_6064,N_7006);
xnor U8699 (N_8699,N_6409,N_6519);
or U8700 (N_8700,N_6180,N_6685);
nand U8701 (N_8701,N_7157,N_6699);
or U8702 (N_8702,N_7344,N_6810);
nand U8703 (N_8703,N_6114,N_6703);
nor U8704 (N_8704,N_7060,N_7400);
or U8705 (N_8705,N_7419,N_6131);
nand U8706 (N_8706,N_6878,N_6512);
and U8707 (N_8707,N_7221,N_6392);
or U8708 (N_8708,N_6695,N_7173);
nand U8709 (N_8709,N_6773,N_6497);
or U8710 (N_8710,N_7125,N_7070);
nor U8711 (N_8711,N_6956,N_6715);
and U8712 (N_8712,N_7282,N_6071);
or U8713 (N_8713,N_6965,N_7206);
and U8714 (N_8714,N_6979,N_6938);
and U8715 (N_8715,N_7370,N_6353);
xor U8716 (N_8716,N_6447,N_6551);
nor U8717 (N_8717,N_7162,N_7269);
nand U8718 (N_8718,N_6476,N_7461);
or U8719 (N_8719,N_6139,N_7154);
and U8720 (N_8720,N_6175,N_6461);
and U8721 (N_8721,N_6910,N_6056);
and U8722 (N_8722,N_6792,N_7498);
nand U8723 (N_8723,N_6259,N_6503);
and U8724 (N_8724,N_6619,N_6312);
nand U8725 (N_8725,N_6624,N_6217);
or U8726 (N_8726,N_6083,N_6827);
nand U8727 (N_8727,N_7038,N_6149);
nor U8728 (N_8728,N_6649,N_6617);
nand U8729 (N_8729,N_6189,N_7479);
nor U8730 (N_8730,N_6185,N_7293);
nor U8731 (N_8731,N_6188,N_6936);
nand U8732 (N_8732,N_7142,N_6501);
nand U8733 (N_8733,N_6176,N_6810);
or U8734 (N_8734,N_7068,N_6039);
and U8735 (N_8735,N_6039,N_7424);
nand U8736 (N_8736,N_6287,N_7411);
xnor U8737 (N_8737,N_7060,N_6173);
nor U8738 (N_8738,N_6189,N_6269);
and U8739 (N_8739,N_6500,N_7242);
nand U8740 (N_8740,N_6046,N_7284);
nor U8741 (N_8741,N_6869,N_6712);
nand U8742 (N_8742,N_7051,N_7132);
nand U8743 (N_8743,N_7129,N_6665);
nand U8744 (N_8744,N_6826,N_7431);
and U8745 (N_8745,N_6692,N_7165);
xor U8746 (N_8746,N_6186,N_6766);
xor U8747 (N_8747,N_6252,N_6622);
nor U8748 (N_8748,N_6864,N_6872);
nand U8749 (N_8749,N_6865,N_6026);
nand U8750 (N_8750,N_6978,N_6562);
or U8751 (N_8751,N_6240,N_7429);
nor U8752 (N_8752,N_7433,N_6535);
and U8753 (N_8753,N_6731,N_6287);
nand U8754 (N_8754,N_7330,N_6976);
and U8755 (N_8755,N_6818,N_6072);
or U8756 (N_8756,N_6154,N_7099);
and U8757 (N_8757,N_7488,N_6050);
or U8758 (N_8758,N_7403,N_6143);
nand U8759 (N_8759,N_7146,N_6429);
or U8760 (N_8760,N_7330,N_7198);
nand U8761 (N_8761,N_7240,N_6917);
nand U8762 (N_8762,N_6817,N_7431);
nand U8763 (N_8763,N_6075,N_6039);
or U8764 (N_8764,N_6130,N_7497);
nand U8765 (N_8765,N_7081,N_7336);
and U8766 (N_8766,N_6725,N_7251);
nor U8767 (N_8767,N_6796,N_7345);
and U8768 (N_8768,N_6879,N_7406);
and U8769 (N_8769,N_7089,N_6698);
xor U8770 (N_8770,N_6234,N_7077);
or U8771 (N_8771,N_6117,N_7482);
or U8772 (N_8772,N_7235,N_7105);
or U8773 (N_8773,N_6521,N_7335);
nor U8774 (N_8774,N_6079,N_6176);
or U8775 (N_8775,N_6558,N_7023);
and U8776 (N_8776,N_7307,N_7449);
nand U8777 (N_8777,N_6908,N_7446);
nor U8778 (N_8778,N_6099,N_6638);
nor U8779 (N_8779,N_6760,N_6653);
nand U8780 (N_8780,N_6493,N_7318);
nand U8781 (N_8781,N_6368,N_6644);
nand U8782 (N_8782,N_6367,N_6363);
or U8783 (N_8783,N_6514,N_6962);
or U8784 (N_8784,N_6276,N_6031);
nor U8785 (N_8785,N_7124,N_6996);
or U8786 (N_8786,N_6992,N_7218);
nand U8787 (N_8787,N_6793,N_6585);
and U8788 (N_8788,N_6509,N_6767);
or U8789 (N_8789,N_6481,N_7249);
xor U8790 (N_8790,N_7263,N_6771);
nor U8791 (N_8791,N_6028,N_7162);
nor U8792 (N_8792,N_6292,N_6112);
or U8793 (N_8793,N_6268,N_6168);
nand U8794 (N_8794,N_6078,N_6233);
or U8795 (N_8795,N_6099,N_7010);
and U8796 (N_8796,N_6942,N_6033);
or U8797 (N_8797,N_6002,N_7319);
and U8798 (N_8798,N_6507,N_6102);
or U8799 (N_8799,N_6681,N_7282);
and U8800 (N_8800,N_7366,N_7192);
nor U8801 (N_8801,N_7230,N_6012);
nand U8802 (N_8802,N_7366,N_6309);
or U8803 (N_8803,N_6266,N_6862);
nor U8804 (N_8804,N_6788,N_6973);
nor U8805 (N_8805,N_6198,N_6832);
nand U8806 (N_8806,N_7378,N_7171);
and U8807 (N_8807,N_6380,N_6377);
nand U8808 (N_8808,N_6421,N_7285);
xnor U8809 (N_8809,N_6941,N_7197);
nand U8810 (N_8810,N_6943,N_6950);
and U8811 (N_8811,N_7067,N_6028);
and U8812 (N_8812,N_6511,N_6413);
or U8813 (N_8813,N_6587,N_7150);
or U8814 (N_8814,N_7312,N_6849);
or U8815 (N_8815,N_6573,N_6679);
or U8816 (N_8816,N_6178,N_6156);
and U8817 (N_8817,N_6219,N_6698);
nor U8818 (N_8818,N_7019,N_6985);
nor U8819 (N_8819,N_6594,N_7335);
nand U8820 (N_8820,N_6783,N_6671);
or U8821 (N_8821,N_6702,N_6238);
or U8822 (N_8822,N_6979,N_6147);
nand U8823 (N_8823,N_7015,N_6595);
and U8824 (N_8824,N_7042,N_6795);
and U8825 (N_8825,N_6227,N_6848);
nor U8826 (N_8826,N_6781,N_7066);
or U8827 (N_8827,N_7477,N_7403);
nor U8828 (N_8828,N_6030,N_6449);
nand U8829 (N_8829,N_6273,N_7071);
and U8830 (N_8830,N_6440,N_7309);
nor U8831 (N_8831,N_7054,N_6851);
or U8832 (N_8832,N_6219,N_7423);
and U8833 (N_8833,N_7272,N_6788);
nand U8834 (N_8834,N_6996,N_6680);
and U8835 (N_8835,N_7235,N_6037);
or U8836 (N_8836,N_6980,N_6879);
nor U8837 (N_8837,N_6000,N_7119);
and U8838 (N_8838,N_6412,N_6959);
nor U8839 (N_8839,N_7279,N_6160);
xnor U8840 (N_8840,N_7022,N_6315);
nor U8841 (N_8841,N_6980,N_7057);
nand U8842 (N_8842,N_6655,N_7084);
nand U8843 (N_8843,N_6706,N_6083);
or U8844 (N_8844,N_6403,N_6772);
or U8845 (N_8845,N_6894,N_6027);
nor U8846 (N_8846,N_6694,N_6117);
and U8847 (N_8847,N_6067,N_6853);
and U8848 (N_8848,N_7135,N_6615);
nor U8849 (N_8849,N_6745,N_7156);
nor U8850 (N_8850,N_6606,N_6469);
nor U8851 (N_8851,N_7075,N_6747);
and U8852 (N_8852,N_7117,N_6276);
nor U8853 (N_8853,N_7327,N_6996);
nand U8854 (N_8854,N_6261,N_6603);
or U8855 (N_8855,N_6947,N_6562);
nand U8856 (N_8856,N_7259,N_6760);
nand U8857 (N_8857,N_6094,N_6380);
nand U8858 (N_8858,N_7287,N_6094);
and U8859 (N_8859,N_6026,N_6444);
or U8860 (N_8860,N_7329,N_6270);
or U8861 (N_8861,N_6401,N_6284);
and U8862 (N_8862,N_7257,N_6939);
or U8863 (N_8863,N_6195,N_6514);
and U8864 (N_8864,N_6688,N_7134);
nand U8865 (N_8865,N_7325,N_6130);
and U8866 (N_8866,N_6651,N_7039);
nand U8867 (N_8867,N_7001,N_6399);
and U8868 (N_8868,N_6276,N_7310);
nand U8869 (N_8869,N_6758,N_6797);
nor U8870 (N_8870,N_6390,N_6620);
and U8871 (N_8871,N_6910,N_6821);
or U8872 (N_8872,N_6561,N_6060);
nand U8873 (N_8873,N_6946,N_7262);
nor U8874 (N_8874,N_7196,N_6293);
and U8875 (N_8875,N_7125,N_7297);
and U8876 (N_8876,N_6262,N_7298);
xor U8877 (N_8877,N_6893,N_6841);
nand U8878 (N_8878,N_6996,N_7050);
nand U8879 (N_8879,N_7411,N_6546);
nor U8880 (N_8880,N_7083,N_6885);
or U8881 (N_8881,N_6593,N_7449);
or U8882 (N_8882,N_6276,N_6560);
and U8883 (N_8883,N_7193,N_6005);
and U8884 (N_8884,N_6973,N_6714);
nand U8885 (N_8885,N_6969,N_6745);
nand U8886 (N_8886,N_6211,N_7295);
or U8887 (N_8887,N_7478,N_7180);
nor U8888 (N_8888,N_6494,N_7481);
nand U8889 (N_8889,N_6335,N_7197);
and U8890 (N_8890,N_7081,N_7115);
or U8891 (N_8891,N_7303,N_6263);
or U8892 (N_8892,N_6388,N_6326);
nor U8893 (N_8893,N_6571,N_6459);
nand U8894 (N_8894,N_6471,N_6313);
nor U8895 (N_8895,N_6515,N_7128);
and U8896 (N_8896,N_6850,N_7305);
nand U8897 (N_8897,N_7339,N_6784);
and U8898 (N_8898,N_7319,N_6242);
nor U8899 (N_8899,N_6384,N_6446);
and U8900 (N_8900,N_6657,N_6474);
nor U8901 (N_8901,N_6161,N_7259);
xor U8902 (N_8902,N_6917,N_6591);
xnor U8903 (N_8903,N_6179,N_6569);
nand U8904 (N_8904,N_6525,N_6341);
xnor U8905 (N_8905,N_6694,N_7349);
nor U8906 (N_8906,N_6253,N_7302);
or U8907 (N_8907,N_6742,N_6054);
or U8908 (N_8908,N_6676,N_6492);
nor U8909 (N_8909,N_7287,N_6548);
or U8910 (N_8910,N_6274,N_7104);
and U8911 (N_8911,N_6945,N_6515);
nor U8912 (N_8912,N_6916,N_6909);
nor U8913 (N_8913,N_6237,N_7320);
and U8914 (N_8914,N_7387,N_6166);
nor U8915 (N_8915,N_6087,N_7385);
nand U8916 (N_8916,N_6490,N_7453);
and U8917 (N_8917,N_6605,N_6043);
and U8918 (N_8918,N_6706,N_7422);
or U8919 (N_8919,N_6621,N_6731);
and U8920 (N_8920,N_7132,N_7329);
nand U8921 (N_8921,N_6575,N_7154);
and U8922 (N_8922,N_6960,N_6374);
xnor U8923 (N_8923,N_6494,N_7179);
or U8924 (N_8924,N_6200,N_6011);
nor U8925 (N_8925,N_7284,N_7079);
nor U8926 (N_8926,N_6832,N_7231);
nor U8927 (N_8927,N_7084,N_6840);
nor U8928 (N_8928,N_7493,N_7381);
nand U8929 (N_8929,N_6986,N_7095);
and U8930 (N_8930,N_6834,N_7289);
and U8931 (N_8931,N_6236,N_6973);
nor U8932 (N_8932,N_6125,N_6435);
nor U8933 (N_8933,N_7381,N_6368);
and U8934 (N_8934,N_7309,N_6481);
nand U8935 (N_8935,N_6917,N_7336);
or U8936 (N_8936,N_7366,N_6250);
and U8937 (N_8937,N_7232,N_6158);
and U8938 (N_8938,N_7128,N_6224);
nor U8939 (N_8939,N_6338,N_7362);
nor U8940 (N_8940,N_7219,N_7469);
nand U8941 (N_8941,N_6107,N_6483);
and U8942 (N_8942,N_6068,N_7476);
and U8943 (N_8943,N_6918,N_6869);
and U8944 (N_8944,N_6390,N_7279);
and U8945 (N_8945,N_6168,N_6208);
or U8946 (N_8946,N_7223,N_6824);
or U8947 (N_8947,N_7428,N_7206);
and U8948 (N_8948,N_7030,N_6922);
nand U8949 (N_8949,N_7259,N_7211);
nand U8950 (N_8950,N_7393,N_7317);
nand U8951 (N_8951,N_6580,N_6765);
or U8952 (N_8952,N_6119,N_7105);
or U8953 (N_8953,N_7341,N_6501);
xor U8954 (N_8954,N_7222,N_7411);
and U8955 (N_8955,N_6348,N_6979);
nor U8956 (N_8956,N_6466,N_6489);
and U8957 (N_8957,N_7131,N_6511);
and U8958 (N_8958,N_6802,N_6886);
nand U8959 (N_8959,N_6278,N_6268);
nor U8960 (N_8960,N_6276,N_6239);
nor U8961 (N_8961,N_6155,N_6967);
nand U8962 (N_8962,N_6940,N_7499);
nand U8963 (N_8963,N_7146,N_7299);
or U8964 (N_8964,N_6295,N_6724);
nor U8965 (N_8965,N_6073,N_6366);
nor U8966 (N_8966,N_6208,N_6726);
nor U8967 (N_8967,N_6321,N_6886);
nand U8968 (N_8968,N_7415,N_6487);
and U8969 (N_8969,N_6537,N_6966);
nor U8970 (N_8970,N_6261,N_6910);
or U8971 (N_8971,N_6659,N_6139);
nand U8972 (N_8972,N_6189,N_7390);
and U8973 (N_8973,N_6751,N_6054);
and U8974 (N_8974,N_6645,N_7238);
and U8975 (N_8975,N_6870,N_6720);
nor U8976 (N_8976,N_6825,N_6313);
and U8977 (N_8977,N_6132,N_6898);
xor U8978 (N_8978,N_6723,N_7459);
nand U8979 (N_8979,N_7412,N_6225);
and U8980 (N_8980,N_7084,N_6854);
or U8981 (N_8981,N_7199,N_7369);
nand U8982 (N_8982,N_6694,N_6123);
nor U8983 (N_8983,N_6891,N_6165);
or U8984 (N_8984,N_6974,N_6240);
nor U8985 (N_8985,N_6421,N_7216);
xor U8986 (N_8986,N_6098,N_6915);
nand U8987 (N_8987,N_6384,N_6445);
nand U8988 (N_8988,N_6348,N_6615);
nor U8989 (N_8989,N_6672,N_7459);
nand U8990 (N_8990,N_7454,N_7487);
or U8991 (N_8991,N_6781,N_6201);
and U8992 (N_8992,N_7425,N_6316);
or U8993 (N_8993,N_6079,N_6795);
and U8994 (N_8994,N_6273,N_6205);
nand U8995 (N_8995,N_6330,N_6438);
and U8996 (N_8996,N_7021,N_6183);
and U8997 (N_8997,N_7477,N_6381);
or U8998 (N_8998,N_6739,N_6834);
nand U8999 (N_8999,N_7398,N_7172);
nand U9000 (N_9000,N_8260,N_8019);
or U9001 (N_9001,N_8505,N_8738);
xor U9002 (N_9002,N_8681,N_8925);
or U9003 (N_9003,N_7743,N_8776);
xor U9004 (N_9004,N_8911,N_8364);
or U9005 (N_9005,N_8033,N_8435);
xor U9006 (N_9006,N_7756,N_8090);
and U9007 (N_9007,N_8469,N_7935);
and U9008 (N_9008,N_8450,N_8839);
nand U9009 (N_9009,N_7505,N_8516);
or U9010 (N_9010,N_8646,N_7624);
or U9011 (N_9011,N_8181,N_8695);
nand U9012 (N_9012,N_8000,N_8825);
or U9013 (N_9013,N_7778,N_8352);
xor U9014 (N_9014,N_8863,N_8936);
nor U9015 (N_9015,N_8390,N_8196);
nand U9016 (N_9016,N_8359,N_8793);
nor U9017 (N_9017,N_8787,N_7798);
nor U9018 (N_9018,N_8739,N_8576);
or U9019 (N_9019,N_7563,N_8586);
nand U9020 (N_9020,N_8676,N_7758);
or U9021 (N_9021,N_8741,N_7615);
or U9022 (N_9022,N_8256,N_7827);
xor U9023 (N_9023,N_7905,N_8305);
nor U9024 (N_9024,N_8126,N_8687);
nor U9025 (N_9025,N_7873,N_7625);
nand U9026 (N_9026,N_8963,N_7507);
and U9027 (N_9027,N_8265,N_8210);
nand U9028 (N_9028,N_7752,N_8209);
or U9029 (N_9029,N_8086,N_8229);
nor U9030 (N_9030,N_8225,N_8473);
nand U9031 (N_9031,N_8749,N_8991);
and U9032 (N_9032,N_8021,N_7828);
nand U9033 (N_9033,N_8951,N_8246);
and U9034 (N_9034,N_7973,N_8341);
nor U9035 (N_9035,N_7786,N_7989);
nor U9036 (N_9036,N_8923,N_7518);
nor U9037 (N_9037,N_8531,N_7682);
nand U9038 (N_9038,N_7939,N_8819);
and U9039 (N_9039,N_8623,N_8185);
or U9040 (N_9040,N_8812,N_8616);
xor U9041 (N_9041,N_8611,N_8729);
nor U9042 (N_9042,N_7603,N_8072);
nor U9043 (N_9043,N_7692,N_8133);
or U9044 (N_9044,N_8277,N_8891);
nor U9045 (N_9045,N_8808,N_8999);
nand U9046 (N_9046,N_7705,N_8145);
nor U9047 (N_9047,N_7753,N_8737);
nor U9048 (N_9048,N_7799,N_8029);
nor U9049 (N_9049,N_7796,N_8409);
nand U9050 (N_9050,N_7944,N_7695);
and U9051 (N_9051,N_8655,N_7814);
nand U9052 (N_9052,N_7803,N_8660);
xor U9053 (N_9053,N_8966,N_8781);
or U9054 (N_9054,N_8924,N_7820);
and U9055 (N_9055,N_8322,N_8448);
nor U9056 (N_9056,N_8498,N_8003);
and U9057 (N_9057,N_8691,N_7713);
or U9058 (N_9058,N_8226,N_7815);
and U9059 (N_9059,N_7931,N_8288);
and U9060 (N_9060,N_7593,N_8247);
nand U9061 (N_9061,N_8961,N_8700);
nand U9062 (N_9062,N_8854,N_7629);
or U9063 (N_9063,N_7754,N_8666);
nor U9064 (N_9064,N_8369,N_8249);
nor U9065 (N_9065,N_8201,N_8600);
nor U9066 (N_9066,N_8460,N_7541);
nor U9067 (N_9067,N_7678,N_7821);
and U9068 (N_9068,N_8363,N_7960);
and U9069 (N_9069,N_7703,N_8751);
nand U9070 (N_9070,N_8451,N_8091);
or U9071 (N_9071,N_8774,N_7601);
or U9072 (N_9072,N_7787,N_8767);
xor U9073 (N_9073,N_8822,N_7697);
nand U9074 (N_9074,N_8960,N_8790);
nor U9075 (N_9075,N_8765,N_7774);
nor U9076 (N_9076,N_8942,N_8922);
nor U9077 (N_9077,N_8862,N_8372);
xnor U9078 (N_9078,N_8099,N_7914);
or U9079 (N_9079,N_8235,N_8909);
nand U9080 (N_9080,N_8928,N_8568);
nor U9081 (N_9081,N_7992,N_7804);
and U9082 (N_9082,N_8647,N_7599);
nor U9083 (N_9083,N_8754,N_8710);
or U9084 (N_9084,N_7902,N_8971);
or U9085 (N_9085,N_7915,N_7959);
or U9086 (N_9086,N_7951,N_8782);
or U9087 (N_9087,N_7763,N_8335);
nor U9088 (N_9088,N_8107,N_7515);
or U9089 (N_9089,N_7958,N_7702);
nand U9090 (N_9090,N_7779,N_7894);
nor U9091 (N_9091,N_8548,N_8533);
nor U9092 (N_9092,N_8920,N_7529);
nand U9093 (N_9093,N_7592,N_7604);
or U9094 (N_9094,N_8477,N_8183);
nor U9095 (N_9095,N_8441,N_7848);
nand U9096 (N_9096,N_7572,N_7687);
and U9097 (N_9097,N_8538,N_8638);
or U9098 (N_9098,N_8397,N_8910);
xnor U9099 (N_9099,N_8306,N_7516);
nand U9100 (N_9100,N_8811,N_7963);
nand U9101 (N_9101,N_8299,N_8574);
or U9102 (N_9102,N_8261,N_8759);
and U9103 (N_9103,N_8468,N_8395);
or U9104 (N_9104,N_8817,N_8304);
nor U9105 (N_9105,N_7871,N_7974);
and U9106 (N_9106,N_7680,N_8603);
or U9107 (N_9107,N_7933,N_7907);
and U9108 (N_9108,N_7596,N_7977);
and U9109 (N_9109,N_8207,N_8258);
and U9110 (N_9110,N_7920,N_7877);
nand U9111 (N_9111,N_8431,N_8715);
and U9112 (N_9112,N_8311,N_8938);
or U9113 (N_9113,N_7860,N_7720);
nand U9114 (N_9114,N_8296,N_8972);
xnor U9115 (N_9115,N_7998,N_7547);
nor U9116 (N_9116,N_8837,N_7564);
or U9117 (N_9117,N_7940,N_8481);
and U9118 (N_9118,N_7630,N_8186);
and U9119 (N_9119,N_8279,N_8724);
and U9120 (N_9120,N_7502,N_8785);
nand U9121 (N_9121,N_8407,N_8382);
and U9122 (N_9122,N_7673,N_8705);
and U9123 (N_9123,N_8570,N_8897);
and U9124 (N_9124,N_8998,N_7932);
or U9125 (N_9125,N_8992,N_8536);
nand U9126 (N_9126,N_7688,N_7700);
or U9127 (N_9127,N_8772,N_8731);
nor U9128 (N_9128,N_7679,N_7729);
or U9129 (N_9129,N_8499,N_8973);
nand U9130 (N_9130,N_8243,N_8042);
or U9131 (N_9131,N_8561,N_7972);
nor U9132 (N_9132,N_8876,N_7837);
nand U9133 (N_9133,N_7793,N_7643);
nand U9134 (N_9134,N_7723,N_7922);
nor U9135 (N_9135,N_8177,N_8110);
and U9136 (N_9136,N_8321,N_7993);
and U9137 (N_9137,N_7842,N_8057);
or U9138 (N_9138,N_7560,N_7737);
nor U9139 (N_9139,N_8904,N_8065);
nor U9140 (N_9140,N_8262,N_7708);
and U9141 (N_9141,N_8983,N_8147);
and U9142 (N_9142,N_7947,N_8254);
and U9143 (N_9143,N_7768,N_7942);
or U9144 (N_9144,N_8712,N_8330);
nor U9145 (N_9145,N_8327,N_7988);
nand U9146 (N_9146,N_8948,N_8282);
nor U9147 (N_9147,N_7704,N_8682);
nor U9148 (N_9148,N_7943,N_8523);
nand U9149 (N_9149,N_8230,N_7900);
and U9150 (N_9150,N_8146,N_7542);
nand U9151 (N_9151,N_8708,N_7623);
nor U9152 (N_9152,N_7990,N_8613);
nor U9153 (N_9153,N_8612,N_8888);
nor U9154 (N_9154,N_8379,N_7864);
nand U9155 (N_9155,N_8138,N_8485);
or U9156 (N_9156,N_8573,N_7675);
or U9157 (N_9157,N_7612,N_7795);
and U9158 (N_9158,N_7783,N_8475);
nand U9159 (N_9159,N_8271,N_7689);
and U9160 (N_9160,N_7584,N_8281);
nand U9161 (N_9161,N_8076,N_7657);
and U9162 (N_9162,N_7818,N_8610);
or U9163 (N_9163,N_7747,N_8771);
or U9164 (N_9164,N_8530,N_7762);
or U9165 (N_9165,N_8707,N_7765);
or U9166 (N_9166,N_8667,N_8024);
or U9167 (N_9167,N_8001,N_7548);
or U9168 (N_9168,N_7903,N_8168);
or U9169 (N_9169,N_8663,N_8117);
or U9170 (N_9170,N_7714,N_8840);
and U9171 (N_9171,N_8664,N_7641);
xor U9172 (N_9172,N_7767,N_8263);
nand U9173 (N_9173,N_7773,N_7982);
nor U9174 (N_9174,N_8366,N_8040);
or U9175 (N_9175,N_8717,N_8137);
and U9176 (N_9176,N_8894,N_8870);
and U9177 (N_9177,N_7984,N_8511);
nor U9178 (N_9178,N_8711,N_8416);
nor U9179 (N_9179,N_8257,N_8845);
and U9180 (N_9180,N_7588,N_8276);
or U9181 (N_9181,N_7552,N_7709);
nand U9182 (N_9182,N_8208,N_8425);
nor U9183 (N_9183,N_7707,N_7750);
and U9184 (N_9184,N_7851,N_8496);
nand U9185 (N_9185,N_7965,N_7736);
nand U9186 (N_9186,N_8007,N_8555);
nand U9187 (N_9187,N_8240,N_8732);
nor U9188 (N_9188,N_8943,N_8786);
and U9189 (N_9189,N_8355,N_8347);
or U9190 (N_9190,N_8111,N_8908);
and U9191 (N_9191,N_8039,N_7893);
or U9192 (N_9192,N_8688,N_8527);
xnor U9193 (N_9193,N_7545,N_7841);
nor U9194 (N_9194,N_8965,N_7978);
and U9195 (N_9195,N_8976,N_8340);
or U9196 (N_9196,N_8471,N_7957);
nor U9197 (N_9197,N_8643,N_8608);
or U9198 (N_9198,N_8830,N_8482);
nor U9199 (N_9199,N_8606,N_8443);
and U9200 (N_9200,N_8761,N_7927);
or U9201 (N_9201,N_8518,N_8010);
nor U9202 (N_9202,N_8987,N_8075);
nand U9203 (N_9203,N_8402,N_8026);
or U9204 (N_9204,N_7807,N_8709);
and U9205 (N_9205,N_8859,N_7501);
nand U9206 (N_9206,N_8752,N_8385);
nand U9207 (N_9207,N_8821,N_7825);
nand U9208 (N_9208,N_8952,N_7954);
or U9209 (N_9209,N_8406,N_8978);
nand U9210 (N_9210,N_7632,N_7658);
xor U9211 (N_9211,N_8275,N_7946);
nand U9212 (N_9212,N_7976,N_8962);
and U9213 (N_9213,N_7538,N_7718);
nand U9214 (N_9214,N_8377,N_7544);
and U9215 (N_9215,N_8351,N_7757);
and U9216 (N_9216,N_7581,N_8946);
nor U9217 (N_9217,N_7797,N_8092);
and U9218 (N_9218,N_8582,N_7636);
nand U9219 (N_9219,N_8939,N_8684);
nor U9220 (N_9220,N_7967,N_7667);
and U9221 (N_9221,N_8805,N_8017);
and U9222 (N_9222,N_7923,N_8045);
xnor U9223 (N_9223,N_8634,N_8081);
or U9224 (N_9224,N_7832,N_8062);
and U9225 (N_9225,N_8134,N_7732);
nand U9226 (N_9226,N_8728,N_8216);
xnor U9227 (N_9227,N_8599,N_8622);
and U9228 (N_9228,N_8926,N_7626);
nor U9229 (N_9229,N_8101,N_8456);
or U9230 (N_9230,N_8480,N_7906);
and U9231 (N_9231,N_7761,N_7878);
nor U9232 (N_9232,N_8993,N_8047);
or U9233 (N_9233,N_7513,N_7634);
nor U9234 (N_9234,N_8815,N_8627);
nor U9235 (N_9235,N_8083,N_7857);
or U9236 (N_9236,N_7840,N_8342);
or U9237 (N_9237,N_8562,N_8144);
or U9238 (N_9238,N_8766,N_7606);
nor U9239 (N_9239,N_8585,N_7711);
and U9240 (N_9240,N_7845,N_8565);
nand U9241 (N_9241,N_7831,N_8637);
and U9242 (N_9242,N_8266,N_8064);
or U9243 (N_9243,N_7770,N_8620);
and U9244 (N_9244,N_8604,N_8847);
and U9245 (N_9245,N_8584,N_8806);
nor U9246 (N_9246,N_7554,N_8872);
or U9247 (N_9247,N_7605,N_8002);
xnor U9248 (N_9248,N_8566,N_8319);
or U9249 (N_9249,N_7670,N_7671);
or U9250 (N_9250,N_7609,N_7503);
nor U9251 (N_9251,N_8726,N_8470);
nor U9252 (N_9252,N_7706,N_7537);
or U9253 (N_9253,N_8861,N_7504);
and U9254 (N_9254,N_7867,N_7861);
or U9255 (N_9255,N_7874,N_7610);
and U9256 (N_9256,N_7622,N_8095);
and U9257 (N_9257,N_8412,N_8866);
nor U9258 (N_9258,N_7510,N_8896);
or U9259 (N_9259,N_8336,N_7668);
nand U9260 (N_9260,N_8802,N_8697);
nand U9261 (N_9261,N_8339,N_8238);
and U9262 (N_9262,N_7508,N_8621);
nor U9263 (N_9263,N_7512,N_8769);
nand U9264 (N_9264,N_7574,N_8334);
nand U9265 (N_9265,N_8832,N_8905);
and U9266 (N_9266,N_8102,N_8510);
and U9267 (N_9267,N_8014,N_8673);
and U9268 (N_9268,N_8831,N_8857);
and U9269 (N_9269,N_8295,N_8828);
and U9270 (N_9270,N_8778,N_8730);
and U9271 (N_9271,N_8959,N_7628);
nor U9272 (N_9272,N_8968,N_7777);
or U9273 (N_9273,N_8479,N_8085);
and U9274 (N_9274,N_7859,N_8239);
nor U9275 (N_9275,N_7524,N_8096);
or U9276 (N_9276,N_7566,N_7698);
nor U9277 (N_9277,N_8362,N_7608);
nor U9278 (N_9278,N_8692,N_8388);
nor U9279 (N_9279,N_8956,N_8423);
nor U9280 (N_9280,N_8411,N_7971);
or U9281 (N_9281,N_7746,N_8344);
nand U9282 (N_9282,N_8494,N_7968);
or U9283 (N_9283,N_8829,N_8596);
nor U9284 (N_9284,N_8841,N_7808);
nor U9285 (N_9285,N_7633,N_7745);
xor U9286 (N_9286,N_8259,N_7567);
nor U9287 (N_9287,N_7600,N_7966);
and U9288 (N_9288,N_8994,N_8320);
nand U9289 (N_9289,N_8650,N_8124);
and U9290 (N_9290,N_7721,N_8457);
nand U9291 (N_9291,N_8540,N_7526);
or U9292 (N_9292,N_7728,N_7997);
or U9293 (N_9293,N_8253,N_8383);
nand U9294 (N_9294,N_8036,N_8777);
nor U9295 (N_9295,N_8656,N_7817);
nor U9296 (N_9296,N_7776,N_7514);
nand U9297 (N_9297,N_8106,N_8583);
nand U9298 (N_9298,N_7500,N_8486);
and U9299 (N_9299,N_8345,N_7986);
nand U9300 (N_9300,N_8580,N_8399);
nand U9301 (N_9301,N_8324,N_8602);
xor U9302 (N_9302,N_8720,N_7693);
nor U9303 (N_9303,N_7550,N_7562);
or U9304 (N_9304,N_8293,N_8489);
xnor U9305 (N_9305,N_7930,N_8686);
nor U9306 (N_9306,N_8192,N_7956);
and U9307 (N_9307,N_8524,N_8696);
and U9308 (N_9308,N_8337,N_8278);
or U9309 (N_9309,N_8454,N_8300);
and U9310 (N_9310,N_8661,N_8179);
nor U9311 (N_9311,N_7525,N_7666);
or U9312 (N_9312,N_8043,N_7573);
and U9313 (N_9313,N_8375,N_8316);
and U9314 (N_9314,N_8917,N_8556);
and U9315 (N_9315,N_8414,N_8898);
nand U9316 (N_9316,N_7784,N_8564);
and U9317 (N_9317,N_8329,N_7921);
and U9318 (N_9318,N_8970,N_7901);
nand U9319 (N_9319,N_8690,N_8374);
nor U9320 (N_9320,N_8025,N_8312);
and U9321 (N_9321,N_8105,N_7645);
nand U9322 (N_9322,N_8784,N_7888);
nand U9323 (N_9323,N_7892,N_8463);
nor U9324 (N_9324,N_7647,N_8109);
and U9325 (N_9325,N_7897,N_8503);
nor U9326 (N_9326,N_8255,N_8947);
and U9327 (N_9327,N_8141,N_8877);
or U9328 (N_9328,N_8698,N_7568);
xnor U9329 (N_9329,N_7809,N_8733);
nand U9330 (N_9330,N_8988,N_7898);
and U9331 (N_9331,N_8071,N_8795);
nor U9332 (N_9332,N_8796,N_8171);
and U9333 (N_9333,N_8858,N_8685);
nor U9334 (N_9334,N_8886,N_8537);
nor U9335 (N_9335,N_8895,N_7913);
xnor U9336 (N_9336,N_7816,N_7724);
and U9337 (N_9337,N_8162,N_8572);
or U9338 (N_9338,N_8442,N_7640);
nand U9339 (N_9339,N_7543,N_7755);
nand U9340 (N_9340,N_8885,N_8308);
or U9341 (N_9341,N_8515,N_7691);
xor U9342 (N_9342,N_8860,N_8597);
nor U9343 (N_9343,N_8955,N_8982);
and U9344 (N_9344,N_8031,N_7621);
nor U9345 (N_9345,N_7686,N_7889);
nor U9346 (N_9346,N_8581,N_8497);
or U9347 (N_9347,N_7551,N_8267);
or U9348 (N_9348,N_8615,N_8069);
or U9349 (N_9349,N_7590,N_8929);
and U9350 (N_9350,N_8674,N_8338);
nor U9351 (N_9351,N_7996,N_8020);
nor U9352 (N_9352,N_8689,N_7852);
xor U9353 (N_9353,N_8163,N_7938);
nor U9354 (N_9354,N_8986,N_8325);
nand U9355 (N_9355,N_8763,N_8918);
xnor U9356 (N_9356,N_8549,N_7523);
and U9357 (N_9357,N_7883,N_8804);
nand U9358 (N_9358,N_7530,N_7683);
nand U9359 (N_9359,N_8871,N_8504);
and U9360 (N_9360,N_8426,N_8360);
xnor U9361 (N_9361,N_8838,N_7659);
xor U9362 (N_9362,N_7789,N_8120);
nand U9363 (N_9363,N_8501,N_8487);
and U9364 (N_9364,N_8723,N_8170);
nand U9365 (N_9365,N_7533,N_8438);
xnor U9366 (N_9366,N_8328,N_8849);
and U9367 (N_9367,N_8315,N_8493);
and U9368 (N_9368,N_8157,N_7904);
nor U9369 (N_9369,N_8964,N_8571);
xor U9370 (N_9370,N_7655,N_8892);
xor U9371 (N_9371,N_8213,N_7571);
and U9372 (N_9372,N_7646,N_7911);
nand U9373 (N_9373,N_8483,N_8748);
nand U9374 (N_9374,N_8151,N_7811);
nand U9375 (N_9375,N_8507,N_7881);
or U9376 (N_9376,N_7969,N_8403);
nand U9377 (N_9377,N_8419,N_8089);
nand U9378 (N_9378,N_8757,N_7802);
and U9379 (N_9379,N_7854,N_8143);
or U9380 (N_9380,N_7865,N_7654);
nand U9381 (N_9381,N_7690,N_8104);
or U9382 (N_9382,N_8444,N_8668);
and U9383 (N_9383,N_8750,N_8669);
nor U9384 (N_9384,N_8553,N_8373);
or U9385 (N_9385,N_8657,N_8756);
or U9386 (N_9386,N_8394,N_8234);
nor U9387 (N_9387,N_8810,N_8464);
nand U9388 (N_9388,N_8123,N_7810);
xnor U9389 (N_9389,N_7649,N_7651);
or U9390 (N_9390,N_8902,N_8048);
nor U9391 (N_9391,N_8066,N_8563);
nand U9392 (N_9392,N_8368,N_7598);
or U9393 (N_9393,N_8792,N_8678);
and U9394 (N_9394,N_8365,N_8220);
xor U9395 (N_9395,N_8940,N_8636);
and U9396 (N_9396,N_7672,N_8618);
or U9397 (N_9397,N_8607,N_8309);
nor U9398 (N_9398,N_8990,N_7511);
or U9399 (N_9399,N_8714,N_8557);
and U9400 (N_9400,N_8915,N_7800);
nor U9401 (N_9401,N_8827,N_8227);
nor U9402 (N_9402,N_8197,N_8156);
nand U9403 (N_9403,N_7918,N_8791);
and U9404 (N_9404,N_7521,N_8430);
or U9405 (N_9405,N_7839,N_7909);
nor U9406 (N_9406,N_8848,N_8881);
nand U9407 (N_9407,N_8508,N_8914);
and U9408 (N_9408,N_8153,N_8041);
nand U9409 (N_9409,N_7639,N_7715);
or U9410 (N_9410,N_8758,N_8051);
nor U9411 (N_9411,N_7937,N_8193);
and U9412 (N_9412,N_8052,N_7980);
and U9413 (N_9413,N_8250,N_8798);
nand U9414 (N_9414,N_8060,N_7587);
nor U9415 (N_9415,N_8176,N_8058);
nand U9416 (N_9416,N_7764,N_8880);
or U9417 (N_9417,N_7570,N_8842);
nor U9418 (N_9418,N_8073,N_8114);
nand U9419 (N_9419,N_8921,N_8624);
or U9420 (N_9420,N_8658,N_7549);
nor U9421 (N_9421,N_8059,N_8474);
and U9422 (N_9422,N_7858,N_8601);
or U9423 (N_9423,N_8651,N_7785);
and U9424 (N_9424,N_8298,N_8850);
or U9425 (N_9425,N_7577,N_8514);
nor U9426 (N_9426,N_8617,N_8670);
nor U9427 (N_9427,N_7701,N_8165);
nand U9428 (N_9428,N_8544,N_8466);
or U9429 (N_9429,N_8361,N_8941);
or U9430 (N_9430,N_7546,N_8354);
nand U9431 (N_9431,N_8814,N_8834);
nand U9432 (N_9432,N_8706,N_8011);
or U9433 (N_9433,N_8937,N_7970);
nor U9434 (N_9434,N_8386,N_8116);
nor U9435 (N_9435,N_8252,N_8461);
nand U9436 (N_9436,N_7635,N_8317);
and U9437 (N_9437,N_7579,N_8135);
and U9438 (N_9438,N_7813,N_8653);
nand U9439 (N_9439,N_8716,N_7561);
xnor U9440 (N_9440,N_8182,N_8439);
xnor U9441 (N_9441,N_8422,N_8526);
and U9442 (N_9442,N_8376,N_8727);
nand U9443 (N_9443,N_8996,N_7620);
and U9444 (N_9444,N_7602,N_7586);
and U9445 (N_9445,N_7739,N_8434);
nor U9446 (N_9446,N_8520,N_7744);
and U9447 (N_9447,N_8878,N_7677);
and U9448 (N_9448,N_7528,N_8313);
nand U9449 (N_9449,N_7642,N_7652);
or U9450 (N_9450,N_8626,N_7945);
nor U9451 (N_9451,N_7519,N_7725);
nor U9452 (N_9452,N_7589,N_7834);
and U9453 (N_9453,N_7847,N_7637);
and U9454 (N_9454,N_8191,N_8077);
or U9455 (N_9455,N_8773,N_8559);
nor U9456 (N_9456,N_7722,N_8635);
nand U9457 (N_9457,N_8142,N_7981);
nand U9458 (N_9458,N_8242,N_8558);
nand U9459 (N_9459,N_8541,N_8890);
nor U9460 (N_9460,N_8949,N_7955);
or U9461 (N_9461,N_8935,N_8084);
nand U9462 (N_9462,N_8887,N_8893);
nand U9463 (N_9463,N_8189,N_7539);
and U9464 (N_9464,N_8542,N_7506);
or U9465 (N_9465,N_8067,N_8953);
nor U9466 (N_9466,N_8108,N_8833);
xnor U9467 (N_9467,N_8579,N_8428);
xnor U9468 (N_9468,N_8211,N_8818);
nand U9469 (N_9469,N_8172,N_8053);
and U9470 (N_9470,N_7522,N_7788);
or U9471 (N_9471,N_7853,N_8215);
xnor U9472 (N_9472,N_7726,N_8136);
or U9473 (N_9473,N_8588,N_7880);
or U9474 (N_9474,N_8224,N_8703);
or U9475 (N_9475,N_8005,N_7648);
nor U9476 (N_9476,N_8453,N_8056);
or U9477 (N_9477,N_8868,N_7638);
xnor U9478 (N_9478,N_8662,N_8578);
nand U9479 (N_9479,N_8916,N_8346);
and U9480 (N_9480,N_8743,N_8869);
nor U9481 (N_9481,N_7850,N_7712);
nand U9482 (N_9482,N_8121,N_8264);
nor U9483 (N_9483,N_8035,N_7771);
xor U9484 (N_9484,N_8004,N_8699);
nor U9485 (N_9485,N_8356,N_8413);
nand U9486 (N_9486,N_8645,N_8221);
and U9487 (N_9487,N_7616,N_8274);
nand U9488 (N_9488,N_8855,N_8467);
nand U9489 (N_9489,N_8502,N_7532);
or U9490 (N_9490,N_7742,N_7890);
nor U9491 (N_9491,N_8797,N_8476);
or U9492 (N_9492,N_8150,N_8323);
and U9493 (N_9493,N_8899,N_8619);
and U9494 (N_9494,N_8694,N_8721);
and U9495 (N_9495,N_8852,N_7917);
xnor U9496 (N_9496,N_7936,N_8205);
or U9497 (N_9497,N_7509,N_8314);
nand U9498 (N_9498,N_8985,N_7979);
or U9499 (N_9499,N_8237,N_8012);
nand U9500 (N_9500,N_8418,N_7597);
nand U9501 (N_9501,N_8396,N_8560);
or U9502 (N_9502,N_8753,N_8631);
nor U9503 (N_9503,N_8659,N_8028);
nor U9504 (N_9504,N_8800,N_8592);
or U9505 (N_9505,N_8843,N_8233);
nor U9506 (N_9506,N_8577,N_8100);
or U9507 (N_9507,N_7925,N_8044);
xnor U9508 (N_9508,N_8648,N_8358);
nor U9509 (N_9509,N_8975,N_8977);
and U9510 (N_9510,N_8050,N_8302);
nand U9511 (N_9511,N_8519,N_7835);
nand U9512 (N_9512,N_8589,N_8155);
xnor U9513 (N_9513,N_7740,N_8149);
nand U9514 (N_9514,N_8310,N_8630);
or U9515 (N_9515,N_8160,N_7676);
nor U9516 (N_9516,N_8292,N_8129);
or U9517 (N_9517,N_8174,N_8068);
and U9518 (N_9518,N_8140,N_7520);
and U9519 (N_9519,N_7812,N_8780);
nand U9520 (N_9520,N_8979,N_8984);
or U9521 (N_9521,N_7849,N_8639);
nand U9522 (N_9522,N_8521,N_7607);
or U9523 (N_9523,N_8649,N_8289);
or U9524 (N_9524,N_7836,N_8879);
and U9525 (N_9525,N_7727,N_7833);
nand U9526 (N_9526,N_8823,N_7948);
or U9527 (N_9527,N_8115,N_7760);
nand U9528 (N_9528,N_8594,N_8417);
xor U9529 (N_9529,N_7733,N_8332);
and U9530 (N_9530,N_8190,N_8022);
nand U9531 (N_9531,N_7791,N_7595);
nand U9532 (N_9532,N_7619,N_8273);
nor U9533 (N_9533,N_7631,N_8906);
or U9534 (N_9534,N_8932,N_7844);
nor U9535 (N_9535,N_7822,N_8628);
or U9536 (N_9536,N_8683,N_8718);
and U9537 (N_9537,N_8127,N_8410);
nand U9538 (N_9538,N_8184,N_8595);
and U9539 (N_9539,N_8957,N_7819);
and U9540 (N_9540,N_8164,N_8472);
or U9541 (N_9541,N_8934,N_7866);
nand U9542 (N_9542,N_8128,N_7716);
nand U9543 (N_9543,N_7887,N_8462);
and U9544 (N_9544,N_8532,N_8447);
and U9545 (N_9545,N_8919,N_7962);
nand U9546 (N_9546,N_7749,N_8343);
or U9547 (N_9547,N_8125,N_7627);
and U9548 (N_9548,N_7801,N_8291);
nor U9549 (N_9549,N_7856,N_8495);
or U9550 (N_9550,N_7995,N_8546);
xor U9551 (N_9551,N_8794,N_8404);
xnor U9552 (N_9552,N_7926,N_8551);
or U9553 (N_9553,N_8903,N_7964);
or U9554 (N_9554,N_8865,N_8175);
or U9555 (N_9555,N_8452,N_7794);
and U9556 (N_9556,N_7994,N_8445);
xnor U9557 (N_9557,N_8799,N_8113);
xnor U9558 (N_9558,N_8119,N_7661);
nor U9559 (N_9559,N_7838,N_8006);
nor U9560 (N_9560,N_8132,N_8736);
nor U9561 (N_9561,N_8567,N_8398);
nor U9562 (N_9562,N_7910,N_7983);
nand U9563 (N_9563,N_7879,N_7660);
nor U9564 (N_9564,N_8082,N_7806);
or U9565 (N_9565,N_8640,N_7941);
and U9566 (N_9566,N_8206,N_8768);
nand U9567 (N_9567,N_8008,N_8517);
nor U9568 (N_9568,N_8764,N_8642);
and U9569 (N_9569,N_8875,N_8954);
nor U9570 (N_9570,N_7823,N_8384);
nor U9571 (N_9571,N_8693,N_8590);
or U9572 (N_9572,N_8874,N_8251);
and U9573 (N_9573,N_8037,N_7751);
or U9574 (N_9574,N_8883,N_7517);
and U9575 (N_9575,N_8535,N_7665);
or U9576 (N_9576,N_8087,N_8844);
nor U9577 (N_9577,N_7775,N_7576);
and U9578 (N_9578,N_8195,N_8745);
xor U9579 (N_9579,N_8188,N_7559);
nand U9580 (N_9580,N_8746,N_7719);
nor U9581 (N_9581,N_8747,N_7830);
and U9582 (N_9582,N_8629,N_8930);
or U9583 (N_9583,N_7614,N_7580);
nor U9584 (N_9584,N_7540,N_8492);
xnor U9585 (N_9585,N_7759,N_7862);
nor U9586 (N_9586,N_8178,N_7681);
or U9587 (N_9587,N_8199,N_8459);
nor U9588 (N_9588,N_8389,N_8803);
xnor U9589 (N_9589,N_7985,N_8200);
nand U9590 (N_9590,N_8488,N_8927);
nand U9591 (N_9591,N_8401,N_8826);
xnor U9592 (N_9592,N_8490,N_8248);
and U9593 (N_9593,N_8704,N_8370);
and U9594 (N_9594,N_8809,N_8813);
nand U9595 (N_9595,N_8788,N_8884);
nor U9596 (N_9596,N_8427,N_8569);
and U9597 (N_9597,N_8440,N_8734);
nand U9598 (N_9598,N_8286,N_8824);
and U9599 (N_9599,N_7578,N_8228);
nand U9600 (N_9600,N_8236,N_8166);
or U9601 (N_9601,N_7805,N_8380);
or U9602 (N_9602,N_7782,N_8770);
nand U9603 (N_9603,N_8078,N_8679);
nand U9604 (N_9604,N_7829,N_8097);
or U9605 (N_9605,N_7896,N_7908);
and U9606 (N_9606,N_8755,N_8093);
nor U9607 (N_9607,N_7694,N_7569);
or U9608 (N_9608,N_8283,N_8198);
xnor U9609 (N_9609,N_7975,N_7899);
nand U9610 (N_9610,N_8722,N_8644);
xnor U9611 (N_9611,N_8027,N_8701);
nand U9612 (N_9612,N_8013,N_8491);
or U9613 (N_9613,N_7891,N_8307);
or U9614 (N_9614,N_8677,N_8539);
nor U9615 (N_9615,N_7991,N_7895);
or U9616 (N_9616,N_8326,N_8543);
nand U9617 (N_9617,N_8900,N_8901);
nor U9618 (N_9618,N_8522,N_7558);
nand U9619 (N_9619,N_8015,N_7780);
nand U9620 (N_9620,N_8974,N_8154);
nor U9621 (N_9621,N_8446,N_8484);
or U9622 (N_9622,N_8882,N_7882);
nand U9623 (N_9623,N_8270,N_7582);
nor U9624 (N_9624,N_7662,N_7617);
and U9625 (N_9625,N_8458,N_8873);
nand U9626 (N_9626,N_8867,N_8223);
and U9627 (N_9627,N_8614,N_8161);
and U9628 (N_9628,N_8836,N_8725);
nand U9629 (N_9629,N_7912,N_8641);
or U9630 (N_9630,N_8944,N_8118);
nor U9631 (N_9631,N_7674,N_8420);
nor U9632 (N_9632,N_8222,N_8214);
nor U9633 (N_9633,N_8632,N_8074);
nand U9634 (N_9634,N_7884,N_8500);
nor U9635 (N_9635,N_8030,N_8913);
or U9636 (N_9636,N_7790,N_8719);
nor U9637 (N_9637,N_8393,N_8285);
nor U9638 (N_9638,N_8512,N_7781);
or U9639 (N_9639,N_8625,N_8244);
xor U9640 (N_9640,N_7929,N_8598);
or U9641 (N_9641,N_8449,N_8587);
nor U9642 (N_9642,N_8112,N_8680);
or U9643 (N_9643,N_8169,N_8268);
and U9644 (N_9644,N_8212,N_8835);
or U9645 (N_9645,N_8152,N_8204);
xor U9646 (N_9646,N_8301,N_8070);
nor U9647 (N_9647,N_8981,N_8421);
and U9648 (N_9648,N_8232,N_7734);
nand U9649 (N_9649,N_7876,N_8187);
nor U9650 (N_9650,N_7536,N_7594);
and U9651 (N_9651,N_8591,N_8016);
nor U9652 (N_9652,N_8672,N_8465);
nand U9653 (N_9653,N_8436,N_7869);
nor U9654 (N_9654,N_8742,N_7650);
xor U9655 (N_9655,N_8593,N_8034);
or U9656 (N_9656,N_8429,N_8049);
nand U9657 (N_9657,N_7999,N_8094);
or U9658 (N_9658,N_8801,N_8202);
or U9659 (N_9659,N_7928,N_8353);
nor U9660 (N_9660,N_8912,N_8378);
nand U9661 (N_9661,N_7557,N_8529);
nand U9662 (N_9662,N_7613,N_7949);
or U9663 (N_9663,N_7685,N_7710);
or U9664 (N_9664,N_8272,N_8654);
and U9665 (N_9665,N_8061,N_7855);
xnor U9666 (N_9666,N_7611,N_7919);
nor U9667 (N_9667,N_7953,N_8424);
nor U9668 (N_9668,N_8303,N_7669);
xor U9669 (N_9669,N_7824,N_8455);
or U9670 (N_9670,N_8851,N_8297);
or U9671 (N_9671,N_8605,N_8241);
nor U9672 (N_9672,N_8367,N_7717);
nor U9673 (N_9673,N_7885,N_8405);
nand U9674 (N_9674,N_7735,N_8381);
or U9675 (N_9675,N_7738,N_7699);
or U9676 (N_9676,N_8290,N_8408);
or U9677 (N_9677,N_8775,N_8575);
nand U9678 (N_9678,N_8506,N_8392);
or U9679 (N_9679,N_8387,N_8180);
nand U9680 (N_9680,N_8098,N_7870);
and U9681 (N_9681,N_8009,N_8552);
nand U9682 (N_9682,N_8652,N_8995);
and U9683 (N_9683,N_8167,N_8760);
and U9684 (N_9684,N_8931,N_7553);
and U9685 (N_9685,N_8148,N_7527);
or U9686 (N_9686,N_8294,N_8853);
nor U9687 (N_9687,N_8534,N_7843);
nand U9688 (N_9688,N_7924,N_7731);
nor U9689 (N_9689,N_7585,N_7916);
or U9690 (N_9690,N_8046,N_8945);
nor U9691 (N_9691,N_7696,N_8054);
nand U9692 (N_9692,N_8789,N_8528);
or U9693 (N_9693,N_8554,N_8967);
or U9694 (N_9694,N_8864,N_7766);
nand U9695 (N_9695,N_8779,N_8219);
or U9696 (N_9696,N_8744,N_7950);
nand U9697 (N_9697,N_8702,N_8609);
and U9698 (N_9698,N_7575,N_8350);
and U9699 (N_9699,N_8269,N_7846);
nand U9700 (N_9700,N_8371,N_8063);
nor U9701 (N_9701,N_8997,N_7535);
or U9702 (N_9702,N_7664,N_8103);
or U9703 (N_9703,N_8348,N_8023);
and U9704 (N_9704,N_8131,N_8122);
and U9705 (N_9705,N_8284,N_8231);
nor U9706 (N_9706,N_8203,N_8547);
or U9707 (N_9707,N_8550,N_8762);
and U9708 (N_9708,N_7591,N_8509);
nor U9709 (N_9709,N_7663,N_8950);
nand U9710 (N_9710,N_8080,N_8437);
nand U9711 (N_9711,N_8318,N_8989);
nand U9712 (N_9712,N_8173,N_8331);
nor U9713 (N_9713,N_7644,N_7875);
nand U9714 (N_9714,N_8139,N_8735);
and U9715 (N_9715,N_8513,N_7872);
or U9716 (N_9716,N_8055,N_8159);
nand U9717 (N_9717,N_7556,N_8969);
nand U9718 (N_9718,N_8889,N_7555);
xnor U9719 (N_9719,N_8933,N_8713);
and U9720 (N_9720,N_8194,N_8958);
or U9721 (N_9721,N_8783,N_8130);
or U9722 (N_9722,N_7583,N_8018);
nor U9723 (N_9723,N_7748,N_7792);
xor U9724 (N_9724,N_7684,N_8740);
nand U9725 (N_9725,N_7531,N_7730);
and U9726 (N_9726,N_7961,N_8633);
nor U9727 (N_9727,N_8432,N_8820);
nand U9728 (N_9728,N_8088,N_8217);
or U9729 (N_9729,N_8545,N_7565);
and U9730 (N_9730,N_8816,N_8280);
or U9731 (N_9731,N_7741,N_8907);
or U9732 (N_9732,N_7656,N_7769);
nand U9733 (N_9733,N_7952,N_8287);
and U9734 (N_9734,N_8846,N_7886);
and U9735 (N_9735,N_7618,N_8333);
or U9736 (N_9736,N_8357,N_7826);
or U9737 (N_9737,N_8218,N_7772);
nor U9738 (N_9738,N_8807,N_8415);
or U9739 (N_9739,N_8671,N_8675);
nor U9740 (N_9740,N_7534,N_8245);
or U9741 (N_9741,N_8525,N_8433);
xnor U9742 (N_9742,N_8158,N_7863);
or U9743 (N_9743,N_8391,N_7934);
and U9744 (N_9744,N_7653,N_7868);
and U9745 (N_9745,N_8038,N_8079);
or U9746 (N_9746,N_8478,N_8856);
nor U9747 (N_9747,N_7987,N_8400);
nor U9748 (N_9748,N_8980,N_8032);
nand U9749 (N_9749,N_8349,N_8665);
nor U9750 (N_9750,N_8140,N_8254);
and U9751 (N_9751,N_7857,N_8468);
xnor U9752 (N_9752,N_8801,N_8391);
and U9753 (N_9753,N_8424,N_8675);
nand U9754 (N_9754,N_7970,N_7639);
nand U9755 (N_9755,N_8700,N_8400);
or U9756 (N_9756,N_8441,N_8432);
or U9757 (N_9757,N_8747,N_8123);
and U9758 (N_9758,N_8983,N_7865);
nor U9759 (N_9759,N_8694,N_7613);
nor U9760 (N_9760,N_8363,N_8289);
and U9761 (N_9761,N_8769,N_8947);
nand U9762 (N_9762,N_8781,N_7714);
nor U9763 (N_9763,N_7555,N_8305);
or U9764 (N_9764,N_8596,N_8170);
or U9765 (N_9765,N_8042,N_7501);
nor U9766 (N_9766,N_8018,N_8747);
or U9767 (N_9767,N_8810,N_8723);
nor U9768 (N_9768,N_8777,N_8846);
nand U9769 (N_9769,N_8454,N_7975);
nand U9770 (N_9770,N_8086,N_8289);
and U9771 (N_9771,N_8597,N_8343);
or U9772 (N_9772,N_8195,N_8412);
and U9773 (N_9773,N_7584,N_8383);
or U9774 (N_9774,N_7540,N_8112);
and U9775 (N_9775,N_8659,N_8478);
nor U9776 (N_9776,N_8801,N_8881);
or U9777 (N_9777,N_7703,N_7668);
nand U9778 (N_9778,N_8058,N_8095);
nor U9779 (N_9779,N_7595,N_8019);
nor U9780 (N_9780,N_8345,N_8453);
or U9781 (N_9781,N_7617,N_8662);
and U9782 (N_9782,N_8472,N_8639);
nor U9783 (N_9783,N_8926,N_7658);
nand U9784 (N_9784,N_7834,N_8552);
or U9785 (N_9785,N_7844,N_8584);
or U9786 (N_9786,N_8806,N_7779);
or U9787 (N_9787,N_7930,N_8433);
and U9788 (N_9788,N_8465,N_8956);
nor U9789 (N_9789,N_8534,N_8825);
nor U9790 (N_9790,N_8945,N_8310);
nand U9791 (N_9791,N_7547,N_7535);
nand U9792 (N_9792,N_7870,N_7667);
nor U9793 (N_9793,N_7911,N_7614);
nor U9794 (N_9794,N_7677,N_8913);
xor U9795 (N_9795,N_8968,N_8317);
or U9796 (N_9796,N_7603,N_8918);
or U9797 (N_9797,N_7785,N_8789);
or U9798 (N_9798,N_8612,N_8414);
nand U9799 (N_9799,N_8718,N_8798);
nor U9800 (N_9800,N_7763,N_8830);
nor U9801 (N_9801,N_8266,N_8416);
and U9802 (N_9802,N_8778,N_8417);
and U9803 (N_9803,N_8428,N_7646);
nand U9804 (N_9804,N_8061,N_7736);
and U9805 (N_9805,N_8742,N_8084);
nor U9806 (N_9806,N_7911,N_7525);
xnor U9807 (N_9807,N_7714,N_8580);
xnor U9808 (N_9808,N_7948,N_8656);
and U9809 (N_9809,N_8909,N_7765);
nor U9810 (N_9810,N_8226,N_7968);
nor U9811 (N_9811,N_8580,N_8699);
xor U9812 (N_9812,N_8222,N_8499);
or U9813 (N_9813,N_8263,N_7553);
nand U9814 (N_9814,N_8856,N_7793);
nand U9815 (N_9815,N_7648,N_7701);
and U9816 (N_9816,N_7969,N_8647);
or U9817 (N_9817,N_8286,N_8042);
and U9818 (N_9818,N_8898,N_8815);
nand U9819 (N_9819,N_8570,N_8902);
nand U9820 (N_9820,N_8958,N_7809);
nand U9821 (N_9821,N_8162,N_8013);
and U9822 (N_9822,N_8710,N_8491);
nand U9823 (N_9823,N_8280,N_8795);
or U9824 (N_9824,N_8077,N_8581);
xnor U9825 (N_9825,N_8752,N_8365);
and U9826 (N_9826,N_8720,N_8617);
xnor U9827 (N_9827,N_7511,N_8928);
or U9828 (N_9828,N_8200,N_8508);
nand U9829 (N_9829,N_8551,N_8951);
nand U9830 (N_9830,N_8316,N_8614);
nor U9831 (N_9831,N_7673,N_8458);
or U9832 (N_9832,N_7905,N_8919);
xnor U9833 (N_9833,N_8312,N_8303);
nor U9834 (N_9834,N_8281,N_8067);
or U9835 (N_9835,N_7567,N_8587);
nor U9836 (N_9836,N_8051,N_8762);
nand U9837 (N_9837,N_8666,N_8064);
nor U9838 (N_9838,N_8593,N_7518);
and U9839 (N_9839,N_7710,N_8712);
nand U9840 (N_9840,N_8152,N_8256);
and U9841 (N_9841,N_7669,N_8439);
nand U9842 (N_9842,N_8171,N_8319);
or U9843 (N_9843,N_8038,N_8134);
nor U9844 (N_9844,N_7995,N_8579);
or U9845 (N_9845,N_7937,N_7823);
xnor U9846 (N_9846,N_8718,N_8100);
or U9847 (N_9847,N_8012,N_8677);
nor U9848 (N_9848,N_7707,N_7907);
and U9849 (N_9849,N_8553,N_8041);
and U9850 (N_9850,N_8992,N_8901);
and U9851 (N_9851,N_8558,N_8485);
nand U9852 (N_9852,N_8274,N_8013);
and U9853 (N_9853,N_8126,N_7614);
or U9854 (N_9854,N_8750,N_8096);
nand U9855 (N_9855,N_8074,N_8795);
nor U9856 (N_9856,N_8207,N_8383);
and U9857 (N_9857,N_8722,N_8741);
nor U9858 (N_9858,N_8571,N_7804);
nand U9859 (N_9859,N_8272,N_7584);
or U9860 (N_9860,N_8021,N_8677);
nand U9861 (N_9861,N_8266,N_7679);
and U9862 (N_9862,N_7521,N_8806);
or U9863 (N_9863,N_8364,N_8788);
and U9864 (N_9864,N_8450,N_7620);
nand U9865 (N_9865,N_8973,N_8991);
nand U9866 (N_9866,N_8921,N_8504);
nand U9867 (N_9867,N_8534,N_8588);
and U9868 (N_9868,N_8181,N_8142);
nor U9869 (N_9869,N_8550,N_7820);
and U9870 (N_9870,N_8857,N_8641);
nand U9871 (N_9871,N_7639,N_7534);
nor U9872 (N_9872,N_8202,N_8527);
or U9873 (N_9873,N_7788,N_8993);
or U9874 (N_9874,N_7965,N_8277);
nor U9875 (N_9875,N_8316,N_8286);
or U9876 (N_9876,N_8528,N_8919);
nor U9877 (N_9877,N_7556,N_8263);
nor U9878 (N_9878,N_8882,N_7906);
and U9879 (N_9879,N_8449,N_8429);
nor U9880 (N_9880,N_7837,N_8049);
and U9881 (N_9881,N_7740,N_8233);
nor U9882 (N_9882,N_8852,N_8644);
or U9883 (N_9883,N_8115,N_8634);
and U9884 (N_9884,N_8329,N_8916);
and U9885 (N_9885,N_8054,N_8233);
nand U9886 (N_9886,N_8001,N_7655);
nor U9887 (N_9887,N_8372,N_8421);
nor U9888 (N_9888,N_7871,N_7959);
nand U9889 (N_9889,N_7725,N_8814);
nand U9890 (N_9890,N_8863,N_8325);
nor U9891 (N_9891,N_8210,N_7656);
xnor U9892 (N_9892,N_7896,N_8961);
nor U9893 (N_9893,N_8185,N_8621);
xnor U9894 (N_9894,N_7984,N_8040);
or U9895 (N_9895,N_8774,N_8483);
and U9896 (N_9896,N_8036,N_8154);
xor U9897 (N_9897,N_8441,N_7509);
nand U9898 (N_9898,N_8735,N_7727);
or U9899 (N_9899,N_7726,N_7632);
nor U9900 (N_9900,N_7896,N_8405);
nor U9901 (N_9901,N_8075,N_8019);
or U9902 (N_9902,N_8783,N_8733);
and U9903 (N_9903,N_8765,N_7828);
xnor U9904 (N_9904,N_7796,N_7631);
and U9905 (N_9905,N_8849,N_8979);
or U9906 (N_9906,N_8066,N_8948);
nand U9907 (N_9907,N_8595,N_7665);
and U9908 (N_9908,N_8289,N_8189);
and U9909 (N_9909,N_7913,N_8206);
nor U9910 (N_9910,N_8569,N_8804);
or U9911 (N_9911,N_8810,N_7530);
nand U9912 (N_9912,N_8260,N_8827);
nand U9913 (N_9913,N_8833,N_7638);
or U9914 (N_9914,N_8167,N_8714);
nor U9915 (N_9915,N_8672,N_8017);
or U9916 (N_9916,N_8061,N_7849);
nand U9917 (N_9917,N_7888,N_7875);
nor U9918 (N_9918,N_8230,N_8292);
nand U9919 (N_9919,N_8347,N_7696);
nor U9920 (N_9920,N_7623,N_8569);
and U9921 (N_9921,N_7642,N_7821);
xor U9922 (N_9922,N_7863,N_8220);
nand U9923 (N_9923,N_7686,N_7529);
nand U9924 (N_9924,N_8488,N_8075);
and U9925 (N_9925,N_7864,N_7902);
xor U9926 (N_9926,N_8682,N_7917);
nor U9927 (N_9927,N_7982,N_8833);
nand U9928 (N_9928,N_8100,N_8418);
and U9929 (N_9929,N_8131,N_8785);
or U9930 (N_9930,N_7655,N_8649);
xor U9931 (N_9931,N_7789,N_7824);
and U9932 (N_9932,N_7832,N_8625);
or U9933 (N_9933,N_7776,N_7614);
and U9934 (N_9934,N_8179,N_7994);
and U9935 (N_9935,N_7713,N_8355);
nor U9936 (N_9936,N_8280,N_7712);
nand U9937 (N_9937,N_8429,N_8286);
and U9938 (N_9938,N_8115,N_7669);
nand U9939 (N_9939,N_8012,N_7514);
nand U9940 (N_9940,N_8986,N_7567);
and U9941 (N_9941,N_8472,N_8204);
nor U9942 (N_9942,N_8248,N_8355);
or U9943 (N_9943,N_8977,N_8563);
nor U9944 (N_9944,N_7933,N_8995);
nand U9945 (N_9945,N_8847,N_8255);
nand U9946 (N_9946,N_8757,N_8279);
and U9947 (N_9947,N_8064,N_8244);
and U9948 (N_9948,N_7789,N_8698);
nand U9949 (N_9949,N_8788,N_8578);
or U9950 (N_9950,N_8771,N_8153);
and U9951 (N_9951,N_8027,N_8374);
nand U9952 (N_9952,N_7655,N_8453);
nand U9953 (N_9953,N_8470,N_8592);
and U9954 (N_9954,N_8315,N_7567);
nand U9955 (N_9955,N_8005,N_8195);
and U9956 (N_9956,N_8636,N_8458);
and U9957 (N_9957,N_8960,N_7607);
or U9958 (N_9958,N_8575,N_8468);
nand U9959 (N_9959,N_8803,N_7928);
nand U9960 (N_9960,N_8689,N_8878);
nand U9961 (N_9961,N_7936,N_7727);
nor U9962 (N_9962,N_7747,N_7531);
nor U9963 (N_9963,N_8424,N_8749);
and U9964 (N_9964,N_8656,N_7739);
or U9965 (N_9965,N_8810,N_7901);
or U9966 (N_9966,N_7522,N_8988);
and U9967 (N_9967,N_8803,N_8897);
nor U9968 (N_9968,N_8818,N_7569);
and U9969 (N_9969,N_7591,N_8486);
xnor U9970 (N_9970,N_8554,N_8956);
xnor U9971 (N_9971,N_7720,N_8909);
nor U9972 (N_9972,N_8551,N_8648);
or U9973 (N_9973,N_8755,N_8173);
and U9974 (N_9974,N_8563,N_8848);
nor U9975 (N_9975,N_8810,N_7560);
or U9976 (N_9976,N_8065,N_8586);
and U9977 (N_9977,N_7885,N_8400);
nand U9978 (N_9978,N_8716,N_7773);
or U9979 (N_9979,N_8284,N_7718);
xnor U9980 (N_9980,N_8386,N_8532);
nand U9981 (N_9981,N_7610,N_8529);
or U9982 (N_9982,N_8074,N_7573);
and U9983 (N_9983,N_8499,N_8229);
or U9984 (N_9984,N_7648,N_7798);
or U9985 (N_9985,N_8877,N_7812);
nand U9986 (N_9986,N_8922,N_7504);
or U9987 (N_9987,N_8324,N_7953);
or U9988 (N_9988,N_8786,N_7630);
or U9989 (N_9989,N_7776,N_8303);
or U9990 (N_9990,N_8564,N_8886);
nor U9991 (N_9991,N_8313,N_7789);
or U9992 (N_9992,N_8431,N_8470);
nor U9993 (N_9993,N_8947,N_7993);
nand U9994 (N_9994,N_8100,N_7555);
nor U9995 (N_9995,N_7759,N_8728);
or U9996 (N_9996,N_7687,N_8641);
and U9997 (N_9997,N_8312,N_8479);
and U9998 (N_9998,N_8864,N_7576);
and U9999 (N_9999,N_8242,N_8233);
nand U10000 (N_10000,N_8390,N_7772);
nand U10001 (N_10001,N_8338,N_8047);
and U10002 (N_10002,N_8808,N_7743);
nand U10003 (N_10003,N_7798,N_8794);
nand U10004 (N_10004,N_7666,N_8077);
nand U10005 (N_10005,N_8235,N_8733);
or U10006 (N_10006,N_8022,N_8253);
or U10007 (N_10007,N_8532,N_8118);
or U10008 (N_10008,N_7846,N_7643);
nor U10009 (N_10009,N_7693,N_7555);
nand U10010 (N_10010,N_8743,N_8572);
nor U10011 (N_10011,N_8719,N_7576);
nor U10012 (N_10012,N_7547,N_7672);
and U10013 (N_10013,N_8101,N_8669);
nand U10014 (N_10014,N_7858,N_8491);
nor U10015 (N_10015,N_8664,N_8746);
xnor U10016 (N_10016,N_7825,N_7545);
and U10017 (N_10017,N_8896,N_8812);
and U10018 (N_10018,N_8344,N_7654);
xor U10019 (N_10019,N_7646,N_8800);
and U10020 (N_10020,N_8733,N_7648);
or U10021 (N_10021,N_7708,N_7602);
or U10022 (N_10022,N_7710,N_8790);
nand U10023 (N_10023,N_8832,N_8107);
nor U10024 (N_10024,N_8842,N_8657);
or U10025 (N_10025,N_8282,N_8796);
nand U10026 (N_10026,N_8899,N_7760);
or U10027 (N_10027,N_7777,N_8678);
nor U10028 (N_10028,N_8093,N_8937);
and U10029 (N_10029,N_8717,N_8227);
or U10030 (N_10030,N_8685,N_7666);
nor U10031 (N_10031,N_8920,N_8075);
nor U10032 (N_10032,N_7848,N_8394);
xor U10033 (N_10033,N_7673,N_8350);
and U10034 (N_10034,N_8360,N_7961);
nand U10035 (N_10035,N_8079,N_8919);
or U10036 (N_10036,N_7525,N_8127);
nand U10037 (N_10037,N_8210,N_8477);
xor U10038 (N_10038,N_7621,N_7527);
nor U10039 (N_10039,N_7589,N_8862);
nand U10040 (N_10040,N_8129,N_7672);
nand U10041 (N_10041,N_7857,N_8744);
and U10042 (N_10042,N_8036,N_7507);
nor U10043 (N_10043,N_7946,N_8789);
and U10044 (N_10044,N_7531,N_8683);
nand U10045 (N_10045,N_7945,N_7805);
nand U10046 (N_10046,N_8906,N_7667);
nand U10047 (N_10047,N_8940,N_8699);
nor U10048 (N_10048,N_8712,N_7599);
or U10049 (N_10049,N_8076,N_8211);
nor U10050 (N_10050,N_8051,N_8840);
nor U10051 (N_10051,N_7754,N_8773);
xor U10052 (N_10052,N_7664,N_8086);
xor U10053 (N_10053,N_7519,N_8601);
nor U10054 (N_10054,N_8323,N_8419);
and U10055 (N_10055,N_8500,N_7900);
nor U10056 (N_10056,N_7846,N_7545);
and U10057 (N_10057,N_8399,N_7775);
nand U10058 (N_10058,N_8049,N_7609);
xnor U10059 (N_10059,N_7965,N_7918);
nand U10060 (N_10060,N_8085,N_8617);
nand U10061 (N_10061,N_8283,N_7818);
and U10062 (N_10062,N_8907,N_8924);
xor U10063 (N_10063,N_8621,N_8414);
nand U10064 (N_10064,N_8285,N_8791);
or U10065 (N_10065,N_7958,N_8770);
xnor U10066 (N_10066,N_8740,N_8357);
or U10067 (N_10067,N_8360,N_7673);
nor U10068 (N_10068,N_8776,N_8672);
nand U10069 (N_10069,N_8731,N_7924);
nand U10070 (N_10070,N_7639,N_8245);
nor U10071 (N_10071,N_7860,N_7602);
nor U10072 (N_10072,N_8598,N_8748);
nand U10073 (N_10073,N_8902,N_8516);
nor U10074 (N_10074,N_7948,N_7910);
and U10075 (N_10075,N_8145,N_8703);
and U10076 (N_10076,N_7838,N_8576);
or U10077 (N_10077,N_8767,N_8198);
and U10078 (N_10078,N_7827,N_8397);
nor U10079 (N_10079,N_7926,N_8418);
nor U10080 (N_10080,N_8869,N_7843);
xor U10081 (N_10081,N_7757,N_7830);
and U10082 (N_10082,N_8409,N_8262);
xnor U10083 (N_10083,N_7577,N_7745);
or U10084 (N_10084,N_7605,N_7935);
nor U10085 (N_10085,N_8752,N_8202);
or U10086 (N_10086,N_7565,N_8096);
and U10087 (N_10087,N_8265,N_7934);
and U10088 (N_10088,N_8312,N_8005);
and U10089 (N_10089,N_7644,N_8177);
and U10090 (N_10090,N_8759,N_7627);
nor U10091 (N_10091,N_7517,N_7850);
nor U10092 (N_10092,N_8922,N_8440);
nor U10093 (N_10093,N_8342,N_7589);
nand U10094 (N_10094,N_7592,N_7555);
and U10095 (N_10095,N_8737,N_7891);
xnor U10096 (N_10096,N_8776,N_8368);
nand U10097 (N_10097,N_7887,N_7933);
xor U10098 (N_10098,N_8554,N_8306);
nand U10099 (N_10099,N_7874,N_7586);
or U10100 (N_10100,N_7873,N_8904);
nand U10101 (N_10101,N_7604,N_8254);
nor U10102 (N_10102,N_8071,N_8512);
nor U10103 (N_10103,N_8411,N_7508);
or U10104 (N_10104,N_7981,N_7681);
and U10105 (N_10105,N_7712,N_8705);
nand U10106 (N_10106,N_8131,N_7650);
nor U10107 (N_10107,N_8084,N_7685);
or U10108 (N_10108,N_8334,N_8956);
and U10109 (N_10109,N_8047,N_8261);
and U10110 (N_10110,N_7957,N_8066);
or U10111 (N_10111,N_8962,N_8243);
nand U10112 (N_10112,N_8783,N_8223);
nand U10113 (N_10113,N_7559,N_8811);
nand U10114 (N_10114,N_8270,N_8922);
nand U10115 (N_10115,N_7869,N_8454);
or U10116 (N_10116,N_8157,N_8144);
nand U10117 (N_10117,N_7568,N_7513);
and U10118 (N_10118,N_8141,N_8710);
and U10119 (N_10119,N_7566,N_8009);
and U10120 (N_10120,N_8544,N_8770);
xor U10121 (N_10121,N_8012,N_8846);
or U10122 (N_10122,N_8575,N_7795);
nor U10123 (N_10123,N_8637,N_8943);
or U10124 (N_10124,N_7878,N_7669);
and U10125 (N_10125,N_8651,N_8730);
and U10126 (N_10126,N_8666,N_8674);
nor U10127 (N_10127,N_8558,N_8563);
nand U10128 (N_10128,N_8388,N_8913);
nand U10129 (N_10129,N_8688,N_8438);
and U10130 (N_10130,N_8020,N_7921);
xor U10131 (N_10131,N_8399,N_8955);
nor U10132 (N_10132,N_8850,N_8714);
nor U10133 (N_10133,N_7709,N_7780);
nor U10134 (N_10134,N_7618,N_8885);
nand U10135 (N_10135,N_7694,N_8539);
and U10136 (N_10136,N_8593,N_8413);
xnor U10137 (N_10137,N_8006,N_7959);
nor U10138 (N_10138,N_8754,N_7561);
nand U10139 (N_10139,N_8573,N_8484);
nor U10140 (N_10140,N_8209,N_7559);
and U10141 (N_10141,N_8899,N_7516);
nand U10142 (N_10142,N_8568,N_7749);
nor U10143 (N_10143,N_8477,N_8179);
nand U10144 (N_10144,N_7763,N_8098);
or U10145 (N_10145,N_8105,N_8013);
nand U10146 (N_10146,N_8473,N_7576);
or U10147 (N_10147,N_8100,N_7557);
nor U10148 (N_10148,N_8249,N_8239);
or U10149 (N_10149,N_8124,N_8589);
and U10150 (N_10150,N_7877,N_7664);
or U10151 (N_10151,N_8893,N_8543);
xor U10152 (N_10152,N_8754,N_7816);
xnor U10153 (N_10153,N_7951,N_8902);
or U10154 (N_10154,N_8831,N_7594);
and U10155 (N_10155,N_8152,N_8659);
or U10156 (N_10156,N_8104,N_7696);
and U10157 (N_10157,N_8302,N_8418);
nor U10158 (N_10158,N_7923,N_7911);
or U10159 (N_10159,N_8921,N_7850);
nand U10160 (N_10160,N_8104,N_8740);
and U10161 (N_10161,N_7814,N_8700);
nor U10162 (N_10162,N_7800,N_8392);
nor U10163 (N_10163,N_8723,N_8626);
nand U10164 (N_10164,N_8588,N_8842);
nand U10165 (N_10165,N_8776,N_7588);
or U10166 (N_10166,N_8688,N_8583);
nand U10167 (N_10167,N_7627,N_7553);
nor U10168 (N_10168,N_7544,N_7932);
or U10169 (N_10169,N_7521,N_8712);
and U10170 (N_10170,N_8163,N_8492);
nor U10171 (N_10171,N_8764,N_7695);
nor U10172 (N_10172,N_7539,N_7970);
nand U10173 (N_10173,N_8454,N_8318);
and U10174 (N_10174,N_7753,N_7966);
or U10175 (N_10175,N_7814,N_8441);
nor U10176 (N_10176,N_8706,N_8382);
nor U10177 (N_10177,N_7596,N_7518);
or U10178 (N_10178,N_8763,N_8382);
nor U10179 (N_10179,N_8550,N_7558);
nand U10180 (N_10180,N_8289,N_8519);
and U10181 (N_10181,N_7902,N_8573);
or U10182 (N_10182,N_8111,N_8900);
nor U10183 (N_10183,N_7574,N_7597);
xor U10184 (N_10184,N_8683,N_8047);
or U10185 (N_10185,N_8041,N_8058);
nand U10186 (N_10186,N_7757,N_7954);
or U10187 (N_10187,N_7527,N_8368);
or U10188 (N_10188,N_7799,N_8842);
nand U10189 (N_10189,N_8526,N_8495);
nand U10190 (N_10190,N_8914,N_7659);
xnor U10191 (N_10191,N_8534,N_8425);
and U10192 (N_10192,N_8154,N_7780);
and U10193 (N_10193,N_8636,N_8591);
or U10194 (N_10194,N_8834,N_8006);
and U10195 (N_10195,N_8748,N_7635);
and U10196 (N_10196,N_8087,N_8835);
xor U10197 (N_10197,N_7861,N_7618);
nor U10198 (N_10198,N_8443,N_8474);
nor U10199 (N_10199,N_8962,N_7520);
or U10200 (N_10200,N_8333,N_8277);
nand U10201 (N_10201,N_8830,N_7515);
nand U10202 (N_10202,N_7787,N_8698);
or U10203 (N_10203,N_8430,N_8434);
nand U10204 (N_10204,N_8648,N_7859);
and U10205 (N_10205,N_8631,N_8276);
xnor U10206 (N_10206,N_8303,N_7511);
xor U10207 (N_10207,N_8727,N_8482);
nand U10208 (N_10208,N_8747,N_8630);
or U10209 (N_10209,N_7516,N_7936);
nand U10210 (N_10210,N_7933,N_8955);
nand U10211 (N_10211,N_8529,N_7908);
nand U10212 (N_10212,N_8530,N_8629);
xnor U10213 (N_10213,N_8940,N_7582);
xor U10214 (N_10214,N_8162,N_8235);
or U10215 (N_10215,N_8368,N_7901);
nand U10216 (N_10216,N_7705,N_8917);
and U10217 (N_10217,N_7559,N_8143);
nand U10218 (N_10218,N_8470,N_8389);
and U10219 (N_10219,N_7549,N_8485);
nor U10220 (N_10220,N_7962,N_7716);
nand U10221 (N_10221,N_8352,N_8253);
or U10222 (N_10222,N_8010,N_7730);
nand U10223 (N_10223,N_8326,N_7741);
and U10224 (N_10224,N_8727,N_7799);
or U10225 (N_10225,N_7988,N_8665);
nor U10226 (N_10226,N_8950,N_8967);
and U10227 (N_10227,N_8026,N_8090);
and U10228 (N_10228,N_8315,N_8900);
nor U10229 (N_10229,N_8241,N_7960);
and U10230 (N_10230,N_7787,N_7713);
nor U10231 (N_10231,N_8549,N_8189);
and U10232 (N_10232,N_8188,N_7892);
nor U10233 (N_10233,N_7848,N_7618);
nor U10234 (N_10234,N_7966,N_7852);
and U10235 (N_10235,N_8682,N_7598);
nand U10236 (N_10236,N_7691,N_7710);
or U10237 (N_10237,N_8009,N_7909);
nor U10238 (N_10238,N_7756,N_8530);
or U10239 (N_10239,N_8669,N_8293);
nand U10240 (N_10240,N_7620,N_7938);
nor U10241 (N_10241,N_8920,N_8998);
xor U10242 (N_10242,N_7978,N_7596);
or U10243 (N_10243,N_7818,N_8900);
nand U10244 (N_10244,N_8026,N_8801);
or U10245 (N_10245,N_8847,N_8818);
nor U10246 (N_10246,N_8492,N_8153);
nor U10247 (N_10247,N_8783,N_7773);
or U10248 (N_10248,N_8606,N_8491);
nand U10249 (N_10249,N_8519,N_8811);
and U10250 (N_10250,N_8830,N_8405);
and U10251 (N_10251,N_7518,N_8294);
xnor U10252 (N_10252,N_7669,N_8498);
nand U10253 (N_10253,N_8631,N_8939);
or U10254 (N_10254,N_8320,N_8814);
or U10255 (N_10255,N_8973,N_8231);
and U10256 (N_10256,N_8195,N_7974);
nor U10257 (N_10257,N_7972,N_8500);
xnor U10258 (N_10258,N_8874,N_8867);
or U10259 (N_10259,N_7504,N_8467);
nor U10260 (N_10260,N_8724,N_8769);
or U10261 (N_10261,N_8946,N_7524);
and U10262 (N_10262,N_8903,N_7547);
nor U10263 (N_10263,N_7721,N_8436);
or U10264 (N_10264,N_7720,N_7717);
nor U10265 (N_10265,N_7998,N_7567);
or U10266 (N_10266,N_8744,N_8266);
nand U10267 (N_10267,N_8941,N_8496);
or U10268 (N_10268,N_7823,N_7925);
and U10269 (N_10269,N_8461,N_8753);
or U10270 (N_10270,N_8311,N_8999);
nor U10271 (N_10271,N_8121,N_8462);
nor U10272 (N_10272,N_8475,N_8865);
and U10273 (N_10273,N_8922,N_7762);
or U10274 (N_10274,N_7887,N_8430);
nand U10275 (N_10275,N_8301,N_8231);
nor U10276 (N_10276,N_8856,N_7750);
nor U10277 (N_10277,N_7510,N_8437);
and U10278 (N_10278,N_8190,N_7889);
and U10279 (N_10279,N_7641,N_8036);
nand U10280 (N_10280,N_8450,N_8800);
nand U10281 (N_10281,N_8224,N_8589);
and U10282 (N_10282,N_8760,N_8248);
nand U10283 (N_10283,N_8206,N_8584);
or U10284 (N_10284,N_7763,N_8872);
nand U10285 (N_10285,N_7595,N_7810);
nor U10286 (N_10286,N_8403,N_8171);
and U10287 (N_10287,N_8286,N_7733);
nor U10288 (N_10288,N_8642,N_8564);
and U10289 (N_10289,N_8251,N_7553);
nand U10290 (N_10290,N_7612,N_7604);
or U10291 (N_10291,N_7589,N_8236);
nor U10292 (N_10292,N_8304,N_7779);
nor U10293 (N_10293,N_7806,N_8430);
nor U10294 (N_10294,N_8525,N_7569);
and U10295 (N_10295,N_8883,N_8184);
and U10296 (N_10296,N_8323,N_8162);
and U10297 (N_10297,N_8140,N_8421);
nand U10298 (N_10298,N_8002,N_8156);
and U10299 (N_10299,N_7956,N_8276);
and U10300 (N_10300,N_8903,N_7753);
nor U10301 (N_10301,N_8332,N_8511);
nand U10302 (N_10302,N_7822,N_7673);
nor U10303 (N_10303,N_8149,N_7812);
nand U10304 (N_10304,N_7701,N_8273);
xor U10305 (N_10305,N_8164,N_8908);
nor U10306 (N_10306,N_7916,N_7724);
and U10307 (N_10307,N_8546,N_8233);
nor U10308 (N_10308,N_8630,N_8923);
and U10309 (N_10309,N_7870,N_7929);
nor U10310 (N_10310,N_8313,N_8257);
nor U10311 (N_10311,N_8835,N_8070);
nor U10312 (N_10312,N_7589,N_8420);
xnor U10313 (N_10313,N_8255,N_8911);
or U10314 (N_10314,N_8419,N_7995);
nand U10315 (N_10315,N_8559,N_8218);
and U10316 (N_10316,N_8713,N_8695);
nor U10317 (N_10317,N_8062,N_8955);
and U10318 (N_10318,N_7570,N_7730);
and U10319 (N_10319,N_8906,N_8349);
nand U10320 (N_10320,N_7694,N_8969);
nand U10321 (N_10321,N_8687,N_8036);
nor U10322 (N_10322,N_7772,N_7973);
or U10323 (N_10323,N_7658,N_8972);
or U10324 (N_10324,N_8812,N_8305);
nand U10325 (N_10325,N_8253,N_7812);
nor U10326 (N_10326,N_8175,N_7737);
and U10327 (N_10327,N_7893,N_7867);
xor U10328 (N_10328,N_8506,N_7774);
nand U10329 (N_10329,N_7637,N_8702);
nand U10330 (N_10330,N_8219,N_7954);
or U10331 (N_10331,N_7691,N_7600);
nor U10332 (N_10332,N_7566,N_8784);
nand U10333 (N_10333,N_8970,N_7603);
nand U10334 (N_10334,N_8276,N_8364);
xor U10335 (N_10335,N_7621,N_7573);
or U10336 (N_10336,N_8931,N_8780);
and U10337 (N_10337,N_8617,N_8639);
nor U10338 (N_10338,N_8993,N_8635);
nand U10339 (N_10339,N_8958,N_8893);
and U10340 (N_10340,N_8110,N_8274);
nor U10341 (N_10341,N_8432,N_8145);
and U10342 (N_10342,N_8145,N_8748);
nand U10343 (N_10343,N_7732,N_8375);
nand U10344 (N_10344,N_8429,N_8559);
and U10345 (N_10345,N_7628,N_8757);
or U10346 (N_10346,N_7787,N_7880);
nor U10347 (N_10347,N_8665,N_8280);
nor U10348 (N_10348,N_7618,N_8467);
and U10349 (N_10349,N_8650,N_7821);
xor U10350 (N_10350,N_8617,N_8785);
or U10351 (N_10351,N_7651,N_8005);
xnor U10352 (N_10352,N_7528,N_7910);
or U10353 (N_10353,N_8616,N_8054);
or U10354 (N_10354,N_8953,N_8470);
nor U10355 (N_10355,N_8061,N_8001);
and U10356 (N_10356,N_7769,N_7593);
nor U10357 (N_10357,N_7963,N_7689);
xor U10358 (N_10358,N_7552,N_8906);
nand U10359 (N_10359,N_8602,N_8432);
nand U10360 (N_10360,N_7583,N_8466);
nand U10361 (N_10361,N_8979,N_7919);
nand U10362 (N_10362,N_7655,N_8851);
nand U10363 (N_10363,N_8394,N_8264);
or U10364 (N_10364,N_7594,N_8855);
or U10365 (N_10365,N_8245,N_8942);
nor U10366 (N_10366,N_8867,N_7952);
and U10367 (N_10367,N_8488,N_8976);
and U10368 (N_10368,N_8579,N_8294);
nor U10369 (N_10369,N_7866,N_7963);
nand U10370 (N_10370,N_8143,N_8963);
nand U10371 (N_10371,N_7647,N_7929);
xnor U10372 (N_10372,N_8159,N_7856);
and U10373 (N_10373,N_8101,N_8555);
and U10374 (N_10374,N_8295,N_7639);
nand U10375 (N_10375,N_8154,N_7957);
and U10376 (N_10376,N_8177,N_7895);
nor U10377 (N_10377,N_8816,N_7897);
nand U10378 (N_10378,N_8508,N_7727);
nand U10379 (N_10379,N_8514,N_7814);
and U10380 (N_10380,N_8323,N_7626);
and U10381 (N_10381,N_8409,N_8737);
or U10382 (N_10382,N_7937,N_8641);
or U10383 (N_10383,N_8308,N_7787);
nor U10384 (N_10384,N_8302,N_7737);
or U10385 (N_10385,N_8294,N_8478);
xnor U10386 (N_10386,N_8498,N_7582);
nand U10387 (N_10387,N_8421,N_8350);
nand U10388 (N_10388,N_8006,N_8812);
and U10389 (N_10389,N_7788,N_7924);
nor U10390 (N_10390,N_8855,N_8412);
nor U10391 (N_10391,N_8007,N_8544);
nand U10392 (N_10392,N_7674,N_8881);
nand U10393 (N_10393,N_7772,N_7873);
xnor U10394 (N_10394,N_8350,N_8756);
nor U10395 (N_10395,N_7699,N_8469);
or U10396 (N_10396,N_7972,N_7812);
nand U10397 (N_10397,N_8846,N_8799);
and U10398 (N_10398,N_8419,N_8601);
nand U10399 (N_10399,N_8523,N_8388);
or U10400 (N_10400,N_8210,N_8179);
or U10401 (N_10401,N_8803,N_8231);
nand U10402 (N_10402,N_8604,N_8233);
and U10403 (N_10403,N_8920,N_7707);
nor U10404 (N_10404,N_8170,N_8371);
nor U10405 (N_10405,N_8202,N_7805);
nor U10406 (N_10406,N_8233,N_8200);
nor U10407 (N_10407,N_8916,N_8650);
and U10408 (N_10408,N_8780,N_7614);
xnor U10409 (N_10409,N_8166,N_8724);
nor U10410 (N_10410,N_8246,N_8722);
nand U10411 (N_10411,N_8598,N_8235);
and U10412 (N_10412,N_7631,N_7521);
nor U10413 (N_10413,N_7610,N_8231);
nor U10414 (N_10414,N_7816,N_8807);
xor U10415 (N_10415,N_8707,N_8397);
or U10416 (N_10416,N_8236,N_7818);
and U10417 (N_10417,N_8235,N_7703);
nand U10418 (N_10418,N_8603,N_8539);
nor U10419 (N_10419,N_8826,N_7975);
nor U10420 (N_10420,N_8983,N_7558);
nand U10421 (N_10421,N_8021,N_7807);
xnor U10422 (N_10422,N_7740,N_8240);
nor U10423 (N_10423,N_7777,N_8993);
or U10424 (N_10424,N_7647,N_8633);
nand U10425 (N_10425,N_8424,N_8631);
nor U10426 (N_10426,N_7736,N_7545);
xnor U10427 (N_10427,N_8171,N_7572);
or U10428 (N_10428,N_8715,N_7667);
nand U10429 (N_10429,N_7885,N_8761);
nand U10430 (N_10430,N_7520,N_8102);
xnor U10431 (N_10431,N_8179,N_8876);
nor U10432 (N_10432,N_8934,N_8157);
nand U10433 (N_10433,N_7901,N_8562);
or U10434 (N_10434,N_8306,N_8907);
or U10435 (N_10435,N_8885,N_8361);
and U10436 (N_10436,N_8207,N_7814);
and U10437 (N_10437,N_8895,N_7968);
nor U10438 (N_10438,N_8565,N_7690);
or U10439 (N_10439,N_8999,N_7998);
or U10440 (N_10440,N_7597,N_8728);
nand U10441 (N_10441,N_8754,N_7900);
nand U10442 (N_10442,N_7979,N_8469);
and U10443 (N_10443,N_8868,N_7765);
or U10444 (N_10444,N_8159,N_8383);
nor U10445 (N_10445,N_8841,N_8101);
xor U10446 (N_10446,N_8276,N_8921);
nor U10447 (N_10447,N_8700,N_8082);
or U10448 (N_10448,N_8382,N_8734);
and U10449 (N_10449,N_7886,N_7969);
or U10450 (N_10450,N_8086,N_8041);
xor U10451 (N_10451,N_8202,N_8911);
nand U10452 (N_10452,N_8754,N_7858);
nor U10453 (N_10453,N_8120,N_7837);
and U10454 (N_10454,N_8678,N_8685);
and U10455 (N_10455,N_8438,N_8245);
or U10456 (N_10456,N_8462,N_7577);
and U10457 (N_10457,N_8039,N_8022);
nand U10458 (N_10458,N_8321,N_7862);
xnor U10459 (N_10459,N_7853,N_8993);
xnor U10460 (N_10460,N_7670,N_8294);
nand U10461 (N_10461,N_8917,N_8299);
and U10462 (N_10462,N_8794,N_8912);
xor U10463 (N_10463,N_7622,N_8487);
nor U10464 (N_10464,N_8706,N_8207);
and U10465 (N_10465,N_8141,N_7858);
nor U10466 (N_10466,N_8576,N_7771);
or U10467 (N_10467,N_7751,N_7916);
and U10468 (N_10468,N_7621,N_8260);
nor U10469 (N_10469,N_8061,N_8600);
nor U10470 (N_10470,N_7584,N_7995);
nor U10471 (N_10471,N_8321,N_8723);
nor U10472 (N_10472,N_7888,N_7941);
or U10473 (N_10473,N_8626,N_7541);
nor U10474 (N_10474,N_7758,N_8673);
or U10475 (N_10475,N_8079,N_8151);
nand U10476 (N_10476,N_8793,N_7708);
nand U10477 (N_10477,N_8080,N_8576);
nand U10478 (N_10478,N_7907,N_8252);
and U10479 (N_10479,N_8529,N_7957);
nand U10480 (N_10480,N_8820,N_8712);
nand U10481 (N_10481,N_8428,N_8273);
and U10482 (N_10482,N_8011,N_8782);
and U10483 (N_10483,N_8072,N_8241);
nor U10484 (N_10484,N_8210,N_7724);
and U10485 (N_10485,N_8991,N_8997);
nand U10486 (N_10486,N_8531,N_8545);
or U10487 (N_10487,N_8086,N_7549);
and U10488 (N_10488,N_8010,N_8908);
nor U10489 (N_10489,N_7697,N_8693);
xor U10490 (N_10490,N_8266,N_7583);
or U10491 (N_10491,N_8940,N_8910);
and U10492 (N_10492,N_8784,N_8673);
and U10493 (N_10493,N_8195,N_7610);
nor U10494 (N_10494,N_7648,N_8960);
nand U10495 (N_10495,N_8401,N_8965);
and U10496 (N_10496,N_8960,N_7895);
and U10497 (N_10497,N_8003,N_8379);
xnor U10498 (N_10498,N_8005,N_7934);
xnor U10499 (N_10499,N_8736,N_8382);
nand U10500 (N_10500,N_9946,N_9578);
or U10501 (N_10501,N_9563,N_10295);
or U10502 (N_10502,N_9020,N_10340);
nor U10503 (N_10503,N_9721,N_10100);
nor U10504 (N_10504,N_9664,N_9099);
and U10505 (N_10505,N_9419,N_9189);
nor U10506 (N_10506,N_9488,N_9276);
or U10507 (N_10507,N_10071,N_9512);
nor U10508 (N_10508,N_9595,N_10087);
nand U10509 (N_10509,N_10183,N_10229);
xnor U10510 (N_10510,N_10239,N_9536);
xor U10511 (N_10511,N_9299,N_9628);
or U10512 (N_10512,N_9001,N_9669);
nor U10513 (N_10513,N_9989,N_10434);
and U10514 (N_10514,N_9702,N_9275);
or U10515 (N_10515,N_9928,N_10163);
or U10516 (N_10516,N_9591,N_10221);
and U10517 (N_10517,N_9371,N_9794);
and U10518 (N_10518,N_9178,N_10277);
or U10519 (N_10519,N_9881,N_9040);
or U10520 (N_10520,N_9801,N_10098);
nor U10521 (N_10521,N_9997,N_9498);
and U10522 (N_10522,N_9703,N_9974);
nand U10523 (N_10523,N_9747,N_10290);
and U10524 (N_10524,N_10132,N_10164);
or U10525 (N_10525,N_9463,N_9384);
nor U10526 (N_10526,N_9435,N_9095);
and U10527 (N_10527,N_10218,N_9165);
and U10528 (N_10528,N_9810,N_9667);
and U10529 (N_10529,N_10155,N_10175);
xnor U10530 (N_10530,N_9056,N_9665);
xor U10531 (N_10531,N_9147,N_10390);
nor U10532 (N_10532,N_10343,N_9119);
and U10533 (N_10533,N_9107,N_10212);
and U10534 (N_10534,N_9809,N_9472);
or U10535 (N_10535,N_10234,N_9888);
nand U10536 (N_10536,N_9755,N_9060);
or U10537 (N_10537,N_10368,N_9726);
nand U10538 (N_10538,N_9865,N_9109);
or U10539 (N_10539,N_9210,N_9115);
or U10540 (N_10540,N_9994,N_9399);
or U10541 (N_10541,N_9026,N_9112);
xor U10542 (N_10542,N_9678,N_10282);
or U10543 (N_10543,N_9104,N_9295);
nor U10544 (N_10544,N_9693,N_10425);
xnor U10545 (N_10545,N_9137,N_10211);
or U10546 (N_10546,N_9013,N_9367);
and U10547 (N_10547,N_10418,N_9677);
and U10548 (N_10548,N_9818,N_9303);
or U10549 (N_10549,N_9788,N_9535);
and U10550 (N_10550,N_9869,N_10244);
nor U10551 (N_10551,N_10464,N_10350);
or U10552 (N_10552,N_9637,N_9722);
or U10553 (N_10553,N_10353,N_10135);
and U10554 (N_10554,N_9028,N_9938);
or U10555 (N_10555,N_10025,N_9904);
nand U10556 (N_10556,N_9256,N_9993);
and U10557 (N_10557,N_9270,N_9448);
and U10558 (N_10558,N_10344,N_9142);
xnor U10559 (N_10559,N_10382,N_9460);
and U10560 (N_10560,N_10176,N_10120);
and U10561 (N_10561,N_9261,N_10199);
or U10562 (N_10562,N_9288,N_10379);
nand U10563 (N_10563,N_9380,N_9279);
or U10564 (N_10564,N_9239,N_10012);
nor U10565 (N_10565,N_9530,N_9616);
or U10566 (N_10566,N_9424,N_10480);
nand U10567 (N_10567,N_10483,N_9971);
and U10568 (N_10568,N_10319,N_9635);
nor U10569 (N_10569,N_9324,N_9871);
and U10570 (N_10570,N_10198,N_9429);
and U10571 (N_10571,N_9127,N_10287);
nor U10572 (N_10572,N_9094,N_10044);
nand U10573 (N_10573,N_10494,N_9996);
nor U10574 (N_10574,N_10256,N_10424);
or U10575 (N_10575,N_9922,N_9786);
or U10576 (N_10576,N_9695,N_10197);
and U10577 (N_10577,N_9412,N_10479);
nor U10578 (N_10578,N_9929,N_9731);
nor U10579 (N_10579,N_9526,N_10094);
nor U10580 (N_10580,N_10193,N_9956);
or U10581 (N_10581,N_9668,N_9909);
and U10582 (N_10582,N_9290,N_10170);
nor U10583 (N_10583,N_9333,N_9305);
nor U10584 (N_10584,N_9552,N_9574);
nand U10585 (N_10585,N_9216,N_9255);
or U10586 (N_10586,N_9620,N_9840);
or U10587 (N_10587,N_9874,N_9245);
nor U10588 (N_10588,N_9402,N_9204);
nor U10589 (N_10589,N_10016,N_9867);
nor U10590 (N_10590,N_9209,N_9543);
nand U10591 (N_10591,N_9066,N_10428);
nor U10592 (N_10592,N_9999,N_10405);
xor U10593 (N_10593,N_9807,N_9579);
nand U10594 (N_10594,N_9700,N_9038);
nor U10595 (N_10595,N_9983,N_9483);
nor U10596 (N_10596,N_9467,N_9527);
and U10597 (N_10597,N_9666,N_9771);
nand U10598 (N_10598,N_9004,N_9886);
nor U10599 (N_10599,N_9051,N_9091);
and U10600 (N_10600,N_9745,N_10158);
nand U10601 (N_10601,N_9877,N_9344);
nor U10602 (N_10602,N_9798,N_9751);
nand U10603 (N_10603,N_9792,N_9141);
nand U10604 (N_10604,N_9673,N_9507);
nand U10605 (N_10605,N_10326,N_10118);
nor U10606 (N_10606,N_9846,N_10476);
or U10607 (N_10607,N_9200,N_10145);
or U10608 (N_10608,N_9732,N_10048);
and U10609 (N_10609,N_9738,N_9817);
or U10610 (N_10610,N_10423,N_9052);
and U10611 (N_10611,N_10219,N_9496);
nand U10612 (N_10612,N_10288,N_10137);
nand U10613 (N_10613,N_9864,N_10125);
nand U10614 (N_10614,N_10254,N_9943);
nand U10615 (N_10615,N_9674,N_10099);
and U10616 (N_10616,N_9553,N_9849);
nand U10617 (N_10617,N_9319,N_9699);
or U10618 (N_10618,N_9682,N_10307);
and U10619 (N_10619,N_9735,N_9623);
or U10620 (N_10620,N_9075,N_9005);
or U10621 (N_10621,N_9639,N_9898);
or U10622 (N_10622,N_9885,N_9833);
and U10623 (N_10623,N_9910,N_9438);
or U10624 (N_10624,N_9879,N_10299);
nor U10625 (N_10625,N_10462,N_9044);
nor U10626 (N_10626,N_9514,N_10124);
and U10627 (N_10627,N_9559,N_9876);
and U10628 (N_10628,N_9318,N_10321);
and U10629 (N_10629,N_9736,N_9440);
nor U10630 (N_10630,N_9043,N_9234);
nand U10631 (N_10631,N_9450,N_9133);
or U10632 (N_10632,N_9227,N_10113);
and U10633 (N_10633,N_9891,N_9401);
or U10634 (N_10634,N_9174,N_10066);
nand U10635 (N_10635,N_10093,N_9139);
or U10636 (N_10636,N_9701,N_10136);
nand U10637 (N_10637,N_10196,N_9734);
nor U10638 (N_10638,N_9847,N_9582);
or U10639 (N_10639,N_9179,N_9346);
and U10640 (N_10640,N_9158,N_9901);
nand U10641 (N_10641,N_9236,N_9386);
nand U10642 (N_10642,N_10156,N_10081);
nand U10643 (N_10643,N_9936,N_9378);
nand U10644 (N_10644,N_9832,N_10452);
and U10645 (N_10645,N_9336,N_9787);
xnor U10646 (N_10646,N_9980,N_9972);
nor U10647 (N_10647,N_10067,N_10465);
nand U10648 (N_10648,N_9311,N_9057);
and U10649 (N_10649,N_9638,N_10259);
and U10650 (N_10650,N_10057,N_9614);
nand U10651 (N_10651,N_10192,N_10236);
nand U10652 (N_10652,N_9949,N_9557);
or U10653 (N_10653,N_9629,N_10317);
nand U10654 (N_10654,N_9266,N_10050);
or U10655 (N_10655,N_10128,N_9073);
nor U10656 (N_10656,N_9491,N_9660);
or U10657 (N_10657,N_9358,N_9392);
nor U10658 (N_10658,N_10252,N_9328);
or U10659 (N_10659,N_9892,N_10348);
nor U10660 (N_10660,N_9243,N_9042);
or U10661 (N_10661,N_9015,N_9352);
and U10662 (N_10662,N_9457,N_10331);
and U10663 (N_10663,N_9377,N_9769);
or U10664 (N_10664,N_9500,N_9381);
nand U10665 (N_10665,N_9445,N_9636);
and U10666 (N_10666,N_9214,N_9171);
xnor U10667 (N_10667,N_9645,N_9173);
xor U10668 (N_10668,N_10130,N_10035);
nor U10669 (N_10669,N_10154,N_9505);
nand U10670 (N_10670,N_9430,N_10209);
or U10671 (N_10671,N_9725,N_9634);
nand U10672 (N_10672,N_9625,N_10274);
or U10673 (N_10673,N_10451,N_9427);
nor U10674 (N_10674,N_9215,N_10246);
xnor U10675 (N_10675,N_9195,N_9720);
or U10676 (N_10676,N_9785,N_9519);
or U10677 (N_10677,N_9254,N_9306);
and U10678 (N_10678,N_10381,N_9990);
nand U10679 (N_10679,N_9588,N_9393);
and U10680 (N_10680,N_9587,N_9548);
and U10681 (N_10681,N_10141,N_9838);
nor U10682 (N_10682,N_9229,N_10079);
and U10683 (N_10683,N_10315,N_9207);
nor U10684 (N_10684,N_9803,N_10126);
nand U10685 (N_10685,N_9768,N_9932);
or U10686 (N_10686,N_10449,N_9053);
and U10687 (N_10687,N_9325,N_10247);
xor U10688 (N_10688,N_10261,N_10152);
xor U10689 (N_10689,N_10284,N_9580);
nand U10690 (N_10690,N_9469,N_10408);
xnor U10691 (N_10691,N_9024,N_10371);
nor U10692 (N_10692,N_9744,N_9055);
or U10693 (N_10693,N_9630,N_9839);
and U10694 (N_10694,N_9296,N_10028);
or U10695 (N_10695,N_10024,N_9193);
nor U10696 (N_10696,N_10092,N_9062);
or U10697 (N_10697,N_10454,N_9281);
nand U10698 (N_10698,N_9723,N_9120);
or U10699 (N_10699,N_10358,N_9866);
xor U10700 (N_10700,N_10401,N_9259);
nand U10701 (N_10701,N_10032,N_10478);
nand U10702 (N_10702,N_9068,N_10351);
and U10703 (N_10703,N_10090,N_9230);
and U10704 (N_10704,N_10105,N_9691);
or U10705 (N_10705,N_10160,N_9389);
or U10706 (N_10706,N_10324,N_10460);
and U10707 (N_10707,N_10232,N_9730);
xor U10708 (N_10708,N_9397,N_9883);
nor U10709 (N_10709,N_10322,N_10265);
and U10710 (N_10710,N_9640,N_9233);
or U10711 (N_10711,N_9777,N_9036);
and U10712 (N_10712,N_10041,N_9117);
or U10713 (N_10713,N_9544,N_9627);
nor U10714 (N_10714,N_10360,N_9716);
and U10715 (N_10715,N_9237,N_10419);
nor U10716 (N_10716,N_9799,N_9379);
nor U10717 (N_10717,N_9287,N_10151);
or U10718 (N_10718,N_9485,N_9184);
and U10719 (N_10719,N_10139,N_10293);
nand U10720 (N_10720,N_9136,N_9610);
nand U10721 (N_10721,N_9258,N_9297);
nand U10722 (N_10722,N_9850,N_10409);
nand U10723 (N_10723,N_9729,N_10171);
and U10724 (N_10724,N_9415,N_9495);
and U10725 (N_10725,N_10332,N_9571);
nand U10726 (N_10726,N_9606,N_9294);
and U10727 (N_10727,N_9915,N_9513);
and U10728 (N_10728,N_9170,N_10091);
nor U10729 (N_10729,N_9684,N_10426);
nor U10730 (N_10730,N_10227,N_9893);
and U10731 (N_10731,N_9811,N_9025);
nand U10732 (N_10732,N_10445,N_9081);
or U10733 (N_10733,N_9742,N_9824);
nor U10734 (N_10734,N_9903,N_9454);
and U10735 (N_10735,N_10251,N_9219);
or U10736 (N_10736,N_9315,N_9965);
and U10737 (N_10737,N_9208,N_9451);
nor U10738 (N_10738,N_10365,N_9316);
or U10739 (N_10739,N_9187,N_9842);
xnor U10740 (N_10740,N_10301,N_9271);
and U10741 (N_10741,N_9941,N_10179);
nor U10742 (N_10742,N_9767,N_10297);
nor U10743 (N_10743,N_9308,N_9948);
nor U10744 (N_10744,N_9781,N_10377);
or U10745 (N_10745,N_10439,N_9672);
xor U10746 (N_10746,N_10202,N_9688);
or U10747 (N_10747,N_9641,N_9357);
nand U10748 (N_10748,N_10009,N_10159);
nor U10749 (N_10749,N_9719,N_9861);
or U10750 (N_10750,N_9851,N_9696);
xnor U10751 (N_10751,N_9649,N_9033);
nand U10752 (N_10752,N_9776,N_9520);
xor U10753 (N_10753,N_9128,N_9391);
nor U10754 (N_10754,N_9360,N_9772);
nand U10755 (N_10755,N_9177,N_9067);
or U10756 (N_10756,N_9671,N_9464);
nand U10757 (N_10757,N_10482,N_9329);
nor U10758 (N_10758,N_9549,N_10200);
nand U10759 (N_10759,N_10253,N_9164);
and U10760 (N_10760,N_9492,N_9930);
nand U10761 (N_10761,N_9282,N_9528);
nor U10762 (N_10762,N_9452,N_10069);
and U10763 (N_10763,N_9594,N_9059);
and U10764 (N_10764,N_9301,N_9356);
nand U10765 (N_10765,N_10280,N_9576);
nand U10766 (N_10766,N_9525,N_9349);
nand U10767 (N_10767,N_10468,N_9369);
nand U10768 (N_10768,N_9683,N_10108);
nand U10769 (N_10769,N_10134,N_10435);
or U10770 (N_10770,N_9420,N_9063);
nor U10771 (N_10771,N_9368,N_9065);
or U10772 (N_10772,N_10021,N_9285);
and U10773 (N_10773,N_10165,N_9134);
nor U10774 (N_10774,N_9516,N_9714);
nor U10775 (N_10775,N_10484,N_10260);
nor U10776 (N_10776,N_10363,N_10142);
nor U10777 (N_10777,N_9774,N_9345);
or U10778 (N_10778,N_9250,N_9704);
xor U10779 (N_10779,N_9531,N_10162);
nor U10780 (N_10780,N_9562,N_9650);
nand U10781 (N_10781,N_9564,N_9035);
nand U10782 (N_10782,N_9348,N_9278);
nor U10783 (N_10783,N_9960,N_9289);
and U10784 (N_10784,N_9432,N_10276);
xor U10785 (N_10785,N_10110,N_10248);
nor U10786 (N_10786,N_9532,N_10475);
nor U10787 (N_10787,N_9533,N_10138);
nand U10788 (N_10788,N_9858,N_9083);
or U10789 (N_10789,N_10308,N_10393);
nor U10790 (N_10790,N_9262,N_9405);
and U10791 (N_10791,N_10088,N_9022);
nor U10792 (N_10792,N_10316,N_10148);
or U10793 (N_10793,N_10008,N_10086);
xor U10794 (N_10794,N_9332,N_9154);
nand U10795 (N_10795,N_9221,N_9201);
nand U10796 (N_10796,N_9727,N_9018);
or U10797 (N_10797,N_10497,N_9124);
nand U10798 (N_10798,N_10489,N_9449);
and U10799 (N_10799,N_9937,N_10399);
nor U10800 (N_10800,N_10122,N_9383);
nor U10801 (N_10801,N_9192,N_9205);
nor U10802 (N_10802,N_9880,N_9621);
nor U10803 (N_10803,N_10047,N_9927);
or U10804 (N_10804,N_9309,N_9508);
or U10805 (N_10805,N_10242,N_10373);
nand U10806 (N_10806,N_9103,N_9280);
nor U10807 (N_10807,N_9084,N_9515);
nor U10808 (N_10808,N_9416,N_10346);
and U10809 (N_10809,N_9988,N_10492);
nand U10810 (N_10810,N_10034,N_9475);
and U10811 (N_10811,N_9815,N_10329);
and U10812 (N_10812,N_9653,N_10235);
nand U10813 (N_10813,N_9327,N_9455);
nor U10814 (N_10814,N_9370,N_9908);
nor U10815 (N_10815,N_9570,N_9599);
nand U10816 (N_10816,N_10463,N_10112);
nor U10817 (N_10817,N_9374,N_9945);
xnor U10818 (N_10818,N_9172,N_9976);
nand U10819 (N_10819,N_10469,N_9111);
or U10820 (N_10820,N_10204,N_10430);
nor U10821 (N_10821,N_9135,N_9434);
and U10822 (N_10822,N_9875,N_10013);
nor U10823 (N_10823,N_9292,N_9086);
nor U10824 (N_10824,N_9087,N_9584);
nor U10825 (N_10825,N_9778,N_10045);
or U10826 (N_10826,N_9050,N_9470);
and U10827 (N_10827,N_10187,N_9797);
nor U10828 (N_10828,N_9439,N_9619);
nor U10829 (N_10829,N_10472,N_10068);
or U10830 (N_10830,N_9631,N_9382);
or U10831 (N_10831,N_9835,N_9633);
nand U10832 (N_10832,N_10231,N_9330);
and U10833 (N_10833,N_9146,N_9979);
nor U10834 (N_10834,N_9597,N_10084);
nand U10835 (N_10835,N_10063,N_10306);
or U10836 (N_10836,N_10216,N_9555);
nor U10837 (N_10837,N_10062,N_10300);
xor U10838 (N_10838,N_9148,N_10291);
xor U10839 (N_10839,N_10194,N_9912);
xor U10840 (N_10840,N_9009,N_9933);
and U10841 (N_10841,N_9156,N_10037);
and U10842 (N_10842,N_9821,N_9034);
nor U10843 (N_10843,N_9446,N_9373);
nor U10844 (N_10844,N_10285,N_9685);
or U10845 (N_10845,N_10040,N_9958);
or U10846 (N_10846,N_10039,N_10072);
and U10847 (N_10847,N_9998,N_9642);
nor U10848 (N_10848,N_9493,N_9413);
nor U10849 (N_10849,N_10129,N_9426);
nand U10850 (N_10850,N_9581,N_9870);
or U10851 (N_10851,N_9228,N_9312);
nor U10852 (N_10852,N_9873,N_10364);
nor U10853 (N_10853,N_10206,N_10031);
and U10854 (N_10854,N_9728,N_9845);
and U10855 (N_10855,N_9252,N_10049);
nor U10856 (N_10856,N_10349,N_9074);
or U10857 (N_10857,N_10119,N_9923);
xnor U10858 (N_10858,N_9918,N_9765);
xnor U10859 (N_10859,N_9715,N_10168);
and U10860 (N_10860,N_10133,N_9286);
nor U10861 (N_10861,N_10441,N_9149);
or U10862 (N_10862,N_9456,N_9011);
nor U10863 (N_10863,N_9697,N_9089);
or U10864 (N_10864,N_10309,N_10085);
and U10865 (N_10865,N_9705,N_9114);
and U10866 (N_10866,N_10262,N_9853);
nand U10867 (N_10867,N_10017,N_10064);
nand U10868 (N_10868,N_9407,N_10178);
xnor U10869 (N_10869,N_9390,N_9072);
and U10870 (N_10870,N_9365,N_10096);
or U10871 (N_10871,N_9986,N_9741);
nor U10872 (N_10872,N_10385,N_9477);
nor U10873 (N_10873,N_10420,N_9820);
xor U10874 (N_10874,N_9414,N_10117);
xnor U10875 (N_10875,N_9760,N_9969);
xnor U10876 (N_10876,N_10302,N_9573);
nand U10877 (N_10877,N_9268,N_10228);
or U10878 (N_10878,N_9342,N_9110);
nand U10879 (N_10879,N_9551,N_9522);
and U10880 (N_10880,N_9939,N_10249);
or U10881 (N_10881,N_9045,N_10359);
and U10882 (N_10882,N_9218,N_9049);
nor U10883 (N_10883,N_9101,N_10189);
and U10884 (N_10884,N_10416,N_10471);
or U10885 (N_10885,N_9654,N_9260);
or U10886 (N_10886,N_10335,N_10082);
and U10887 (N_10887,N_9272,N_9947);
or U10888 (N_10888,N_9572,N_10191);
xor U10889 (N_10889,N_10394,N_9096);
or U10890 (N_10890,N_9304,N_9859);
or U10891 (N_10891,N_10361,N_9894);
nor U10892 (N_10892,N_10432,N_9659);
and U10893 (N_10893,N_10023,N_9082);
nand U10894 (N_10894,N_10226,N_9802);
nand U10895 (N_10895,N_9323,N_10257);
nand U10896 (N_10896,N_9122,N_10002);
or U10897 (N_10897,N_10058,N_9080);
nor U10898 (N_10898,N_9550,N_9466);
and U10899 (N_10899,N_9176,N_10245);
or U10900 (N_10900,N_9899,N_9433);
and U10901 (N_10901,N_9967,N_9589);
or U10902 (N_10902,N_10486,N_10311);
nand U10903 (N_10903,N_9320,N_9441);
or U10904 (N_10904,N_9916,N_10392);
xnor U10905 (N_10905,N_9232,N_9264);
nand U10906 (N_10906,N_9995,N_9486);
and U10907 (N_10907,N_10255,N_10011);
xnor U10908 (N_10908,N_9523,N_10080);
nand U10909 (N_10909,N_9975,N_9828);
and U10910 (N_10910,N_9603,N_10018);
xnor U10911 (N_10911,N_10070,N_9478);
or U10912 (N_10912,N_10333,N_10073);
and U10913 (N_10913,N_9150,N_10342);
nor U10914 (N_10914,N_9887,N_9521);
and U10915 (N_10915,N_10210,N_9534);
nand U10916 (N_10916,N_9852,N_10077);
and U10917 (N_10917,N_9761,N_9724);
nor U10918 (N_10918,N_9746,N_9436);
nor U10919 (N_10919,N_10446,N_9748);
nor U10920 (N_10920,N_9679,N_9577);
or U10921 (N_10921,N_9601,N_10312);
nor U10922 (N_10922,N_9130,N_9253);
nor U10923 (N_10923,N_9425,N_10273);
nand U10924 (N_10924,N_10443,N_10177);
and U10925 (N_10925,N_9652,N_10078);
nand U10926 (N_10926,N_9906,N_9409);
or U10927 (N_10927,N_10400,N_9326);
nor U10928 (N_10928,N_9372,N_9538);
nor U10929 (N_10929,N_10431,N_9759);
or U10930 (N_10930,N_9806,N_9602);
or U10931 (N_10931,N_9152,N_9398);
and U10932 (N_10932,N_9202,N_9197);
nor U10933 (N_10933,N_10466,N_10149);
or U10934 (N_10934,N_10366,N_9565);
or U10935 (N_10935,N_9126,N_9479);
or U10936 (N_10936,N_9468,N_9222);
nand U10937 (N_10937,N_9041,N_10310);
or U10938 (N_10938,N_9175,N_9354);
nand U10939 (N_10939,N_9421,N_9822);
nor U10940 (N_10940,N_10195,N_10474);
and U10941 (N_10941,N_10184,N_9298);
xnor U10942 (N_10942,N_9010,N_10440);
or U10943 (N_10943,N_10286,N_9712);
nand U10944 (N_10944,N_9343,N_9006);
xnor U10945 (N_10945,N_9753,N_10131);
xnor U10946 (N_10946,N_9991,N_9071);
and U10947 (N_10947,N_9644,N_9037);
and U10948 (N_10948,N_9030,N_9890);
or U10949 (N_10949,N_9561,N_9437);
and U10950 (N_10950,N_10325,N_9314);
nor U10951 (N_10951,N_9698,N_9944);
and U10952 (N_10952,N_9284,N_9003);
or U10953 (N_10953,N_9145,N_9966);
xnor U10954 (N_10954,N_9953,N_9277);
and U10955 (N_10955,N_9347,N_10442);
xnor U10956 (N_10956,N_10263,N_9985);
nor U10957 (N_10957,N_9105,N_10404);
and U10958 (N_10958,N_9476,N_10459);
or U10959 (N_10959,N_10225,N_9955);
nor U10960 (N_10960,N_10217,N_9504);
and U10961 (N_10961,N_9957,N_10304);
nand U10962 (N_10962,N_9940,N_9739);
and U10963 (N_10963,N_10174,N_9596);
nand U10964 (N_10964,N_9108,N_10421);
nand U10965 (N_10965,N_9199,N_9837);
nand U10966 (N_10966,N_10453,N_9919);
xor U10967 (N_10967,N_9905,N_10220);
or U10968 (N_10968,N_9125,N_10268);
xnor U10969 (N_10969,N_10330,N_10410);
or U10970 (N_10970,N_10043,N_10101);
nand U10971 (N_10971,N_10387,N_9273);
and U10972 (N_10972,N_9921,N_9740);
nand U10973 (N_10973,N_9032,N_9780);
or U10974 (N_10974,N_10374,N_10015);
and U10975 (N_10975,N_9558,N_9617);
and U10976 (N_10976,N_9014,N_9796);
xor U10977 (N_10977,N_10267,N_9182);
nand U10978 (N_10978,N_10341,N_9106);
or U10979 (N_10979,N_9016,N_9274);
nand U10980 (N_10980,N_10019,N_9529);
or U10981 (N_10981,N_9812,N_9269);
and U10982 (N_10982,N_9524,N_10313);
and U10983 (N_10983,N_10115,N_10493);
xnor U10984 (N_10984,N_10089,N_9952);
and U10985 (N_10985,N_9884,N_9017);
or U10986 (N_10986,N_10275,N_9267);
and U10987 (N_10987,N_9341,N_9689);
or U10988 (N_10988,N_9400,N_10375);
nand U10989 (N_10989,N_9166,N_9293);
and U10990 (N_10990,N_10447,N_9585);
and U10991 (N_10991,N_9090,N_9959);
nor U10992 (N_10992,N_9100,N_9618);
nand U10993 (N_10993,N_10250,N_9102);
and U10994 (N_10994,N_9046,N_9023);
and U10995 (N_10995,N_9542,N_9000);
nor U10996 (N_10996,N_10369,N_10150);
and U10997 (N_10997,N_9539,N_10033);
nand U10998 (N_10998,N_9661,N_9411);
and U10999 (N_10999,N_10395,N_9226);
and U11000 (N_11000,N_10181,N_9706);
xor U11001 (N_11001,N_10357,N_10258);
and U11002 (N_11002,N_9586,N_10323);
or U11003 (N_11003,N_9480,N_9517);
and U11004 (N_11004,N_9647,N_10461);
and U11005 (N_11005,N_9984,N_9658);
and U11006 (N_11006,N_9823,N_9896);
nor U11007 (N_11007,N_9070,N_9604);
and U11008 (N_11008,N_9925,N_10488);
nor U11009 (N_11009,N_9878,N_9396);
and U11010 (N_11010,N_9545,N_10433);
nand U11011 (N_11011,N_9061,N_9681);
nand U11012 (N_11012,N_9687,N_10010);
and U11013 (N_11013,N_10389,N_10143);
or U11014 (N_11014,N_9737,N_10173);
nor U11015 (N_11015,N_9841,N_9962);
nand U11016 (N_11016,N_9217,N_9546);
nor U11017 (N_11017,N_10029,N_9600);
xnor U11018 (N_11018,N_9632,N_9132);
nor U11019 (N_11019,N_9605,N_10157);
xnor U11020 (N_11020,N_10005,N_10411);
nand U11021 (N_11021,N_9913,N_10383);
and U11022 (N_11022,N_10140,N_9646);
nand U11023 (N_11023,N_9151,N_9718);
and U11024 (N_11024,N_10203,N_9615);
nand U11025 (N_11025,N_9098,N_9511);
nand U11026 (N_11026,N_9868,N_10102);
xnor U11027 (N_11027,N_9118,N_9225);
and U11028 (N_11028,N_9143,N_9180);
xor U11029 (N_11029,N_9194,N_9954);
and U11030 (N_11030,N_10074,N_9394);
and U11031 (N_11031,N_9387,N_9247);
and U11032 (N_11032,N_9613,N_9085);
nor U11033 (N_11033,N_9540,N_10166);
nor U11034 (N_11034,N_9404,N_9190);
nor U11035 (N_11035,N_9113,N_9708);
xor U11036 (N_11036,N_10146,N_9461);
nor U11037 (N_11037,N_10487,N_9770);
and U11038 (N_11038,N_10496,N_9951);
and U11039 (N_11039,N_9167,N_9686);
and U11040 (N_11040,N_9779,N_9709);
and U11041 (N_11041,N_10436,N_10347);
and U11042 (N_11042,N_9931,N_9567);
nand U11043 (N_11043,N_9307,N_10458);
nor U11044 (N_11044,N_10121,N_9198);
nand U11045 (N_11045,N_10339,N_10318);
and U11046 (N_11046,N_10388,N_9622);
xor U11047 (N_11047,N_9808,N_9819);
or U11048 (N_11048,N_10237,N_9355);
or U11049 (N_11049,N_10289,N_10083);
and U11050 (N_11050,N_10467,N_10386);
nand U11051 (N_11051,N_9231,N_10294);
or U11052 (N_11052,N_9643,N_9471);
nand U11053 (N_11053,N_9503,N_10104);
and U11054 (N_11054,N_9047,N_10186);
nand U11055 (N_11055,N_10417,N_9509);
and U11056 (N_11056,N_9694,N_9961);
and U11057 (N_11057,N_9453,N_10030);
xnor U11058 (N_11058,N_9804,N_9872);
xor U11059 (N_11059,N_9340,N_10046);
and U11060 (N_11060,N_9185,N_10182);
and U11061 (N_11061,N_10214,N_10014);
nand U11062 (N_11062,N_9743,N_9651);
nor U11063 (N_11063,N_9692,N_9212);
nor U11064 (N_11064,N_10384,N_9447);
nor U11065 (N_11065,N_10380,N_9331);
or U11066 (N_11066,N_9805,N_10205);
or U11067 (N_11067,N_10055,N_10370);
or U11068 (N_11068,N_10328,N_9506);
and U11069 (N_11069,N_9403,N_9069);
nor U11070 (N_11070,N_10283,N_10456);
or U11071 (N_11071,N_9408,N_9364);
nor U11072 (N_11072,N_9733,N_10298);
nor U11073 (N_11073,N_9263,N_10391);
nor U11074 (N_11074,N_9982,N_9240);
and U11075 (N_11075,N_9335,N_9224);
and U11076 (N_11076,N_9339,N_9575);
or U11077 (N_11077,N_10415,N_9855);
nor U11078 (N_11078,N_9857,N_10438);
nor U11079 (N_11079,N_9078,N_10038);
or U11080 (N_11080,N_9241,N_9813);
or U11081 (N_11081,N_10222,N_9568);
nor U11082 (N_11082,N_10271,N_9283);
or U11083 (N_11083,N_9590,N_9556);
nor U11084 (N_11084,N_9914,N_9829);
nor U11085 (N_11085,N_9265,N_9385);
and U11086 (N_11086,N_9690,N_9656);
or U11087 (N_11087,N_10450,N_10026);
nand U11088 (N_11088,N_10305,N_10127);
nor U11089 (N_11089,N_9902,N_9782);
nor U11090 (N_11090,N_10281,N_9310);
or U11091 (N_11091,N_10490,N_9160);
nand U11092 (N_11092,N_10270,N_9058);
nor U11093 (N_11093,N_9321,N_9800);
or U11094 (N_11094,N_10402,N_9981);
nor U11095 (N_11095,N_9612,N_9676);
or U11096 (N_11096,N_9882,N_9624);
nor U11097 (N_11097,N_9499,N_9395);
nor U11098 (N_11098,N_9662,N_9762);
nor U11099 (N_11099,N_9211,N_9465);
or U11100 (N_11100,N_10477,N_9854);
and U11101 (N_11101,N_9593,N_10367);
and U11102 (N_11102,N_9317,N_10223);
and U11103 (N_11103,N_9144,N_9611);
nand U11104 (N_11104,N_9569,N_10378);
and U11105 (N_11105,N_9497,N_10060);
or U11106 (N_11106,N_9406,N_9027);
nand U11107 (N_11107,N_9093,N_9710);
or U11108 (N_11108,N_10185,N_9987);
or U11109 (N_11109,N_9129,N_9758);
nand U11110 (N_11110,N_9002,N_10201);
or U11111 (N_11111,N_10422,N_9186);
and U11112 (N_11112,N_10114,N_10230);
nand U11113 (N_11113,N_9248,N_9831);
or U11114 (N_11114,N_9973,N_9353);
and U11115 (N_11115,N_9300,N_10213);
or U11116 (N_11116,N_10481,N_10243);
nand U11117 (N_11117,N_10042,N_10180);
or U11118 (N_11118,N_10051,N_9121);
xnor U11119 (N_11119,N_10169,N_9816);
or U11120 (N_11120,N_10059,N_9422);
nor U11121 (N_11121,N_9763,N_9351);
or U11122 (N_11122,N_10109,N_10224);
nor U11123 (N_11123,N_10338,N_9942);
nor U11124 (N_11124,N_9789,N_9609);
nand U11125 (N_11125,N_10272,N_9157);
or U11126 (N_11126,N_9196,N_9031);
xor U11127 (N_11127,N_9935,N_9359);
or U11128 (N_11128,N_9754,N_10052);
nor U11129 (N_11129,N_10455,N_10097);
xor U11130 (N_11130,N_10161,N_9423);
nand U11131 (N_11131,N_9161,N_9489);
xnor U11132 (N_11132,N_10320,N_10473);
or U11133 (N_11133,N_10499,N_9749);
xor U11134 (N_11134,N_9482,N_10334);
or U11135 (N_11135,N_10414,N_9092);
nand U11136 (N_11136,N_9766,N_9992);
nand U11137 (N_11137,N_9793,N_9350);
or U11138 (N_11138,N_9431,N_10485);
and U11139 (N_11139,N_10065,N_9191);
or U11140 (N_11140,N_10337,N_9249);
or U11141 (N_11141,N_9021,N_10292);
or U11142 (N_11142,N_10355,N_9675);
nor U11143 (N_11143,N_9246,N_9206);
and U11144 (N_11144,N_9862,N_10107);
or U11145 (N_11145,N_10076,N_10470);
or U11146 (N_11146,N_9163,N_9680);
nand U11147 (N_11147,N_9978,N_9417);
nor U11148 (N_11148,N_9494,N_9220);
or U11149 (N_11149,N_9843,N_9502);
or U11150 (N_11150,N_9048,N_9444);
and U11151 (N_11151,N_9791,N_10006);
nor U11152 (N_11152,N_10075,N_10362);
nor U11153 (N_11153,N_9752,N_9826);
xor U11154 (N_11154,N_9608,N_10007);
nand U11155 (N_11155,N_9648,N_9418);
nor U11156 (N_11156,N_9895,N_10095);
xnor U11157 (N_11157,N_10238,N_9242);
or U11158 (N_11158,N_9291,N_9598);
and U11159 (N_11159,N_10054,N_10457);
and U11160 (N_11160,N_9064,N_9375);
nand U11161 (N_11161,N_9790,N_9443);
or U11162 (N_11162,N_9963,N_9019);
nor U11163 (N_11163,N_9968,N_9213);
nand U11164 (N_11164,N_9924,N_10397);
and U11165 (N_11165,N_9717,N_9863);
or U11166 (N_11166,N_9155,N_9203);
and U11167 (N_11167,N_9934,N_9518);
and U11168 (N_11168,N_9153,N_10406);
and U11169 (N_11169,N_10314,N_9183);
and U11170 (N_11170,N_9458,N_9626);
xnor U11171 (N_11171,N_9008,N_9537);
nor U11172 (N_11172,N_9920,N_9442);
xor U11173 (N_11173,N_9510,N_10279);
or U11174 (N_11174,N_9844,N_9338);
nand U11175 (N_11175,N_9707,N_9964);
xor U11176 (N_11176,N_9784,N_9856);
nand U11177 (N_11177,N_9123,N_9560);
nand U11178 (N_11178,N_9926,N_10354);
nor U11179 (N_11179,N_10264,N_10003);
and U11180 (N_11180,N_10498,N_10427);
nand U11181 (N_11181,N_9711,N_10356);
and U11182 (N_11182,N_9487,N_10296);
nand U11183 (N_11183,N_9076,N_10403);
nor U11184 (N_11184,N_9007,N_9592);
and U11185 (N_11185,N_10144,N_9825);
nand U11186 (N_11186,N_9484,N_9131);
nor U11187 (N_11187,N_9138,N_9583);
or U11188 (N_11188,N_9235,N_9900);
xor U11189 (N_11189,N_9827,N_9897);
and U11190 (N_11190,N_10188,N_9541);
and U11191 (N_11191,N_9376,N_9757);
nand U11192 (N_11192,N_9773,N_9188);
nand U11193 (N_11193,N_9462,N_9547);
or U11194 (N_11194,N_9302,N_9830);
or U11195 (N_11195,N_9554,N_9670);
nand U11196 (N_11196,N_9889,N_10345);
nor U11197 (N_11197,N_10000,N_10429);
and U11198 (N_11198,N_10444,N_10027);
nand U11199 (N_11199,N_9362,N_9088);
or U11200 (N_11200,N_10413,N_9663);
or U11201 (N_11201,N_9029,N_10241);
and U11202 (N_11202,N_9077,N_10153);
or U11203 (N_11203,N_9313,N_9181);
nand U11204 (N_11204,N_9366,N_9836);
xnor U11205 (N_11205,N_9168,N_10004);
or U11206 (N_11206,N_9860,N_10207);
nand U11207 (N_11207,N_9116,N_10491);
nor U11208 (N_11208,N_10372,N_9410);
nand U11209 (N_11209,N_9140,N_10412);
and U11210 (N_11210,N_10327,N_9251);
or U11211 (N_11211,N_10116,N_9756);
nor U11212 (N_11212,N_10020,N_9322);
xnor U11213 (N_11213,N_9713,N_9764);
nor U11214 (N_11214,N_10061,N_10437);
nor U11215 (N_11215,N_10103,N_9162);
and U11216 (N_11216,N_9783,N_10495);
and U11217 (N_11217,N_10396,N_10376);
or U11218 (N_11218,N_10266,N_9473);
and U11219 (N_11219,N_9490,N_9361);
and U11220 (N_11220,N_10167,N_9039);
and U11221 (N_11221,N_10448,N_10398);
nor U11222 (N_11222,N_9223,N_10215);
and U11223 (N_11223,N_9428,N_10036);
or U11224 (N_11224,N_10056,N_9655);
nor U11225 (N_11225,N_9814,N_9054);
nor U11226 (N_11226,N_10172,N_10001);
nand U11227 (N_11227,N_10123,N_10407);
nor U11228 (N_11228,N_9481,N_9169);
and U11229 (N_11229,N_9657,N_9950);
or U11230 (N_11230,N_10208,N_10053);
nand U11231 (N_11231,N_9970,N_9911);
nand U11232 (N_11232,N_9474,N_9834);
nor U11233 (N_11233,N_9257,N_9459);
and U11234 (N_11234,N_10022,N_10240);
and U11235 (N_11235,N_9244,N_10106);
nand U11236 (N_11236,N_10336,N_10303);
nor U11237 (N_11237,N_9363,N_10269);
xor U11238 (N_11238,N_9097,N_9917);
nand U11239 (N_11239,N_9607,N_9566);
or U11240 (N_11240,N_9501,N_9012);
xor U11241 (N_11241,N_9159,N_9977);
nor U11242 (N_11242,N_9238,N_9795);
or U11243 (N_11243,N_9750,N_9907);
nand U11244 (N_11244,N_9337,N_9388);
nand U11245 (N_11245,N_10111,N_9848);
nand U11246 (N_11246,N_10352,N_10233);
and U11247 (N_11247,N_9775,N_10147);
xnor U11248 (N_11248,N_9079,N_10190);
nand U11249 (N_11249,N_10278,N_9334);
or U11250 (N_11250,N_10232,N_9974);
and U11251 (N_11251,N_9888,N_9934);
and U11252 (N_11252,N_9113,N_9537);
nor U11253 (N_11253,N_9967,N_10405);
nor U11254 (N_11254,N_10060,N_10446);
nand U11255 (N_11255,N_10274,N_10261);
or U11256 (N_11256,N_9512,N_10227);
nor U11257 (N_11257,N_9061,N_9555);
xnor U11258 (N_11258,N_9518,N_9848);
and U11259 (N_11259,N_10303,N_9180);
or U11260 (N_11260,N_9474,N_9911);
nor U11261 (N_11261,N_9539,N_9491);
and U11262 (N_11262,N_9499,N_10267);
nor U11263 (N_11263,N_10113,N_10423);
nand U11264 (N_11264,N_10424,N_10435);
nor U11265 (N_11265,N_9632,N_10126);
and U11266 (N_11266,N_9793,N_9185);
xnor U11267 (N_11267,N_9959,N_9884);
or U11268 (N_11268,N_10041,N_9924);
nand U11269 (N_11269,N_9797,N_10324);
or U11270 (N_11270,N_9274,N_9772);
or U11271 (N_11271,N_9601,N_9517);
xor U11272 (N_11272,N_10153,N_9132);
nor U11273 (N_11273,N_9605,N_9488);
or U11274 (N_11274,N_9414,N_9609);
nand U11275 (N_11275,N_9642,N_9664);
nor U11276 (N_11276,N_10075,N_10009);
nor U11277 (N_11277,N_9086,N_9047);
nand U11278 (N_11278,N_9539,N_10097);
or U11279 (N_11279,N_10450,N_10099);
nand U11280 (N_11280,N_9273,N_9834);
nand U11281 (N_11281,N_10433,N_9232);
nand U11282 (N_11282,N_9420,N_10461);
nand U11283 (N_11283,N_9745,N_10180);
or U11284 (N_11284,N_10465,N_9710);
and U11285 (N_11285,N_10283,N_9422);
nand U11286 (N_11286,N_9043,N_9350);
nand U11287 (N_11287,N_10453,N_10487);
xor U11288 (N_11288,N_10219,N_10296);
and U11289 (N_11289,N_10219,N_9067);
and U11290 (N_11290,N_9028,N_10264);
nand U11291 (N_11291,N_9526,N_10365);
xor U11292 (N_11292,N_10365,N_9165);
nor U11293 (N_11293,N_9339,N_10338);
xor U11294 (N_11294,N_9815,N_10216);
or U11295 (N_11295,N_9317,N_10446);
nand U11296 (N_11296,N_9109,N_10365);
nor U11297 (N_11297,N_9383,N_9357);
nor U11298 (N_11298,N_10281,N_9409);
or U11299 (N_11299,N_9947,N_10037);
or U11300 (N_11300,N_9517,N_10104);
nand U11301 (N_11301,N_10422,N_9809);
nand U11302 (N_11302,N_9211,N_10086);
or U11303 (N_11303,N_9726,N_9623);
or U11304 (N_11304,N_9336,N_9027);
or U11305 (N_11305,N_9097,N_9501);
nor U11306 (N_11306,N_10052,N_9538);
nor U11307 (N_11307,N_9131,N_9765);
nand U11308 (N_11308,N_9027,N_9435);
nor U11309 (N_11309,N_9701,N_9014);
nor U11310 (N_11310,N_9003,N_9155);
and U11311 (N_11311,N_10013,N_10273);
nor U11312 (N_11312,N_10074,N_10454);
xnor U11313 (N_11313,N_9603,N_10219);
xnor U11314 (N_11314,N_9784,N_9808);
or U11315 (N_11315,N_10233,N_9861);
nor U11316 (N_11316,N_9910,N_10254);
and U11317 (N_11317,N_9271,N_9202);
nor U11318 (N_11318,N_10295,N_10421);
nor U11319 (N_11319,N_9923,N_9372);
nor U11320 (N_11320,N_10030,N_10377);
and U11321 (N_11321,N_9791,N_9506);
and U11322 (N_11322,N_9440,N_9541);
and U11323 (N_11323,N_9960,N_10062);
or U11324 (N_11324,N_10137,N_9525);
and U11325 (N_11325,N_10480,N_9444);
nand U11326 (N_11326,N_10446,N_9746);
and U11327 (N_11327,N_9466,N_10366);
or U11328 (N_11328,N_10098,N_9170);
nand U11329 (N_11329,N_10077,N_10458);
nor U11330 (N_11330,N_9036,N_9853);
or U11331 (N_11331,N_10030,N_10211);
xor U11332 (N_11332,N_9956,N_9436);
nand U11333 (N_11333,N_9784,N_9766);
nor U11334 (N_11334,N_9470,N_9258);
or U11335 (N_11335,N_9130,N_9584);
or U11336 (N_11336,N_10248,N_9942);
and U11337 (N_11337,N_10081,N_9557);
nor U11338 (N_11338,N_9820,N_9504);
nor U11339 (N_11339,N_9126,N_10263);
nor U11340 (N_11340,N_10429,N_9168);
nand U11341 (N_11341,N_10057,N_9603);
and U11342 (N_11342,N_9832,N_9426);
or U11343 (N_11343,N_10485,N_9878);
and U11344 (N_11344,N_9100,N_9657);
nand U11345 (N_11345,N_9759,N_10030);
or U11346 (N_11346,N_10231,N_9056);
and U11347 (N_11347,N_9608,N_9362);
nand U11348 (N_11348,N_10112,N_9126);
or U11349 (N_11349,N_10280,N_10217);
nor U11350 (N_11350,N_10151,N_9162);
or U11351 (N_11351,N_9097,N_9127);
nor U11352 (N_11352,N_10083,N_9539);
nor U11353 (N_11353,N_9751,N_9982);
xor U11354 (N_11354,N_10317,N_10470);
xor U11355 (N_11355,N_10482,N_10186);
nor U11356 (N_11356,N_9609,N_10336);
or U11357 (N_11357,N_10136,N_10397);
nor U11358 (N_11358,N_9042,N_10312);
and U11359 (N_11359,N_9190,N_9588);
nor U11360 (N_11360,N_10144,N_9619);
nand U11361 (N_11361,N_10151,N_9394);
nand U11362 (N_11362,N_9222,N_10254);
or U11363 (N_11363,N_10453,N_10043);
and U11364 (N_11364,N_9305,N_9006);
and U11365 (N_11365,N_9534,N_9066);
xor U11366 (N_11366,N_10438,N_9641);
and U11367 (N_11367,N_9435,N_9911);
xnor U11368 (N_11368,N_10352,N_10359);
and U11369 (N_11369,N_9543,N_10201);
or U11370 (N_11370,N_9403,N_10061);
nand U11371 (N_11371,N_9897,N_9527);
nand U11372 (N_11372,N_9643,N_10440);
nor U11373 (N_11373,N_9091,N_9595);
and U11374 (N_11374,N_10243,N_9734);
xor U11375 (N_11375,N_9628,N_9547);
nand U11376 (N_11376,N_10217,N_9636);
or U11377 (N_11377,N_9560,N_10196);
and U11378 (N_11378,N_9537,N_9960);
nand U11379 (N_11379,N_10292,N_9012);
nor U11380 (N_11380,N_9426,N_9351);
or U11381 (N_11381,N_9179,N_9661);
and U11382 (N_11382,N_10348,N_10376);
nand U11383 (N_11383,N_9916,N_10022);
nor U11384 (N_11384,N_9753,N_9664);
nand U11385 (N_11385,N_10115,N_9978);
nand U11386 (N_11386,N_9120,N_9749);
or U11387 (N_11387,N_9838,N_9623);
and U11388 (N_11388,N_9899,N_10433);
or U11389 (N_11389,N_9702,N_10384);
and U11390 (N_11390,N_9932,N_9030);
or U11391 (N_11391,N_9333,N_9799);
and U11392 (N_11392,N_9691,N_9854);
and U11393 (N_11393,N_10498,N_9741);
and U11394 (N_11394,N_9413,N_9253);
nor U11395 (N_11395,N_9553,N_9660);
xor U11396 (N_11396,N_10495,N_9189);
nand U11397 (N_11397,N_10109,N_9035);
or U11398 (N_11398,N_9098,N_10056);
or U11399 (N_11399,N_10183,N_9185);
or U11400 (N_11400,N_9708,N_9601);
xnor U11401 (N_11401,N_9831,N_10102);
nor U11402 (N_11402,N_9327,N_9095);
and U11403 (N_11403,N_10033,N_9317);
nor U11404 (N_11404,N_10155,N_9784);
nand U11405 (N_11405,N_10466,N_9027);
nand U11406 (N_11406,N_10168,N_9482);
nand U11407 (N_11407,N_9639,N_9610);
and U11408 (N_11408,N_10469,N_10145);
nor U11409 (N_11409,N_9508,N_9111);
nand U11410 (N_11410,N_9930,N_9830);
nand U11411 (N_11411,N_9759,N_9259);
xnor U11412 (N_11412,N_10374,N_10139);
nor U11413 (N_11413,N_9807,N_9602);
or U11414 (N_11414,N_10228,N_10330);
nor U11415 (N_11415,N_9297,N_10356);
nand U11416 (N_11416,N_9726,N_10402);
xor U11417 (N_11417,N_9459,N_10040);
nor U11418 (N_11418,N_9134,N_9493);
and U11419 (N_11419,N_10249,N_9309);
and U11420 (N_11420,N_9304,N_9193);
nand U11421 (N_11421,N_9537,N_9816);
nor U11422 (N_11422,N_9586,N_10196);
and U11423 (N_11423,N_9905,N_9022);
nand U11424 (N_11424,N_9375,N_9239);
nand U11425 (N_11425,N_9706,N_10021);
nor U11426 (N_11426,N_9982,N_9698);
and U11427 (N_11427,N_9777,N_10368);
nor U11428 (N_11428,N_10324,N_9659);
nor U11429 (N_11429,N_9901,N_9760);
nand U11430 (N_11430,N_9816,N_9989);
nand U11431 (N_11431,N_10199,N_9439);
nand U11432 (N_11432,N_10405,N_9451);
and U11433 (N_11433,N_10026,N_9224);
or U11434 (N_11434,N_9428,N_10019);
and U11435 (N_11435,N_9441,N_9461);
nor U11436 (N_11436,N_9131,N_9574);
nor U11437 (N_11437,N_10273,N_10316);
xor U11438 (N_11438,N_9708,N_9722);
or U11439 (N_11439,N_10382,N_9525);
and U11440 (N_11440,N_9780,N_9051);
or U11441 (N_11441,N_9538,N_9807);
or U11442 (N_11442,N_10162,N_10253);
nor U11443 (N_11443,N_9149,N_9014);
nor U11444 (N_11444,N_9854,N_10311);
nand U11445 (N_11445,N_9961,N_9272);
or U11446 (N_11446,N_10370,N_10027);
or U11447 (N_11447,N_9476,N_9600);
and U11448 (N_11448,N_9569,N_9400);
and U11449 (N_11449,N_9189,N_9872);
nand U11450 (N_11450,N_9548,N_9379);
nand U11451 (N_11451,N_10209,N_9657);
and U11452 (N_11452,N_9125,N_10123);
nand U11453 (N_11453,N_9622,N_9201);
and U11454 (N_11454,N_10247,N_9852);
nand U11455 (N_11455,N_9440,N_9556);
nor U11456 (N_11456,N_9911,N_9350);
nor U11457 (N_11457,N_9685,N_9285);
xor U11458 (N_11458,N_10443,N_9207);
and U11459 (N_11459,N_9216,N_10266);
nand U11460 (N_11460,N_10043,N_9367);
nand U11461 (N_11461,N_9437,N_9672);
and U11462 (N_11462,N_9418,N_9371);
nand U11463 (N_11463,N_10386,N_9219);
or U11464 (N_11464,N_10327,N_9919);
nor U11465 (N_11465,N_9912,N_9369);
or U11466 (N_11466,N_9149,N_9078);
or U11467 (N_11467,N_9529,N_10299);
nand U11468 (N_11468,N_9858,N_9399);
nor U11469 (N_11469,N_9105,N_9263);
nor U11470 (N_11470,N_9105,N_9372);
nor U11471 (N_11471,N_9459,N_9796);
nor U11472 (N_11472,N_9523,N_10162);
nand U11473 (N_11473,N_9519,N_9260);
or U11474 (N_11474,N_9585,N_9431);
and U11475 (N_11475,N_9263,N_9761);
nor U11476 (N_11476,N_9907,N_9634);
or U11477 (N_11477,N_9887,N_9938);
nand U11478 (N_11478,N_9759,N_9736);
nand U11479 (N_11479,N_9899,N_10170);
or U11480 (N_11480,N_9670,N_10315);
and U11481 (N_11481,N_10155,N_9868);
nand U11482 (N_11482,N_9070,N_10116);
nor U11483 (N_11483,N_9911,N_9898);
and U11484 (N_11484,N_9566,N_10273);
nand U11485 (N_11485,N_10105,N_9439);
nand U11486 (N_11486,N_9350,N_10255);
nor U11487 (N_11487,N_9066,N_9743);
nor U11488 (N_11488,N_9228,N_9008);
nand U11489 (N_11489,N_9024,N_9229);
and U11490 (N_11490,N_9519,N_9840);
and U11491 (N_11491,N_9327,N_10151);
xor U11492 (N_11492,N_9939,N_9300);
or U11493 (N_11493,N_9480,N_9125);
xnor U11494 (N_11494,N_9287,N_9939);
xor U11495 (N_11495,N_10151,N_9108);
or U11496 (N_11496,N_9625,N_9715);
xnor U11497 (N_11497,N_9940,N_9427);
or U11498 (N_11498,N_9196,N_9436);
or U11499 (N_11499,N_10298,N_9452);
and U11500 (N_11500,N_9493,N_9902);
xnor U11501 (N_11501,N_9663,N_9642);
nand U11502 (N_11502,N_10108,N_10383);
and U11503 (N_11503,N_9140,N_9186);
or U11504 (N_11504,N_9353,N_9412);
nand U11505 (N_11505,N_10362,N_9673);
xnor U11506 (N_11506,N_9085,N_9565);
nor U11507 (N_11507,N_10399,N_9742);
nand U11508 (N_11508,N_10077,N_9399);
nand U11509 (N_11509,N_10281,N_9927);
or U11510 (N_11510,N_9992,N_9333);
nor U11511 (N_11511,N_9195,N_9749);
nand U11512 (N_11512,N_10181,N_9909);
and U11513 (N_11513,N_9521,N_10495);
nor U11514 (N_11514,N_9585,N_10378);
nor U11515 (N_11515,N_9478,N_10216);
or U11516 (N_11516,N_9654,N_9697);
and U11517 (N_11517,N_9787,N_10025);
or U11518 (N_11518,N_9491,N_9907);
nor U11519 (N_11519,N_9137,N_9859);
and U11520 (N_11520,N_10100,N_10116);
and U11521 (N_11521,N_10333,N_9188);
and U11522 (N_11522,N_9531,N_9612);
nor U11523 (N_11523,N_10233,N_10115);
nand U11524 (N_11524,N_9773,N_9405);
and U11525 (N_11525,N_9098,N_9469);
and U11526 (N_11526,N_9500,N_9799);
nand U11527 (N_11527,N_9177,N_9203);
and U11528 (N_11528,N_9760,N_9514);
and U11529 (N_11529,N_9402,N_10467);
or U11530 (N_11530,N_9829,N_9550);
or U11531 (N_11531,N_9840,N_10346);
nor U11532 (N_11532,N_10271,N_9820);
and U11533 (N_11533,N_9654,N_10196);
nor U11534 (N_11534,N_9743,N_10377);
nand U11535 (N_11535,N_9256,N_9960);
xor U11536 (N_11536,N_10288,N_10044);
nor U11537 (N_11537,N_9685,N_9881);
or U11538 (N_11538,N_9131,N_10324);
nor U11539 (N_11539,N_9283,N_9318);
nand U11540 (N_11540,N_10459,N_9994);
nand U11541 (N_11541,N_9606,N_9605);
or U11542 (N_11542,N_10262,N_10236);
nor U11543 (N_11543,N_10225,N_9342);
and U11544 (N_11544,N_10439,N_9767);
xnor U11545 (N_11545,N_9148,N_9747);
or U11546 (N_11546,N_9519,N_10460);
nor U11547 (N_11547,N_10012,N_9535);
nor U11548 (N_11548,N_9474,N_10066);
nand U11549 (N_11549,N_9478,N_9633);
or U11550 (N_11550,N_9654,N_9200);
nor U11551 (N_11551,N_9895,N_10141);
nor U11552 (N_11552,N_9145,N_9457);
nor U11553 (N_11553,N_9825,N_9245);
or U11554 (N_11554,N_9165,N_10440);
and U11555 (N_11555,N_9592,N_9783);
nor U11556 (N_11556,N_10340,N_9305);
or U11557 (N_11557,N_9015,N_10133);
or U11558 (N_11558,N_10387,N_10094);
nand U11559 (N_11559,N_9619,N_9043);
or U11560 (N_11560,N_9423,N_10165);
xor U11561 (N_11561,N_9351,N_9522);
nand U11562 (N_11562,N_9524,N_9366);
nor U11563 (N_11563,N_10438,N_9582);
or U11564 (N_11564,N_9238,N_9427);
nor U11565 (N_11565,N_10478,N_9959);
nor U11566 (N_11566,N_9394,N_10042);
and U11567 (N_11567,N_9611,N_9097);
nor U11568 (N_11568,N_10383,N_9853);
nor U11569 (N_11569,N_9669,N_9956);
nor U11570 (N_11570,N_9826,N_9275);
nand U11571 (N_11571,N_9136,N_9142);
nand U11572 (N_11572,N_9864,N_9993);
or U11573 (N_11573,N_9280,N_10019);
or U11574 (N_11574,N_9014,N_10445);
nor U11575 (N_11575,N_10093,N_9714);
xnor U11576 (N_11576,N_9684,N_9708);
and U11577 (N_11577,N_9952,N_10273);
nand U11578 (N_11578,N_10217,N_9515);
nor U11579 (N_11579,N_9114,N_9463);
or U11580 (N_11580,N_9753,N_9839);
nor U11581 (N_11581,N_9830,N_9549);
nor U11582 (N_11582,N_9272,N_9919);
xor U11583 (N_11583,N_10032,N_10138);
nor U11584 (N_11584,N_10470,N_9022);
and U11585 (N_11585,N_9150,N_10012);
and U11586 (N_11586,N_9971,N_9148);
xnor U11587 (N_11587,N_9857,N_9172);
and U11588 (N_11588,N_9884,N_9302);
nand U11589 (N_11589,N_9436,N_10213);
xor U11590 (N_11590,N_9821,N_9790);
or U11591 (N_11591,N_9698,N_9556);
nand U11592 (N_11592,N_9524,N_10096);
xor U11593 (N_11593,N_10322,N_10247);
nor U11594 (N_11594,N_9654,N_9573);
nand U11595 (N_11595,N_10105,N_9003);
nor U11596 (N_11596,N_10079,N_9841);
nor U11597 (N_11597,N_9475,N_9865);
nor U11598 (N_11598,N_9487,N_9223);
or U11599 (N_11599,N_10496,N_10461);
or U11600 (N_11600,N_10153,N_9820);
nand U11601 (N_11601,N_9527,N_10387);
xor U11602 (N_11602,N_9968,N_9033);
and U11603 (N_11603,N_9841,N_9956);
or U11604 (N_11604,N_9585,N_9158);
nor U11605 (N_11605,N_10116,N_10102);
xnor U11606 (N_11606,N_9072,N_9559);
or U11607 (N_11607,N_9396,N_10191);
nand U11608 (N_11608,N_9545,N_9093);
nand U11609 (N_11609,N_10467,N_10497);
and U11610 (N_11610,N_9986,N_9043);
or U11611 (N_11611,N_9752,N_9640);
or U11612 (N_11612,N_9118,N_9952);
and U11613 (N_11613,N_9061,N_9235);
xnor U11614 (N_11614,N_9742,N_9142);
and U11615 (N_11615,N_9716,N_10424);
nand U11616 (N_11616,N_9560,N_10473);
nand U11617 (N_11617,N_9283,N_10296);
nor U11618 (N_11618,N_10464,N_9764);
and U11619 (N_11619,N_10442,N_10118);
and U11620 (N_11620,N_9505,N_10305);
and U11621 (N_11621,N_10288,N_10289);
nand U11622 (N_11622,N_10282,N_10169);
or U11623 (N_11623,N_9092,N_9000);
xor U11624 (N_11624,N_9388,N_9129);
and U11625 (N_11625,N_10461,N_9415);
xnor U11626 (N_11626,N_9088,N_9688);
or U11627 (N_11627,N_10167,N_9809);
and U11628 (N_11628,N_10367,N_9603);
or U11629 (N_11629,N_9567,N_9719);
nand U11630 (N_11630,N_9604,N_10077);
or U11631 (N_11631,N_9874,N_9116);
or U11632 (N_11632,N_9540,N_9752);
and U11633 (N_11633,N_9252,N_9554);
nand U11634 (N_11634,N_9837,N_9479);
or U11635 (N_11635,N_9963,N_10004);
or U11636 (N_11636,N_9549,N_10066);
xor U11637 (N_11637,N_9284,N_9477);
xnor U11638 (N_11638,N_9006,N_9648);
xnor U11639 (N_11639,N_9426,N_10498);
nor U11640 (N_11640,N_9107,N_9353);
nor U11641 (N_11641,N_9330,N_9701);
nor U11642 (N_11642,N_9351,N_9468);
nor U11643 (N_11643,N_9494,N_9658);
xor U11644 (N_11644,N_9072,N_10182);
and U11645 (N_11645,N_9577,N_9797);
xnor U11646 (N_11646,N_9932,N_10156);
and U11647 (N_11647,N_9522,N_10006);
nor U11648 (N_11648,N_10422,N_9995);
and U11649 (N_11649,N_9561,N_9032);
or U11650 (N_11650,N_9243,N_9154);
nor U11651 (N_11651,N_9357,N_9156);
or U11652 (N_11652,N_9369,N_9132);
nand U11653 (N_11653,N_9599,N_10352);
nand U11654 (N_11654,N_9403,N_10140);
nor U11655 (N_11655,N_9481,N_10193);
and U11656 (N_11656,N_9196,N_9353);
nor U11657 (N_11657,N_9381,N_9827);
nor U11658 (N_11658,N_9370,N_10105);
nor U11659 (N_11659,N_9567,N_9725);
nor U11660 (N_11660,N_9084,N_9648);
and U11661 (N_11661,N_10028,N_9493);
nor U11662 (N_11662,N_9249,N_9923);
nor U11663 (N_11663,N_10213,N_9714);
nand U11664 (N_11664,N_10400,N_9236);
nor U11665 (N_11665,N_9127,N_9433);
and U11666 (N_11666,N_9647,N_10359);
and U11667 (N_11667,N_9109,N_9919);
or U11668 (N_11668,N_10465,N_9770);
nor U11669 (N_11669,N_10436,N_10434);
and U11670 (N_11670,N_10161,N_9047);
nor U11671 (N_11671,N_9541,N_10435);
or U11672 (N_11672,N_9411,N_9731);
and U11673 (N_11673,N_9985,N_9427);
xor U11674 (N_11674,N_9120,N_9475);
and U11675 (N_11675,N_10161,N_10044);
or U11676 (N_11676,N_9961,N_9295);
nand U11677 (N_11677,N_10464,N_9032);
or U11678 (N_11678,N_9846,N_9905);
and U11679 (N_11679,N_9714,N_10394);
or U11680 (N_11680,N_10068,N_9267);
nor U11681 (N_11681,N_10212,N_9664);
nand U11682 (N_11682,N_9645,N_9827);
or U11683 (N_11683,N_10304,N_9976);
nor U11684 (N_11684,N_10393,N_10116);
or U11685 (N_11685,N_10473,N_9625);
xnor U11686 (N_11686,N_9966,N_9692);
and U11687 (N_11687,N_10179,N_9813);
and U11688 (N_11688,N_9583,N_9982);
and U11689 (N_11689,N_10425,N_9168);
nor U11690 (N_11690,N_9536,N_10254);
nand U11691 (N_11691,N_10278,N_9182);
or U11692 (N_11692,N_9817,N_9504);
nand U11693 (N_11693,N_9880,N_9890);
or U11694 (N_11694,N_9078,N_9214);
or U11695 (N_11695,N_9886,N_9052);
and U11696 (N_11696,N_10011,N_9314);
xnor U11697 (N_11697,N_10015,N_10240);
and U11698 (N_11698,N_9109,N_9480);
nor U11699 (N_11699,N_9214,N_9693);
or U11700 (N_11700,N_9309,N_10490);
or U11701 (N_11701,N_10101,N_9725);
or U11702 (N_11702,N_10297,N_10427);
nand U11703 (N_11703,N_9927,N_10412);
nand U11704 (N_11704,N_9417,N_9259);
xor U11705 (N_11705,N_9816,N_10451);
and U11706 (N_11706,N_9219,N_9284);
and U11707 (N_11707,N_10024,N_10169);
or U11708 (N_11708,N_9034,N_9806);
or U11709 (N_11709,N_9779,N_10401);
or U11710 (N_11710,N_9663,N_9407);
xnor U11711 (N_11711,N_10130,N_9835);
nand U11712 (N_11712,N_9510,N_10196);
or U11713 (N_11713,N_9331,N_10262);
or U11714 (N_11714,N_9208,N_9399);
nor U11715 (N_11715,N_9553,N_9719);
and U11716 (N_11716,N_10253,N_10248);
nand U11717 (N_11717,N_9533,N_9813);
nor U11718 (N_11718,N_10460,N_10105);
and U11719 (N_11719,N_9065,N_9956);
or U11720 (N_11720,N_10163,N_10337);
nor U11721 (N_11721,N_10117,N_10227);
or U11722 (N_11722,N_9374,N_9390);
xor U11723 (N_11723,N_10297,N_9175);
nor U11724 (N_11724,N_10406,N_10068);
xor U11725 (N_11725,N_9337,N_10413);
xnor U11726 (N_11726,N_10230,N_10243);
or U11727 (N_11727,N_9977,N_10440);
nor U11728 (N_11728,N_9795,N_9353);
or U11729 (N_11729,N_9299,N_9547);
and U11730 (N_11730,N_9723,N_10147);
xor U11731 (N_11731,N_9930,N_9963);
and U11732 (N_11732,N_10091,N_9293);
nor U11733 (N_11733,N_10010,N_9355);
or U11734 (N_11734,N_9485,N_9047);
nor U11735 (N_11735,N_10026,N_9002);
or U11736 (N_11736,N_9233,N_9900);
nand U11737 (N_11737,N_10245,N_9675);
nor U11738 (N_11738,N_9956,N_9200);
and U11739 (N_11739,N_9945,N_9210);
or U11740 (N_11740,N_9006,N_10491);
nand U11741 (N_11741,N_9018,N_9023);
nand U11742 (N_11742,N_10424,N_10061);
nand U11743 (N_11743,N_9917,N_9528);
nand U11744 (N_11744,N_9797,N_9007);
xor U11745 (N_11745,N_9518,N_9660);
or U11746 (N_11746,N_10322,N_9864);
or U11747 (N_11747,N_9707,N_9570);
or U11748 (N_11748,N_10058,N_9042);
or U11749 (N_11749,N_9961,N_9478);
xnor U11750 (N_11750,N_10254,N_9378);
nand U11751 (N_11751,N_9703,N_9233);
nor U11752 (N_11752,N_10202,N_9909);
nand U11753 (N_11753,N_9963,N_9387);
and U11754 (N_11754,N_9780,N_10049);
xor U11755 (N_11755,N_10246,N_10472);
nor U11756 (N_11756,N_10058,N_9386);
nor U11757 (N_11757,N_9889,N_10110);
and U11758 (N_11758,N_10454,N_10226);
nor U11759 (N_11759,N_10149,N_9355);
xnor U11760 (N_11760,N_10071,N_9474);
nor U11761 (N_11761,N_10443,N_9055);
nor U11762 (N_11762,N_10144,N_9621);
or U11763 (N_11763,N_9053,N_9315);
and U11764 (N_11764,N_9062,N_9464);
nor U11765 (N_11765,N_9617,N_9027);
nor U11766 (N_11766,N_9952,N_9063);
nor U11767 (N_11767,N_10452,N_9791);
or U11768 (N_11768,N_9026,N_9074);
nor U11769 (N_11769,N_9552,N_10498);
or U11770 (N_11770,N_9282,N_9540);
nor U11771 (N_11771,N_9406,N_9853);
nand U11772 (N_11772,N_9910,N_9074);
and U11773 (N_11773,N_9038,N_9321);
nand U11774 (N_11774,N_9094,N_10328);
nand U11775 (N_11775,N_9586,N_9403);
nor U11776 (N_11776,N_9293,N_10463);
nand U11777 (N_11777,N_9661,N_10214);
and U11778 (N_11778,N_10106,N_9265);
nand U11779 (N_11779,N_10148,N_10130);
or U11780 (N_11780,N_9443,N_9585);
nand U11781 (N_11781,N_9958,N_10098);
nor U11782 (N_11782,N_9797,N_10301);
nor U11783 (N_11783,N_10276,N_10323);
nor U11784 (N_11784,N_9182,N_10177);
nor U11785 (N_11785,N_9062,N_10219);
nand U11786 (N_11786,N_10296,N_9619);
or U11787 (N_11787,N_10366,N_9478);
nor U11788 (N_11788,N_10295,N_9101);
nor U11789 (N_11789,N_9647,N_10440);
nand U11790 (N_11790,N_10406,N_9583);
xnor U11791 (N_11791,N_10156,N_9739);
xor U11792 (N_11792,N_10482,N_10344);
nor U11793 (N_11793,N_9043,N_9399);
and U11794 (N_11794,N_9884,N_9841);
nor U11795 (N_11795,N_9118,N_10252);
and U11796 (N_11796,N_9287,N_10391);
and U11797 (N_11797,N_9855,N_9297);
or U11798 (N_11798,N_10364,N_10396);
or U11799 (N_11799,N_9117,N_9599);
nor U11800 (N_11800,N_9788,N_10086);
nand U11801 (N_11801,N_10304,N_9906);
nand U11802 (N_11802,N_9314,N_9323);
nor U11803 (N_11803,N_9053,N_9535);
and U11804 (N_11804,N_9925,N_9694);
and U11805 (N_11805,N_9432,N_9771);
and U11806 (N_11806,N_10497,N_9222);
or U11807 (N_11807,N_9154,N_9645);
and U11808 (N_11808,N_9099,N_10080);
or U11809 (N_11809,N_9021,N_9872);
nand U11810 (N_11810,N_9818,N_9346);
nand U11811 (N_11811,N_9160,N_9720);
nor U11812 (N_11812,N_10419,N_9771);
nor U11813 (N_11813,N_9535,N_9054);
and U11814 (N_11814,N_9801,N_10320);
and U11815 (N_11815,N_10063,N_10100);
and U11816 (N_11816,N_9132,N_10063);
nor U11817 (N_11817,N_9019,N_9000);
or U11818 (N_11818,N_10022,N_10138);
or U11819 (N_11819,N_10074,N_9281);
and U11820 (N_11820,N_9699,N_9196);
or U11821 (N_11821,N_10211,N_9162);
nand U11822 (N_11822,N_10169,N_9579);
nand U11823 (N_11823,N_9184,N_9054);
nor U11824 (N_11824,N_9912,N_9453);
xnor U11825 (N_11825,N_9093,N_9078);
nand U11826 (N_11826,N_9770,N_9535);
or U11827 (N_11827,N_9464,N_9479);
xor U11828 (N_11828,N_9721,N_9988);
nor U11829 (N_11829,N_10019,N_9678);
and U11830 (N_11830,N_10456,N_10446);
or U11831 (N_11831,N_9166,N_9839);
nor U11832 (N_11832,N_9582,N_10213);
or U11833 (N_11833,N_9915,N_9326);
nor U11834 (N_11834,N_9049,N_10245);
nand U11835 (N_11835,N_9124,N_10239);
and U11836 (N_11836,N_10254,N_9784);
and U11837 (N_11837,N_10152,N_9869);
and U11838 (N_11838,N_9467,N_9733);
nand U11839 (N_11839,N_9582,N_10022);
or U11840 (N_11840,N_9705,N_9909);
or U11841 (N_11841,N_10150,N_9315);
or U11842 (N_11842,N_9695,N_9259);
and U11843 (N_11843,N_9016,N_9508);
nor U11844 (N_11844,N_9518,N_9617);
and U11845 (N_11845,N_9430,N_9453);
nor U11846 (N_11846,N_10284,N_9414);
nand U11847 (N_11847,N_9572,N_9675);
and U11848 (N_11848,N_10341,N_10210);
nand U11849 (N_11849,N_9894,N_9663);
and U11850 (N_11850,N_10022,N_10282);
xor U11851 (N_11851,N_9788,N_10039);
nand U11852 (N_11852,N_9871,N_9044);
and U11853 (N_11853,N_9002,N_9420);
nand U11854 (N_11854,N_10023,N_10442);
or U11855 (N_11855,N_10404,N_9220);
nor U11856 (N_11856,N_9918,N_10476);
nor U11857 (N_11857,N_10114,N_10207);
nand U11858 (N_11858,N_9237,N_9016);
or U11859 (N_11859,N_9998,N_10244);
nand U11860 (N_11860,N_10280,N_9363);
nand U11861 (N_11861,N_9998,N_9835);
and U11862 (N_11862,N_10294,N_9336);
and U11863 (N_11863,N_9661,N_9367);
or U11864 (N_11864,N_9432,N_10173);
nand U11865 (N_11865,N_9110,N_9914);
or U11866 (N_11866,N_10394,N_10322);
and U11867 (N_11867,N_10075,N_9093);
and U11868 (N_11868,N_9454,N_10394);
nand U11869 (N_11869,N_9698,N_9255);
nand U11870 (N_11870,N_9752,N_9428);
nor U11871 (N_11871,N_9082,N_10124);
nand U11872 (N_11872,N_10260,N_9177);
and U11873 (N_11873,N_9826,N_9459);
and U11874 (N_11874,N_9002,N_9293);
and U11875 (N_11875,N_9029,N_10466);
nand U11876 (N_11876,N_10197,N_9596);
nand U11877 (N_11877,N_9275,N_9663);
nand U11878 (N_11878,N_10072,N_9430);
xnor U11879 (N_11879,N_10230,N_9644);
nand U11880 (N_11880,N_9328,N_10364);
or U11881 (N_11881,N_9449,N_9733);
or U11882 (N_11882,N_9751,N_9022);
and U11883 (N_11883,N_9766,N_10450);
nand U11884 (N_11884,N_9648,N_9775);
xor U11885 (N_11885,N_10068,N_10060);
xor U11886 (N_11886,N_10036,N_9059);
nor U11887 (N_11887,N_10474,N_9536);
nor U11888 (N_11888,N_9430,N_10297);
xnor U11889 (N_11889,N_10120,N_9256);
and U11890 (N_11890,N_10421,N_9926);
nor U11891 (N_11891,N_9641,N_9993);
and U11892 (N_11892,N_9091,N_9973);
nor U11893 (N_11893,N_10186,N_9228);
or U11894 (N_11894,N_9755,N_9441);
nand U11895 (N_11895,N_9342,N_10311);
xor U11896 (N_11896,N_9290,N_10498);
nor U11897 (N_11897,N_9032,N_9847);
and U11898 (N_11898,N_10400,N_10470);
nor U11899 (N_11899,N_9717,N_9710);
or U11900 (N_11900,N_9376,N_9142);
or U11901 (N_11901,N_9560,N_10157);
nand U11902 (N_11902,N_9842,N_10235);
nor U11903 (N_11903,N_9701,N_9302);
nand U11904 (N_11904,N_9464,N_10131);
nor U11905 (N_11905,N_10179,N_10474);
and U11906 (N_11906,N_9061,N_10057);
nor U11907 (N_11907,N_9843,N_9091);
and U11908 (N_11908,N_9033,N_9741);
or U11909 (N_11909,N_9751,N_10430);
or U11910 (N_11910,N_9787,N_10323);
and U11911 (N_11911,N_9421,N_9244);
xor U11912 (N_11912,N_9484,N_9444);
nand U11913 (N_11913,N_10484,N_9952);
xnor U11914 (N_11914,N_9311,N_9619);
nor U11915 (N_11915,N_9251,N_9214);
nor U11916 (N_11916,N_9723,N_10287);
xnor U11917 (N_11917,N_9393,N_10488);
nand U11918 (N_11918,N_9999,N_9040);
and U11919 (N_11919,N_9876,N_10126);
nor U11920 (N_11920,N_10112,N_10363);
nor U11921 (N_11921,N_10240,N_9607);
and U11922 (N_11922,N_10478,N_9023);
nand U11923 (N_11923,N_9150,N_9491);
xor U11924 (N_11924,N_10266,N_9187);
or U11925 (N_11925,N_9662,N_10429);
or U11926 (N_11926,N_10368,N_10430);
nand U11927 (N_11927,N_10362,N_10428);
or U11928 (N_11928,N_9096,N_10358);
and U11929 (N_11929,N_10276,N_10166);
or U11930 (N_11930,N_9905,N_9104);
nor U11931 (N_11931,N_9886,N_10068);
and U11932 (N_11932,N_9724,N_10271);
nand U11933 (N_11933,N_9392,N_9763);
nor U11934 (N_11934,N_9095,N_9346);
or U11935 (N_11935,N_9721,N_9314);
and U11936 (N_11936,N_10314,N_9293);
and U11937 (N_11937,N_9733,N_9070);
nor U11938 (N_11938,N_10326,N_9987);
and U11939 (N_11939,N_10399,N_10408);
and U11940 (N_11940,N_9880,N_9198);
nor U11941 (N_11941,N_10103,N_9428);
or U11942 (N_11942,N_10131,N_9121);
or U11943 (N_11943,N_10116,N_9409);
and U11944 (N_11944,N_10317,N_9206);
or U11945 (N_11945,N_10489,N_10451);
and U11946 (N_11946,N_9227,N_10437);
nand U11947 (N_11947,N_10125,N_9844);
and U11948 (N_11948,N_10102,N_10171);
nor U11949 (N_11949,N_10412,N_10463);
or U11950 (N_11950,N_9750,N_9712);
xor U11951 (N_11951,N_9883,N_10190);
or U11952 (N_11952,N_9969,N_10484);
nor U11953 (N_11953,N_9431,N_10094);
and U11954 (N_11954,N_9832,N_9649);
xnor U11955 (N_11955,N_9167,N_10054);
and U11956 (N_11956,N_10243,N_10308);
and U11957 (N_11957,N_9436,N_9787);
and U11958 (N_11958,N_10311,N_9753);
and U11959 (N_11959,N_10112,N_9486);
nor U11960 (N_11960,N_9735,N_9764);
nor U11961 (N_11961,N_10283,N_9147);
or U11962 (N_11962,N_9195,N_9789);
nor U11963 (N_11963,N_10261,N_9567);
and U11964 (N_11964,N_10061,N_9014);
and U11965 (N_11965,N_9257,N_9486);
nand U11966 (N_11966,N_9786,N_9102);
nor U11967 (N_11967,N_9649,N_9416);
nand U11968 (N_11968,N_10324,N_9623);
nand U11969 (N_11969,N_9461,N_10483);
or U11970 (N_11970,N_9355,N_10143);
nand U11971 (N_11971,N_9208,N_9176);
nand U11972 (N_11972,N_9237,N_10227);
nand U11973 (N_11973,N_9049,N_9209);
nand U11974 (N_11974,N_9610,N_10294);
and U11975 (N_11975,N_9721,N_10378);
or U11976 (N_11976,N_9102,N_10122);
nand U11977 (N_11977,N_9242,N_9262);
xor U11978 (N_11978,N_9710,N_9075);
nand U11979 (N_11979,N_10075,N_10210);
or U11980 (N_11980,N_9214,N_9711);
nor U11981 (N_11981,N_9006,N_9798);
nand U11982 (N_11982,N_9053,N_9294);
nand U11983 (N_11983,N_10387,N_10021);
nand U11984 (N_11984,N_9595,N_9089);
and U11985 (N_11985,N_9709,N_9007);
or U11986 (N_11986,N_9827,N_9744);
or U11987 (N_11987,N_9156,N_9188);
or U11988 (N_11988,N_10088,N_10272);
and U11989 (N_11989,N_10385,N_9126);
or U11990 (N_11990,N_9929,N_9090);
xnor U11991 (N_11991,N_9192,N_9275);
or U11992 (N_11992,N_10271,N_9169);
nand U11993 (N_11993,N_9692,N_9956);
nand U11994 (N_11994,N_10178,N_9029);
or U11995 (N_11995,N_10114,N_9313);
xnor U11996 (N_11996,N_9660,N_9963);
or U11997 (N_11997,N_9469,N_10184);
and U11998 (N_11998,N_9210,N_10236);
xor U11999 (N_11999,N_9467,N_9162);
or U12000 (N_12000,N_11239,N_10823);
or U12001 (N_12001,N_10903,N_10831);
nand U12002 (N_12002,N_10885,N_11820);
or U12003 (N_12003,N_11135,N_10884);
nor U12004 (N_12004,N_11380,N_11600);
xor U12005 (N_12005,N_11522,N_11274);
nand U12006 (N_12006,N_10891,N_11310);
and U12007 (N_12007,N_11771,N_10519);
nand U12008 (N_12008,N_11871,N_10778);
xnor U12009 (N_12009,N_10857,N_10717);
nor U12010 (N_12010,N_10787,N_11457);
nand U12011 (N_12011,N_11726,N_11701);
nor U12012 (N_12012,N_11219,N_10541);
and U12013 (N_12013,N_11212,N_11353);
xor U12014 (N_12014,N_11719,N_10575);
and U12015 (N_12015,N_11238,N_11141);
nor U12016 (N_12016,N_11610,N_11288);
or U12017 (N_12017,N_11371,N_11127);
and U12018 (N_12018,N_11104,N_11231);
and U12019 (N_12019,N_11328,N_10629);
nor U12020 (N_12020,N_11080,N_10759);
nor U12021 (N_12021,N_10913,N_11117);
nor U12022 (N_12022,N_11638,N_11533);
nor U12023 (N_12023,N_10525,N_11799);
and U12024 (N_12024,N_10739,N_11076);
nor U12025 (N_12025,N_10639,N_11768);
xor U12026 (N_12026,N_11861,N_11131);
nor U12027 (N_12027,N_11082,N_10950);
nand U12028 (N_12028,N_10731,N_11002);
and U12029 (N_12029,N_11634,N_10988);
and U12030 (N_12030,N_11263,N_10930);
nor U12031 (N_12031,N_11366,N_11460);
nor U12032 (N_12032,N_11195,N_10723);
xor U12033 (N_12033,N_10843,N_10758);
or U12034 (N_12034,N_11254,N_11473);
and U12035 (N_12035,N_10924,N_10509);
or U12036 (N_12036,N_11982,N_10667);
or U12037 (N_12037,N_10669,N_11912);
or U12038 (N_12038,N_11001,N_11168);
nand U12039 (N_12039,N_11869,N_11216);
and U12040 (N_12040,N_11904,N_10646);
or U12041 (N_12041,N_11493,N_11971);
or U12042 (N_12042,N_11287,N_11100);
or U12043 (N_12043,N_10626,N_11857);
or U12044 (N_12044,N_11650,N_10755);
or U12045 (N_12045,N_11077,N_11387);
nand U12046 (N_12046,N_10919,N_11268);
xnor U12047 (N_12047,N_10662,N_10527);
or U12048 (N_12048,N_11188,N_11773);
nor U12049 (N_12049,N_10599,N_10564);
nand U12050 (N_12050,N_11764,N_11792);
or U12051 (N_12051,N_11065,N_11569);
or U12052 (N_12052,N_11936,N_10594);
nor U12053 (N_12053,N_10945,N_11040);
and U12054 (N_12054,N_10867,N_11319);
nor U12055 (N_12055,N_11044,N_10542);
or U12056 (N_12056,N_11558,N_11518);
nor U12057 (N_12057,N_11469,N_10786);
or U12058 (N_12058,N_11616,N_11752);
nand U12059 (N_12059,N_10651,N_10526);
and U12060 (N_12060,N_11261,N_10830);
nor U12061 (N_12061,N_11934,N_11215);
or U12062 (N_12062,N_11047,N_11363);
and U12063 (N_12063,N_11631,N_10794);
xnor U12064 (N_12064,N_10576,N_11580);
nor U12065 (N_12065,N_11759,N_10934);
nor U12066 (N_12066,N_11521,N_11588);
nor U12067 (N_12067,N_10508,N_11273);
nand U12068 (N_12068,N_11136,N_11063);
nand U12069 (N_12069,N_10746,N_11345);
nor U12070 (N_12070,N_11809,N_10502);
nand U12071 (N_12071,N_11028,N_10590);
nand U12072 (N_12072,N_11962,N_11464);
nand U12073 (N_12073,N_11560,N_11480);
and U12074 (N_12074,N_11710,N_10677);
and U12075 (N_12075,N_11488,N_10876);
or U12076 (N_12076,N_11780,N_10954);
xnor U12077 (N_12077,N_11022,N_10998);
and U12078 (N_12078,N_11813,N_11408);
and U12079 (N_12079,N_11005,N_11414);
nand U12080 (N_12080,N_11901,N_10939);
or U12081 (N_12081,N_11333,N_10844);
nand U12082 (N_12082,N_11253,N_11180);
nand U12083 (N_12083,N_11132,N_10745);
nand U12084 (N_12084,N_10562,N_11889);
and U12085 (N_12085,N_11327,N_11921);
nand U12086 (N_12086,N_11171,N_11092);
nor U12087 (N_12087,N_10559,N_11476);
xnor U12088 (N_12088,N_11787,N_11283);
nand U12089 (N_12089,N_11781,N_11386);
or U12090 (N_12090,N_10846,N_10949);
and U12091 (N_12091,N_11743,N_11107);
xnor U12092 (N_12092,N_11264,N_11138);
or U12093 (N_12093,N_11659,N_11983);
nor U12094 (N_12094,N_11206,N_10929);
nor U12095 (N_12095,N_10571,N_10563);
or U12096 (N_12096,N_10583,N_11639);
nand U12097 (N_12097,N_11658,N_11038);
nand U12098 (N_12098,N_11395,N_11917);
or U12099 (N_12099,N_11584,N_10663);
and U12100 (N_12100,N_11008,N_11556);
or U12101 (N_12101,N_11826,N_11794);
and U12102 (N_12102,N_11730,N_11644);
nand U12103 (N_12103,N_10781,N_10753);
or U12104 (N_12104,N_11204,N_10738);
nand U12105 (N_12105,N_11089,N_10771);
nor U12106 (N_12106,N_11401,N_11947);
nand U12107 (N_12107,N_10767,N_10656);
and U12108 (N_12108,N_11672,N_10647);
nand U12109 (N_12109,N_11858,N_11924);
xor U12110 (N_12110,N_11843,N_10572);
or U12111 (N_12111,N_11466,N_10500);
or U12112 (N_12112,N_10806,N_11055);
xnor U12113 (N_12113,N_10592,N_11839);
or U12114 (N_12114,N_10616,N_10588);
nand U12115 (N_12115,N_11611,N_11073);
and U12116 (N_12116,N_11126,N_10896);
nand U12117 (N_12117,N_10586,N_10904);
and U12118 (N_12118,N_11406,N_11834);
nand U12119 (N_12119,N_10504,N_11840);
nand U12120 (N_12120,N_11234,N_11191);
xor U12121 (N_12121,N_11756,N_11472);
nand U12122 (N_12122,N_11045,N_10804);
and U12123 (N_12123,N_10879,N_10899);
nand U12124 (N_12124,N_11693,N_11489);
and U12125 (N_12125,N_10643,N_10754);
nor U12126 (N_12126,N_10932,N_11143);
or U12127 (N_12127,N_11242,N_11437);
and U12128 (N_12128,N_11289,N_10687);
or U12129 (N_12129,N_11657,N_10824);
or U12130 (N_12130,N_10873,N_11897);
nor U12131 (N_12131,N_11281,N_10832);
xor U12132 (N_12132,N_11785,N_11915);
nor U12133 (N_12133,N_11448,N_11715);
xnor U12134 (N_12134,N_11147,N_11999);
and U12135 (N_12135,N_11483,N_11790);
or U12136 (N_12136,N_10727,N_10701);
nor U12137 (N_12137,N_11456,N_11892);
and U12138 (N_12138,N_11425,N_10579);
or U12139 (N_12139,N_11302,N_11583);
and U12140 (N_12140,N_10880,N_11398);
nor U12141 (N_12141,N_10619,N_11882);
nor U12142 (N_12142,N_11895,N_11789);
nor U12143 (N_12143,N_11949,N_11221);
or U12144 (N_12144,N_11338,N_11872);
and U12145 (N_12145,N_11262,N_11649);
and U12146 (N_12146,N_11832,N_11714);
or U12147 (N_12147,N_11067,N_10819);
nor U12148 (N_12148,N_10574,N_11155);
nand U12149 (N_12149,N_11314,N_10697);
nor U12150 (N_12150,N_10972,N_10603);
xnor U12151 (N_12151,N_11898,N_11595);
nor U12152 (N_12152,N_11060,N_11686);
xor U12153 (N_12153,N_10636,N_11545);
nor U12154 (N_12154,N_11462,N_10732);
nand U12155 (N_12155,N_11032,N_11511);
nand U12156 (N_12156,N_11750,N_11244);
or U12157 (N_12157,N_10625,N_11276);
and U12158 (N_12158,N_10751,N_10851);
xor U12159 (N_12159,N_11808,N_11899);
nor U12160 (N_12160,N_10997,N_11442);
and U12161 (N_12161,N_10910,N_10882);
xnor U12162 (N_12162,N_11939,N_10784);
and U12163 (N_12163,N_11849,N_11455);
and U12164 (N_12164,N_11246,N_10868);
or U12165 (N_12165,N_11389,N_10573);
xnor U12166 (N_12166,N_11308,N_11122);
or U12167 (N_12167,N_11252,N_11612);
or U12168 (N_12168,N_10796,N_11515);
and U12169 (N_12169,N_11227,N_10838);
or U12170 (N_12170,N_10975,N_11179);
nor U12171 (N_12171,N_10587,N_10505);
nand U12172 (N_12172,N_10822,N_11670);
and U12173 (N_12173,N_11189,N_10980);
and U12174 (N_12174,N_11602,N_11452);
or U12175 (N_12175,N_10772,N_11029);
nor U12176 (N_12176,N_11667,N_11745);
nand U12177 (N_12177,N_10623,N_11304);
or U12178 (N_12178,N_10691,N_10987);
and U12179 (N_12179,N_10637,N_11011);
nand U12180 (N_12180,N_10769,N_11149);
nor U12181 (N_12181,N_10514,N_11039);
nor U12182 (N_12182,N_10999,N_10718);
xor U12183 (N_12183,N_11876,N_10992);
or U12184 (N_12184,N_11959,N_10604);
xor U12185 (N_12185,N_10577,N_11525);
or U12186 (N_12186,N_10807,N_11512);
nor U12187 (N_12187,N_10631,N_11443);
and U12188 (N_12188,N_11056,N_11669);
nand U12189 (N_12189,N_11050,N_10989);
or U12190 (N_12190,N_11075,N_10561);
and U12191 (N_12191,N_11579,N_10704);
xnor U12192 (N_12192,N_11978,N_11633);
or U12193 (N_12193,N_11110,N_10907);
xnor U12194 (N_12194,N_11852,N_11203);
nor U12195 (N_12195,N_11767,N_11546);
or U12196 (N_12196,N_11628,N_11016);
nand U12197 (N_12197,N_10531,N_10538);
or U12198 (N_12198,N_10721,N_10979);
and U12199 (N_12199,N_10971,N_10560);
nor U12200 (N_12200,N_11927,N_11119);
nand U12201 (N_12201,N_11953,N_11224);
xor U12202 (N_12202,N_11913,N_11435);
nor U12203 (N_12203,N_10863,N_10779);
xnor U12204 (N_12204,N_11361,N_11940);
or U12205 (N_12205,N_11997,N_11996);
nand U12206 (N_12206,N_10618,N_11397);
and U12207 (N_12207,N_11747,N_10711);
and U12208 (N_12208,N_10558,N_11793);
nor U12209 (N_12209,N_11164,N_11950);
and U12210 (N_12210,N_11641,N_11381);
nand U12211 (N_12211,N_11024,N_11175);
nand U12212 (N_12212,N_11585,N_11285);
xor U12213 (N_12213,N_11534,N_11542);
or U12214 (N_12214,N_11705,N_10921);
and U12215 (N_12215,N_11286,N_11935);
xnor U12216 (N_12216,N_11378,N_11417);
nand U12217 (N_12217,N_11259,N_11842);
or U12218 (N_12218,N_11559,N_10617);
nand U12219 (N_12219,N_11689,N_10915);
nor U12220 (N_12220,N_10640,N_10871);
or U12221 (N_12221,N_10817,N_11210);
or U12222 (N_12222,N_10776,N_11294);
nor U12223 (N_12223,N_11961,N_10749);
nor U12224 (N_12224,N_11128,N_10931);
xnor U12225 (N_12225,N_11535,N_11643);
nand U12226 (N_12226,N_11879,N_11567);
or U12227 (N_12227,N_10734,N_11890);
and U12228 (N_12228,N_11405,N_10528);
nor U12229 (N_12229,N_11292,N_11791);
and U12230 (N_12230,N_11860,N_11208);
nor U12231 (N_12231,N_11520,N_10803);
nor U12232 (N_12232,N_11727,N_11181);
nand U12233 (N_12233,N_11150,N_10735);
nor U12234 (N_12234,N_10518,N_11492);
or U12235 (N_12235,N_11440,N_11250);
nor U12236 (N_12236,N_10792,N_11097);
nor U12237 (N_12237,N_10695,N_11249);
nand U12238 (N_12238,N_11571,N_11153);
or U12239 (N_12239,N_10578,N_11035);
nand U12240 (N_12240,N_11906,N_10935);
and U12241 (N_12241,N_11875,N_11527);
or U12242 (N_12242,N_11561,N_11017);
and U12243 (N_12243,N_11444,N_11152);
nor U12244 (N_12244,N_11748,N_11335);
nor U12245 (N_12245,N_11724,N_11903);
xnor U12246 (N_12246,N_11058,N_10596);
nand U12247 (N_12247,N_10535,N_11803);
or U12248 (N_12248,N_11223,N_11332);
xnor U12249 (N_12249,N_10875,N_11736);
nand U12250 (N_12250,N_11679,N_11481);
and U12251 (N_12251,N_10908,N_11360);
or U12252 (N_12252,N_10624,N_11981);
and U12253 (N_12253,N_11270,N_10614);
nand U12254 (N_12254,N_10606,N_11859);
or U12255 (N_12255,N_11680,N_10984);
nor U12256 (N_12256,N_10620,N_10981);
nor U12257 (N_12257,N_10977,N_11108);
nand U12258 (N_12258,N_11233,N_10705);
nand U12259 (N_12259,N_11267,N_11272);
and U12260 (N_12260,N_11735,N_11866);
nand U12261 (N_12261,N_10985,N_11572);
or U12262 (N_12262,N_10568,N_10671);
xnor U12263 (N_12263,N_11677,N_11301);
and U12264 (N_12264,N_10925,N_10696);
and U12265 (N_12265,N_10709,N_10835);
and U12266 (N_12266,N_11887,N_11399);
nor U12267 (N_12267,N_10976,N_10955);
or U12268 (N_12268,N_10549,N_11676);
and U12269 (N_12269,N_10865,N_11433);
nand U12270 (N_12270,N_10657,N_11847);
or U12271 (N_12271,N_11364,N_10893);
or U12272 (N_12272,N_11955,N_10920);
nor U12273 (N_12273,N_11980,N_11691);
nor U12274 (N_12274,N_11937,N_10902);
and U12275 (N_12275,N_11337,N_10861);
nor U12276 (N_12276,N_10548,N_10836);
and U12277 (N_12277,N_11798,N_11954);
or U12278 (N_12278,N_10881,N_10869);
and U12279 (N_12279,N_11322,N_11427);
nand U12280 (N_12280,N_10829,N_11192);
xnor U12281 (N_12281,N_11323,N_10533);
or U12282 (N_12282,N_11966,N_10556);
and U12283 (N_12283,N_11368,N_11574);
or U12284 (N_12284,N_11091,N_11036);
and U12285 (N_12285,N_11685,N_11751);
or U12286 (N_12286,N_11712,N_11217);
nor U12287 (N_12287,N_11963,N_10540);
and U12288 (N_12288,N_11597,N_10911);
nor U12289 (N_12289,N_11877,N_10744);
nand U12290 (N_12290,N_11315,N_11528);
or U12291 (N_12291,N_10760,N_11683);
nor U12292 (N_12292,N_11801,N_11176);
nand U12293 (N_12293,N_10933,N_11404);
and U12294 (N_12294,N_11922,N_10642);
nor U12295 (N_12295,N_11509,N_10849);
nor U12296 (N_12296,N_11213,N_10569);
and U12297 (N_12297,N_10813,N_10591);
nor U12298 (N_12298,N_11833,N_11998);
xor U12299 (N_12299,N_11888,N_10940);
or U12300 (N_12300,N_10644,N_11495);
nand U12301 (N_12301,N_10700,N_11409);
and U12302 (N_12302,N_11721,N_11295);
nor U12303 (N_12303,N_11990,N_10553);
nand U12304 (N_12304,N_11392,N_10510);
and U12305 (N_12305,N_10589,N_10664);
nor U12306 (N_12306,N_11766,N_11451);
nand U12307 (N_12307,N_11873,N_11548);
or U12308 (N_12308,N_11587,N_10650);
nand U12309 (N_12309,N_11737,N_11436);
nand U12310 (N_12310,N_11948,N_11694);
and U12311 (N_12311,N_11486,N_11688);
xor U12312 (N_12312,N_11069,N_10543);
xor U12313 (N_12313,N_10668,N_11053);
nor U12314 (N_12314,N_11566,N_11403);
nor U12315 (N_12315,N_11081,N_11064);
or U12316 (N_12316,N_10546,N_10959);
nor U12317 (N_12317,N_11564,N_11207);
or U12318 (N_12318,N_11358,N_10809);
and U12319 (N_12319,N_10648,N_11115);
or U12320 (N_12320,N_10918,N_11183);
nand U12321 (N_12321,N_11049,N_11532);
and U12322 (N_12322,N_11968,N_11986);
and U12323 (N_12323,N_10886,N_11431);
nand U12324 (N_12324,N_10678,N_11275);
nand U12325 (N_12325,N_11365,N_11151);
nor U12326 (N_12326,N_11988,N_11072);
and U12327 (N_12327,N_11474,N_10748);
nor U12328 (N_12328,N_11084,N_11394);
nand U12329 (N_12329,N_10593,N_11342);
xnor U12330 (N_12330,N_11265,N_10565);
or U12331 (N_12331,N_10845,N_11992);
nand U12332 (N_12332,N_10900,N_11987);
or U12333 (N_12333,N_11426,N_11874);
and U12334 (N_12334,N_11539,N_11795);
xnor U12335 (N_12335,N_11218,N_11868);
nor U12336 (N_12336,N_11823,N_10686);
or U12337 (N_12337,N_10888,N_10737);
or U12338 (N_12338,N_11805,N_11194);
and U12339 (N_12339,N_11979,N_11530);
xor U12340 (N_12340,N_11905,N_10958);
or U12341 (N_12341,N_11505,N_11880);
and U12342 (N_12342,N_11382,N_11837);
and U12343 (N_12343,N_11973,N_10842);
or U12344 (N_12344,N_11484,N_11173);
xnor U12345 (N_12345,N_11157,N_11297);
or U12346 (N_12346,N_10928,N_11606);
nand U12347 (N_12347,N_10922,N_10557);
nand U12348 (N_12348,N_11788,N_10974);
or U12349 (N_12349,N_10555,N_11946);
or U12350 (N_12350,N_11967,N_10513);
nand U12351 (N_12351,N_11819,N_10797);
xor U12352 (N_12352,N_10520,N_11125);
xnor U12353 (N_12353,N_10793,N_10722);
nand U12354 (N_12354,N_11479,N_11449);
nand U12355 (N_12355,N_11507,N_11423);
nand U12356 (N_12356,N_11758,N_11664);
nand U12357 (N_12357,N_10795,N_10665);
nand U12358 (N_12358,N_10715,N_11929);
nand U12359 (N_12359,N_11326,N_10516);
nand U12360 (N_12360,N_11991,N_10774);
nand U12361 (N_12361,N_11516,N_10613);
nand U12362 (N_12362,N_11690,N_11682);
or U12363 (N_12363,N_10775,N_11671);
xor U12364 (N_12364,N_10944,N_11630);
or U12365 (N_12365,N_11111,N_10720);
nand U12366 (N_12366,N_10725,N_11093);
nand U12367 (N_12367,N_10826,N_11867);
or U12368 (N_12368,N_11220,N_11485);
or U12369 (N_12369,N_10982,N_11706);
nand U12370 (N_12370,N_10994,N_11621);
nand U12371 (N_12371,N_11124,N_11487);
nand U12372 (N_12372,N_10653,N_10585);
xnor U12373 (N_12373,N_11186,N_11661);
nor U12374 (N_12374,N_11592,N_11130);
nand U12375 (N_12375,N_11622,N_11148);
nor U12376 (N_12376,N_10978,N_11725);
nor U12377 (N_12377,N_10777,N_11020);
nand U12378 (N_12378,N_11105,N_11279);
nand U12379 (N_12379,N_10580,N_11410);
nand U12380 (N_12380,N_11930,N_11993);
nor U12381 (N_12381,N_10847,N_11825);
xor U12382 (N_12382,N_11477,N_10864);
and U12383 (N_12383,N_11965,N_10675);
nor U12384 (N_12384,N_11298,N_11846);
or U12385 (N_12385,N_11970,N_10507);
and U12386 (N_12386,N_11652,N_11062);
nor U12387 (N_12387,N_11646,N_11578);
or U12388 (N_12388,N_10607,N_11241);
xor U12389 (N_12389,N_10550,N_11741);
nand U12390 (N_12390,N_10598,N_11707);
or U12391 (N_12391,N_10706,N_11114);
and U12392 (N_12392,N_11200,N_10995);
nor U12393 (N_12393,N_11624,N_10716);
or U12394 (N_12394,N_11445,N_11713);
nand U12395 (N_12395,N_10953,N_10901);
xnor U12396 (N_12396,N_11247,N_10570);
or U12397 (N_12397,N_11284,N_11734);
or U12398 (N_12398,N_11334,N_11753);
and U12399 (N_12399,N_11850,N_11178);
nand U12400 (N_12400,N_10756,N_11494);
nor U12401 (N_12401,N_10956,N_11245);
nor U12402 (N_12402,N_10858,N_11708);
nand U12403 (N_12403,N_11617,N_11604);
or U12404 (N_12404,N_11182,N_11829);
xnor U12405 (N_12405,N_10848,N_11818);
nor U12406 (N_12406,N_11197,N_11989);
or U12407 (N_12407,N_11235,N_11391);
nand U12408 (N_12408,N_11418,N_11812);
or U12409 (N_12409,N_11696,N_10503);
nor U12410 (N_12410,N_11305,N_10673);
nand U12411 (N_12411,N_11329,N_11510);
or U12412 (N_12412,N_11291,N_11415);
and U12413 (N_12413,N_10660,N_10814);
and U12414 (N_12414,N_11172,N_11109);
and U12415 (N_12415,N_11942,N_11133);
or U12416 (N_12416,N_10889,N_11786);
or U12417 (N_12417,N_10854,N_10798);
or U12418 (N_12418,N_10757,N_11957);
or U12419 (N_12419,N_11573,N_11662);
nand U12420 (N_12420,N_11156,N_11985);
or U12421 (N_12421,N_11255,N_11718);
nor U12422 (N_12422,N_11923,N_11057);
and U12423 (N_12423,N_10645,N_11884);
xnor U12424 (N_12424,N_10621,N_11467);
nor U12425 (N_12425,N_11607,N_11129);
nand U12426 (N_12426,N_10800,N_11266);
and U12427 (N_12427,N_10713,N_10837);
nand U12428 (N_12428,N_11359,N_10733);
and U12429 (N_12429,N_11190,N_11465);
nor U12430 (N_12430,N_11009,N_11815);
nand U12431 (N_12431,N_11043,N_11531);
nand U12432 (N_12432,N_11441,N_11357);
nor U12433 (N_12433,N_11538,N_11048);
and U12434 (N_12434,N_10581,N_11321);
or U12435 (N_12435,N_11201,N_11598);
nor U12436 (N_12436,N_10966,N_10684);
xnor U12437 (N_12437,N_11269,N_11503);
nor U12438 (N_12438,N_10532,N_11400);
or U12439 (N_12439,N_11593,N_11723);
and U12440 (N_12440,N_10537,N_11900);
xnor U12441 (N_12441,N_11349,N_11103);
nand U12442 (N_12442,N_10708,N_10698);
nand U12443 (N_12443,N_11439,N_11144);
nand U12444 (N_12444,N_10741,N_10655);
xnor U12445 (N_12445,N_11570,N_11344);
and U12446 (N_12446,N_11339,N_11347);
or U12447 (N_12447,N_10785,N_11853);
or U12448 (N_12448,N_11568,N_11372);
nor U12449 (N_12449,N_11916,N_10783);
nor U12450 (N_12450,N_11513,N_11919);
and U12451 (N_12451,N_11716,N_10938);
and U12452 (N_12452,N_10761,N_11774);
xor U12453 (N_12453,N_11722,N_10699);
nand U12454 (N_12454,N_10630,N_11702);
or U12455 (N_12455,N_10895,N_10554);
and U12456 (N_12456,N_11491,N_11088);
nor U12457 (N_12457,N_11810,N_11290);
nand U12458 (N_12458,N_11230,N_11977);
nor U12459 (N_12459,N_11684,N_11331);
nor U12460 (N_12460,N_11421,N_11459);
and U12461 (N_12461,N_11733,N_11083);
nand U12462 (N_12462,N_10685,N_11142);
or U12463 (N_12463,N_11835,N_11783);
nor U12464 (N_12464,N_11023,N_10856);
nor U12465 (N_12465,N_10765,N_11891);
xor U12466 (N_12466,N_10726,N_10963);
and U12467 (N_12467,N_11257,N_11883);
or U12468 (N_12468,N_10534,N_11013);
nor U12469 (N_12469,N_11994,N_11544);
xnor U12470 (N_12470,N_11068,N_11090);
or U12471 (N_12471,N_10529,N_11362);
nor U12472 (N_12472,N_11424,N_10927);
or U12473 (N_12473,N_11434,N_10983);
and U12474 (N_12474,N_11034,N_11390);
or U12475 (N_12475,N_11555,N_10566);
and U12476 (N_12476,N_11933,N_10948);
and U12477 (N_12477,N_11450,N_10602);
and U12478 (N_12478,N_11087,N_11575);
xor U12479 (N_12479,N_11160,N_11817);
nor U12480 (N_12480,N_11827,N_11502);
nor U12481 (N_12481,N_11340,N_11800);
nand U12482 (N_12482,N_10547,N_11393);
xor U12483 (N_12483,N_11594,N_11258);
and U12484 (N_12484,N_11320,N_11864);
and U12485 (N_12485,N_11042,N_11209);
and U12486 (N_12486,N_11551,N_10530);
and U12487 (N_12487,N_11703,N_11653);
and U12488 (N_12488,N_11222,N_11760);
nor U12489 (N_12489,N_11932,N_11941);
and U12490 (N_12490,N_10680,N_11251);
and U12491 (N_12491,N_10605,N_11655);
nand U12492 (N_12492,N_10674,N_11811);
xor U12493 (N_12493,N_11856,N_11865);
or U12494 (N_12494,N_11830,N_11396);
or U12495 (N_12495,N_10912,N_11925);
or U12496 (N_12496,N_11838,N_10883);
nand U12497 (N_12497,N_11779,N_11162);
nor U12498 (N_12498,N_11577,N_11831);
nor U12499 (N_12499,N_11855,N_10991);
nand U12500 (N_12500,N_11836,N_10707);
nand U12501 (N_12501,N_11003,N_10601);
and U12502 (N_12502,N_10612,N_11757);
nor U12503 (N_12503,N_10627,N_11656);
or U12504 (N_12504,N_11052,N_10764);
and U12505 (N_12505,N_11775,N_10658);
and U12506 (N_12506,N_11744,N_10878);
or U12507 (N_12507,N_10782,N_11496);
and U12508 (N_12508,N_11665,N_11563);
or U12509 (N_12509,N_10961,N_11618);
nand U12510 (N_12510,N_11033,N_10894);
nand U12511 (N_12511,N_11540,N_11806);
or U12512 (N_12512,N_11596,N_10649);
nand U12513 (N_12513,N_11214,N_11237);
and U12514 (N_12514,N_10714,N_10752);
nor U12515 (N_12515,N_11316,N_11537);
and U12516 (N_12516,N_10892,N_10916);
and U12517 (N_12517,N_10917,N_11581);
xnor U12518 (N_12518,N_11054,N_11928);
nor U12519 (N_12519,N_10833,N_11199);
and U12520 (N_12520,N_10887,N_11740);
nand U12521 (N_12521,N_10762,N_10633);
nand U12522 (N_12522,N_11026,N_11134);
and U12523 (N_12523,N_10689,N_11166);
nor U12524 (N_12524,N_11278,N_10682);
or U12525 (N_12525,N_11675,N_11909);
and U12526 (N_12526,N_11343,N_11447);
xor U12527 (N_12527,N_10788,N_11776);
or U12528 (N_12528,N_11146,N_10905);
and U12529 (N_12529,N_10703,N_11429);
and U12530 (N_12530,N_11282,N_11139);
nor U12531 (N_12531,N_11796,N_11309);
and U12532 (N_12532,N_11700,N_11958);
or U12533 (N_12533,N_10584,N_11123);
or U12534 (N_12534,N_11271,N_11517);
nand U12535 (N_12535,N_11277,N_11490);
or U12536 (N_12536,N_10816,N_11324);
nor U12537 (N_12537,N_11590,N_11014);
nand U12538 (N_12538,N_11102,N_11770);
nor U12539 (N_12539,N_11198,N_11681);
and U12540 (N_12540,N_11145,N_11772);
nor U12541 (N_12541,N_10789,N_11385);
or U12542 (N_12542,N_11841,N_11018);
and U12543 (N_12543,N_11137,N_10536);
or U12544 (N_12544,N_10724,N_11854);
nand U12545 (N_12545,N_11202,N_11550);
and U12546 (N_12546,N_11101,N_11376);
nor U12547 (N_12547,N_11603,N_11027);
or U12548 (N_12548,N_11699,N_11526);
or U12549 (N_12549,N_11862,N_11851);
or U12550 (N_12550,N_10750,N_10791);
or U12551 (N_12551,N_11453,N_11822);
or U12552 (N_12552,N_11041,N_10812);
nor U12553 (N_12553,N_11070,N_11461);
nor U12554 (N_12554,N_11229,N_10512);
nor U12555 (N_12555,N_11765,N_11243);
and U12556 (N_12556,N_11174,N_11601);
nand U12557 (N_12557,N_11438,N_11498);
nand U12558 (N_12558,N_10693,N_11782);
or U12559 (N_12559,N_11330,N_11549);
nor U12560 (N_12560,N_11373,N_11626);
and U12561 (N_12561,N_10539,N_10692);
and U12562 (N_12562,N_11519,N_10600);
or U12563 (N_12563,N_10805,N_11920);
nor U12564 (N_12564,N_10965,N_10815);
or U12565 (N_12565,N_10679,N_10770);
nand U12566 (N_12566,N_10641,N_11046);
nor U12567 (N_12567,N_11636,N_11613);
and U12568 (N_12568,N_11196,N_11497);
nor U12569 (N_12569,N_11336,N_11777);
xnor U12570 (N_12570,N_10834,N_11910);
or U12571 (N_12571,N_11599,N_11629);
and U12572 (N_12572,N_11761,N_11369);
xor U12573 (N_12573,N_11007,N_11167);
and U12574 (N_12574,N_11902,N_10710);
xor U12575 (N_12575,N_11844,N_11663);
nand U12576 (N_12576,N_11419,N_10973);
or U12577 (N_12577,N_11475,N_10936);
and U12578 (N_12578,N_10632,N_11095);
nand U12579 (N_12579,N_10841,N_10926);
xor U12580 (N_12580,N_11605,N_10799);
and U12581 (N_12581,N_10661,N_11802);
nand U12582 (N_12582,N_11311,N_10952);
xnor U12583 (N_12583,N_10515,N_10968);
or U12584 (N_12584,N_11562,N_11731);
nor U12585 (N_12585,N_10957,N_11673);
and U12586 (N_12586,N_10990,N_11816);
xor U12587 (N_12587,N_11318,N_10962);
or U12588 (N_12588,N_11300,N_10802);
and U12589 (N_12589,N_11500,N_10610);
and U12590 (N_12590,N_10747,N_11379);
nand U12591 (N_12591,N_11367,N_11384);
or U12592 (N_12592,N_11161,N_11969);
nand U12593 (N_12593,N_10943,N_11187);
nand U12594 (N_12594,N_11536,N_11695);
nand U12595 (N_12595,N_11482,N_11021);
nor U12596 (N_12596,N_11096,N_11763);
nand U12597 (N_12597,N_11375,N_11797);
nor U12598 (N_12598,N_11306,N_11059);
and U12599 (N_12599,N_11121,N_10825);
or U12600 (N_12600,N_11845,N_11508);
and U12601 (N_12601,N_11738,N_10551);
xor U12602 (N_12602,N_11821,N_11576);
nand U12603 (N_12603,N_11554,N_11356);
xor U12604 (N_12604,N_10712,N_10736);
or U12605 (N_12605,N_11720,N_10595);
or U12606 (N_12606,N_11975,N_10688);
nand U12607 (N_12607,N_11728,N_10870);
nor U12608 (N_12608,N_11943,N_11742);
nand U12609 (N_12609,N_11351,N_11732);
and U12610 (N_12610,N_11896,N_10860);
nor U12611 (N_12611,N_11642,N_11411);
and U12612 (N_12612,N_10634,N_11640);
xnor U12613 (N_12613,N_11814,N_11893);
or U12614 (N_12614,N_10852,N_11952);
or U12615 (N_12615,N_11698,N_10567);
nor U12616 (N_12616,N_11228,N_10898);
and U12617 (N_12617,N_11704,N_11632);
nor U12618 (N_12618,N_11010,N_11591);
and U12619 (N_12619,N_11529,N_11260);
xor U12620 (N_12620,N_11543,N_11501);
or U12621 (N_12621,N_11422,N_10666);
or U12622 (N_12622,N_11071,N_10608);
nor U12623 (N_12623,N_11004,N_11051);
or U12624 (N_12624,N_10820,N_11651);
nand U12625 (N_12625,N_11755,N_10768);
and U12626 (N_12626,N_11914,N_11355);
or U12627 (N_12627,N_10946,N_10611);
nor U12628 (N_12628,N_11165,N_10790);
xor U12629 (N_12629,N_11177,N_11499);
nand U12630 (N_12630,N_11687,N_10821);
nand U12631 (N_12631,N_11614,N_10969);
nor U12632 (N_12632,N_10694,N_11504);
and U12633 (N_12633,N_11184,N_10937);
and U12634 (N_12634,N_10552,N_11313);
and U12635 (N_12635,N_10690,N_11478);
nor U12636 (N_12636,N_10582,N_10906);
or U12637 (N_12637,N_11886,N_11863);
and U12638 (N_12638,N_11006,N_11413);
and U12639 (N_12639,N_10960,N_11470);
nand U12640 (N_12640,N_11236,N_10521);
nand U12641 (N_12641,N_11000,N_10818);
nand U12642 (N_12642,N_11098,N_11637);
nand U12643 (N_12643,N_11964,N_11402);
or U12644 (N_12644,N_10859,N_10506);
or U12645 (N_12645,N_11240,N_11256);
and U12646 (N_12646,N_11960,N_10523);
nor U12647 (N_12647,N_11754,N_11454);
nand U12648 (N_12648,N_10808,N_11717);
or U12649 (N_12649,N_10862,N_11709);
nor U12650 (N_12650,N_11749,N_11074);
nor U12651 (N_12651,N_11881,N_10544);
nand U12652 (N_12652,N_11894,N_11746);
and U12653 (N_12653,N_11012,N_10866);
nand U12654 (N_12654,N_11154,N_11931);
xor U12655 (N_12655,N_11079,N_10729);
nor U12656 (N_12656,N_10967,N_11407);
nor U12657 (N_12657,N_11807,N_11299);
nand U12658 (N_12658,N_11769,N_11926);
nand U12659 (N_12659,N_11354,N_11066);
nor U12660 (N_12660,N_10766,N_10839);
or U12661 (N_12661,N_11524,N_10970);
nor U12662 (N_12662,N_11296,N_11678);
nor U12663 (N_12663,N_10996,N_11140);
nand U12664 (N_12664,N_11374,N_11565);
xor U12665 (N_12665,N_11471,N_10773);
nor U12666 (N_12666,N_11312,N_10654);
or U12667 (N_12667,N_11293,N_11778);
nand U12668 (N_12668,N_11619,N_11804);
and U12669 (N_12669,N_11120,N_11692);
or U12670 (N_12670,N_11169,N_10909);
or U12671 (N_12671,N_10524,N_10740);
nand U12672 (N_12672,N_11541,N_11116);
nand U12673 (N_12673,N_11648,N_10719);
xor U12674 (N_12674,N_11432,N_11547);
nand U12675 (N_12675,N_10897,N_10947);
nand U12676 (N_12676,N_11938,N_11159);
nor U12677 (N_12677,N_11317,N_11956);
or U12678 (N_12678,N_11352,N_11885);
or U12679 (N_12679,N_11158,N_10877);
or U12680 (N_12680,N_11099,N_11995);
xor U12681 (N_12681,N_11468,N_10853);
or U12682 (N_12682,N_10670,N_11037);
nor U12683 (N_12683,N_11086,N_10676);
nand U12684 (N_12684,N_10941,N_11697);
and U12685 (N_12685,N_10609,N_11303);
nand U12686 (N_12686,N_10659,N_10874);
and U12687 (N_12687,N_11608,N_10872);
and U12688 (N_12688,N_10742,N_11974);
and U12689 (N_12689,N_10840,N_10890);
and U12690 (N_12690,N_10501,N_11113);
nand U12691 (N_12691,N_11907,N_11346);
xnor U12692 (N_12692,N_11586,N_11918);
or U12693 (N_12693,N_11666,N_11582);
nand U12694 (N_12694,N_11325,N_10522);
and U12695 (N_12695,N_11828,N_10728);
nand U12696 (N_12696,N_11870,N_10855);
nand U12697 (N_12697,N_10511,N_11170);
or U12698 (N_12698,N_10545,N_11463);
nor U12699 (N_12699,N_11061,N_10951);
or U12700 (N_12700,N_11446,N_11824);
or U12701 (N_12701,N_10763,N_11711);
xor U12702 (N_12702,N_11078,N_11674);
nor U12703 (N_12703,N_11972,N_11019);
nor U12704 (N_12704,N_10628,N_10850);
xnor U12705 (N_12705,N_11762,N_10635);
nor U12706 (N_12706,N_11350,N_11625);
nand U12707 (N_12707,N_10986,N_10681);
nor U12708 (N_12708,N_10780,N_11557);
xnor U12709 (N_12709,N_10517,N_10652);
nor U12710 (N_12710,N_11383,N_11388);
nand U12711 (N_12711,N_11984,N_10615);
nand U12712 (N_12712,N_11377,N_11430);
nand U12713 (N_12713,N_11620,N_11944);
nor U12714 (N_12714,N_10811,N_10622);
or U12715 (N_12715,N_11951,N_11094);
or U12716 (N_12716,N_10942,N_11412);
and U12717 (N_12717,N_11118,N_11635);
and U12718 (N_12718,N_10801,N_11976);
or U12719 (N_12719,N_10828,N_10683);
and U12720 (N_12720,N_11185,N_11615);
and U12721 (N_12721,N_11668,N_11211);
nand U12722 (N_12722,N_11729,N_10914);
nor U12723 (N_12723,N_11911,N_11878);
or U12724 (N_12724,N_10923,N_10993);
nor U12725 (N_12725,N_11627,N_11654);
nand U12726 (N_12726,N_10672,N_11523);
nor U12727 (N_12727,N_11226,N_10702);
xnor U12728 (N_12728,N_11739,N_11225);
nand U12729 (N_12729,N_11307,N_11908);
or U12730 (N_12730,N_11248,N_11506);
and U12731 (N_12731,N_11848,N_11163);
and U12732 (N_12732,N_11428,N_11660);
or U12733 (N_12733,N_10810,N_10597);
nand U12734 (N_12734,N_11623,N_11193);
or U12735 (N_12735,N_10638,N_11106);
and U12736 (N_12736,N_10730,N_11030);
or U12737 (N_12737,N_10743,N_11370);
nand U12738 (N_12738,N_11552,N_11112);
or U12739 (N_12739,N_11647,N_11232);
and U12740 (N_12740,N_11348,N_11514);
nor U12741 (N_12741,N_11784,N_11205);
or U12742 (N_12742,N_11553,N_11645);
and U12743 (N_12743,N_11031,N_11280);
nor U12744 (N_12744,N_11609,N_10964);
or U12745 (N_12745,N_10827,N_11945);
or U12746 (N_12746,N_11416,N_11025);
nor U12747 (N_12747,N_11341,N_11085);
or U12748 (N_12748,N_11420,N_11589);
or U12749 (N_12749,N_11458,N_11015);
nand U12750 (N_12750,N_11413,N_11243);
and U12751 (N_12751,N_11454,N_10769);
and U12752 (N_12752,N_10707,N_11431);
and U12753 (N_12753,N_11680,N_11119);
nor U12754 (N_12754,N_10943,N_10655);
or U12755 (N_12755,N_10589,N_11847);
nand U12756 (N_12756,N_11614,N_11073);
or U12757 (N_12757,N_11585,N_10709);
xor U12758 (N_12758,N_11205,N_10569);
and U12759 (N_12759,N_11627,N_10985);
nand U12760 (N_12760,N_11891,N_10955);
nand U12761 (N_12761,N_11417,N_10857);
or U12762 (N_12762,N_10662,N_11417);
and U12763 (N_12763,N_11688,N_11509);
nand U12764 (N_12764,N_11265,N_11836);
or U12765 (N_12765,N_11499,N_11126);
or U12766 (N_12766,N_11189,N_10917);
and U12767 (N_12767,N_11128,N_11268);
nor U12768 (N_12768,N_10809,N_10673);
and U12769 (N_12769,N_11309,N_11242);
and U12770 (N_12770,N_11286,N_11146);
or U12771 (N_12771,N_11496,N_10655);
xor U12772 (N_12772,N_10505,N_11096);
nand U12773 (N_12773,N_11960,N_11742);
and U12774 (N_12774,N_11236,N_11080);
and U12775 (N_12775,N_11232,N_11659);
nand U12776 (N_12776,N_10753,N_10935);
nor U12777 (N_12777,N_11093,N_11931);
and U12778 (N_12778,N_10662,N_11203);
nor U12779 (N_12779,N_11299,N_11888);
or U12780 (N_12780,N_11246,N_10858);
or U12781 (N_12781,N_10550,N_10561);
nand U12782 (N_12782,N_11066,N_11603);
nand U12783 (N_12783,N_11961,N_11628);
and U12784 (N_12784,N_11858,N_11105);
xor U12785 (N_12785,N_10703,N_11398);
nand U12786 (N_12786,N_11738,N_11795);
and U12787 (N_12787,N_11094,N_10839);
or U12788 (N_12788,N_10700,N_10630);
nor U12789 (N_12789,N_11865,N_10819);
nor U12790 (N_12790,N_11608,N_10664);
or U12791 (N_12791,N_11607,N_11646);
or U12792 (N_12792,N_11572,N_11379);
and U12793 (N_12793,N_11160,N_11714);
nand U12794 (N_12794,N_10613,N_11019);
nor U12795 (N_12795,N_11665,N_11383);
and U12796 (N_12796,N_10640,N_11298);
or U12797 (N_12797,N_10575,N_11892);
nand U12798 (N_12798,N_11704,N_11858);
or U12799 (N_12799,N_11306,N_11819);
nand U12800 (N_12800,N_11717,N_11776);
xor U12801 (N_12801,N_11991,N_11368);
nor U12802 (N_12802,N_10809,N_11673);
and U12803 (N_12803,N_10754,N_11179);
or U12804 (N_12804,N_11864,N_10972);
nor U12805 (N_12805,N_10955,N_10678);
nand U12806 (N_12806,N_11883,N_10813);
or U12807 (N_12807,N_10835,N_11006);
or U12808 (N_12808,N_11539,N_11293);
or U12809 (N_12809,N_10634,N_10713);
and U12810 (N_12810,N_10576,N_11546);
nand U12811 (N_12811,N_11340,N_11909);
and U12812 (N_12812,N_10573,N_11334);
nand U12813 (N_12813,N_10615,N_11681);
xnor U12814 (N_12814,N_10557,N_11932);
and U12815 (N_12815,N_11509,N_10750);
and U12816 (N_12816,N_11407,N_11262);
and U12817 (N_12817,N_11765,N_11187);
or U12818 (N_12818,N_11332,N_11225);
or U12819 (N_12819,N_11163,N_10863);
nand U12820 (N_12820,N_11601,N_10554);
and U12821 (N_12821,N_10846,N_11836);
nand U12822 (N_12822,N_11550,N_11260);
nand U12823 (N_12823,N_10605,N_11020);
and U12824 (N_12824,N_11849,N_10634);
and U12825 (N_12825,N_11092,N_10547);
nand U12826 (N_12826,N_11735,N_10906);
nor U12827 (N_12827,N_10980,N_11876);
and U12828 (N_12828,N_11437,N_11849);
or U12829 (N_12829,N_10686,N_11614);
nand U12830 (N_12830,N_11565,N_11979);
nor U12831 (N_12831,N_11492,N_11888);
or U12832 (N_12832,N_11501,N_11840);
nor U12833 (N_12833,N_11725,N_11011);
nand U12834 (N_12834,N_11381,N_11213);
or U12835 (N_12835,N_10969,N_11655);
or U12836 (N_12836,N_11794,N_11666);
or U12837 (N_12837,N_10880,N_11155);
xor U12838 (N_12838,N_11816,N_11466);
or U12839 (N_12839,N_10801,N_11941);
and U12840 (N_12840,N_10825,N_11914);
and U12841 (N_12841,N_11742,N_11167);
and U12842 (N_12842,N_11410,N_10626);
or U12843 (N_12843,N_10748,N_10500);
or U12844 (N_12844,N_10594,N_11203);
nor U12845 (N_12845,N_11562,N_11433);
nor U12846 (N_12846,N_11010,N_11863);
nor U12847 (N_12847,N_10691,N_11628);
and U12848 (N_12848,N_11604,N_10964);
or U12849 (N_12849,N_11226,N_10636);
and U12850 (N_12850,N_11417,N_10793);
nand U12851 (N_12851,N_11627,N_11680);
or U12852 (N_12852,N_11004,N_11324);
and U12853 (N_12853,N_11470,N_10813);
nor U12854 (N_12854,N_10977,N_11277);
nand U12855 (N_12855,N_11076,N_11069);
nor U12856 (N_12856,N_10627,N_11980);
xor U12857 (N_12857,N_11590,N_11748);
and U12858 (N_12858,N_11535,N_10509);
and U12859 (N_12859,N_10912,N_11423);
and U12860 (N_12860,N_10666,N_10793);
and U12861 (N_12861,N_10776,N_10880);
and U12862 (N_12862,N_11833,N_11504);
or U12863 (N_12863,N_11212,N_11647);
nor U12864 (N_12864,N_11182,N_11434);
or U12865 (N_12865,N_11200,N_11030);
and U12866 (N_12866,N_10733,N_10985);
nand U12867 (N_12867,N_11344,N_10991);
and U12868 (N_12868,N_10651,N_11326);
or U12869 (N_12869,N_11329,N_11109);
and U12870 (N_12870,N_11340,N_10709);
nor U12871 (N_12871,N_10664,N_11909);
or U12872 (N_12872,N_10820,N_10994);
nor U12873 (N_12873,N_11963,N_10686);
nand U12874 (N_12874,N_11659,N_11463);
and U12875 (N_12875,N_10793,N_10712);
or U12876 (N_12876,N_11305,N_10780);
xnor U12877 (N_12877,N_11673,N_11081);
or U12878 (N_12878,N_11048,N_11130);
and U12879 (N_12879,N_10954,N_11063);
and U12880 (N_12880,N_11310,N_10916);
and U12881 (N_12881,N_11269,N_10860);
or U12882 (N_12882,N_11875,N_10699);
and U12883 (N_12883,N_11704,N_11735);
and U12884 (N_12884,N_11977,N_10722);
nand U12885 (N_12885,N_11299,N_10522);
nand U12886 (N_12886,N_11409,N_11063);
xnor U12887 (N_12887,N_10981,N_11187);
nor U12888 (N_12888,N_11542,N_11520);
nand U12889 (N_12889,N_11937,N_11338);
xor U12890 (N_12890,N_11223,N_10656);
and U12891 (N_12891,N_11558,N_11922);
nor U12892 (N_12892,N_11215,N_11817);
nand U12893 (N_12893,N_10634,N_11907);
nor U12894 (N_12894,N_10526,N_11283);
nand U12895 (N_12895,N_11318,N_11198);
and U12896 (N_12896,N_11905,N_10779);
or U12897 (N_12897,N_10979,N_11662);
and U12898 (N_12898,N_11787,N_10829);
and U12899 (N_12899,N_11235,N_11819);
or U12900 (N_12900,N_11981,N_10868);
or U12901 (N_12901,N_11819,N_11618);
nand U12902 (N_12902,N_11151,N_10726);
nand U12903 (N_12903,N_11823,N_10595);
xor U12904 (N_12904,N_11168,N_11613);
nor U12905 (N_12905,N_11251,N_11800);
or U12906 (N_12906,N_11880,N_10938);
or U12907 (N_12907,N_11994,N_11020);
and U12908 (N_12908,N_10501,N_10953);
and U12909 (N_12909,N_10668,N_10736);
nor U12910 (N_12910,N_11717,N_11184);
or U12911 (N_12911,N_10642,N_11222);
nor U12912 (N_12912,N_10717,N_10660);
nor U12913 (N_12913,N_11604,N_11124);
nand U12914 (N_12914,N_10908,N_11461);
nor U12915 (N_12915,N_11388,N_10501);
and U12916 (N_12916,N_11496,N_10663);
and U12917 (N_12917,N_10659,N_11414);
and U12918 (N_12918,N_10664,N_11798);
xnor U12919 (N_12919,N_10941,N_10823);
or U12920 (N_12920,N_11684,N_10734);
nor U12921 (N_12921,N_10533,N_11901);
or U12922 (N_12922,N_10565,N_10800);
xor U12923 (N_12923,N_11917,N_11715);
nor U12924 (N_12924,N_11333,N_11409);
and U12925 (N_12925,N_10610,N_11659);
or U12926 (N_12926,N_11794,N_10552);
and U12927 (N_12927,N_11649,N_11105);
nand U12928 (N_12928,N_10867,N_10961);
nor U12929 (N_12929,N_11982,N_10578);
nand U12930 (N_12930,N_11030,N_11395);
or U12931 (N_12931,N_11485,N_11556);
and U12932 (N_12932,N_10756,N_11033);
nor U12933 (N_12933,N_11995,N_10783);
xnor U12934 (N_12934,N_10721,N_11805);
and U12935 (N_12935,N_11805,N_10725);
and U12936 (N_12936,N_11432,N_11247);
nand U12937 (N_12937,N_11473,N_11133);
nor U12938 (N_12938,N_11885,N_11671);
and U12939 (N_12939,N_11060,N_11551);
or U12940 (N_12940,N_11024,N_10681);
nor U12941 (N_12941,N_10804,N_10598);
nor U12942 (N_12942,N_11167,N_10509);
and U12943 (N_12943,N_11673,N_10766);
nand U12944 (N_12944,N_11927,N_11480);
nand U12945 (N_12945,N_10616,N_10877);
nand U12946 (N_12946,N_11443,N_10809);
and U12947 (N_12947,N_11763,N_11409);
nand U12948 (N_12948,N_11953,N_11922);
or U12949 (N_12949,N_10548,N_11642);
and U12950 (N_12950,N_11620,N_10810);
nor U12951 (N_12951,N_11100,N_11837);
nand U12952 (N_12952,N_10635,N_11266);
or U12953 (N_12953,N_10776,N_11490);
or U12954 (N_12954,N_10667,N_11086);
nor U12955 (N_12955,N_11881,N_11631);
or U12956 (N_12956,N_11397,N_10815);
or U12957 (N_12957,N_11733,N_11314);
or U12958 (N_12958,N_11539,N_11571);
nor U12959 (N_12959,N_11689,N_11159);
or U12960 (N_12960,N_10511,N_11451);
and U12961 (N_12961,N_10983,N_10964);
nor U12962 (N_12962,N_11121,N_10607);
nand U12963 (N_12963,N_10813,N_11549);
xor U12964 (N_12964,N_11550,N_11429);
and U12965 (N_12965,N_11605,N_11916);
nor U12966 (N_12966,N_11365,N_11997);
nor U12967 (N_12967,N_11293,N_10637);
xor U12968 (N_12968,N_11077,N_10503);
nand U12969 (N_12969,N_11795,N_10977);
nor U12970 (N_12970,N_11445,N_11092);
nor U12971 (N_12971,N_11624,N_11623);
nand U12972 (N_12972,N_11367,N_11593);
and U12973 (N_12973,N_10691,N_10604);
nor U12974 (N_12974,N_11824,N_10736);
or U12975 (N_12975,N_10516,N_11358);
nand U12976 (N_12976,N_11282,N_10777);
nor U12977 (N_12977,N_11487,N_11478);
nor U12978 (N_12978,N_11829,N_10583);
nor U12979 (N_12979,N_11972,N_11925);
nor U12980 (N_12980,N_11279,N_11721);
and U12981 (N_12981,N_11676,N_11299);
nor U12982 (N_12982,N_10662,N_11147);
or U12983 (N_12983,N_11721,N_11002);
nor U12984 (N_12984,N_11801,N_10623);
and U12985 (N_12985,N_11757,N_11762);
and U12986 (N_12986,N_11393,N_11881);
and U12987 (N_12987,N_11154,N_11921);
nor U12988 (N_12988,N_10719,N_11642);
and U12989 (N_12989,N_11684,N_11256);
nor U12990 (N_12990,N_11846,N_11760);
xnor U12991 (N_12991,N_11486,N_11425);
xor U12992 (N_12992,N_11757,N_11773);
or U12993 (N_12993,N_11537,N_11152);
nor U12994 (N_12994,N_10591,N_10818);
nor U12995 (N_12995,N_11258,N_11147);
nand U12996 (N_12996,N_10729,N_10619);
and U12997 (N_12997,N_11856,N_10841);
and U12998 (N_12998,N_10753,N_10694);
nand U12999 (N_12999,N_10869,N_10666);
or U13000 (N_13000,N_10816,N_11890);
or U13001 (N_13001,N_11556,N_11318);
nor U13002 (N_13002,N_11382,N_11901);
and U13003 (N_13003,N_11289,N_10767);
nor U13004 (N_13004,N_10747,N_11555);
xor U13005 (N_13005,N_11920,N_10714);
nor U13006 (N_13006,N_11583,N_11428);
or U13007 (N_13007,N_11919,N_10784);
nor U13008 (N_13008,N_11096,N_10847);
and U13009 (N_13009,N_11095,N_10620);
and U13010 (N_13010,N_11302,N_11680);
xor U13011 (N_13011,N_11780,N_11012);
nand U13012 (N_13012,N_11813,N_11546);
nor U13013 (N_13013,N_10564,N_11442);
xnor U13014 (N_13014,N_11749,N_10893);
nand U13015 (N_13015,N_11183,N_10711);
nand U13016 (N_13016,N_11171,N_11154);
or U13017 (N_13017,N_10530,N_11333);
or U13018 (N_13018,N_11528,N_11617);
or U13019 (N_13019,N_10612,N_10592);
and U13020 (N_13020,N_10725,N_10867);
nor U13021 (N_13021,N_11767,N_10726);
nor U13022 (N_13022,N_11855,N_11316);
or U13023 (N_13023,N_10649,N_11941);
or U13024 (N_13024,N_10524,N_11531);
nand U13025 (N_13025,N_11500,N_11383);
nand U13026 (N_13026,N_11257,N_10577);
nor U13027 (N_13027,N_11940,N_11817);
nand U13028 (N_13028,N_10889,N_11527);
or U13029 (N_13029,N_11453,N_10862);
nor U13030 (N_13030,N_10860,N_11013);
and U13031 (N_13031,N_10662,N_11981);
nand U13032 (N_13032,N_11667,N_10582);
and U13033 (N_13033,N_11799,N_11021);
nand U13034 (N_13034,N_11507,N_11918);
and U13035 (N_13035,N_11823,N_11258);
nor U13036 (N_13036,N_11364,N_10510);
nor U13037 (N_13037,N_11769,N_11020);
nand U13038 (N_13038,N_11921,N_11381);
nand U13039 (N_13039,N_10747,N_10914);
xnor U13040 (N_13040,N_10567,N_11147);
and U13041 (N_13041,N_11013,N_11087);
nand U13042 (N_13042,N_11943,N_11799);
nor U13043 (N_13043,N_11774,N_11228);
nor U13044 (N_13044,N_11659,N_11425);
or U13045 (N_13045,N_11645,N_11987);
or U13046 (N_13046,N_11294,N_11496);
or U13047 (N_13047,N_11962,N_11122);
or U13048 (N_13048,N_11560,N_11590);
nor U13049 (N_13049,N_10539,N_11812);
nand U13050 (N_13050,N_11156,N_11244);
nand U13051 (N_13051,N_11564,N_10803);
nand U13052 (N_13052,N_11727,N_10834);
or U13053 (N_13053,N_11169,N_11262);
nor U13054 (N_13054,N_11090,N_10954);
nor U13055 (N_13055,N_11913,N_11791);
and U13056 (N_13056,N_10721,N_10889);
xor U13057 (N_13057,N_10758,N_11167);
and U13058 (N_13058,N_11181,N_10780);
and U13059 (N_13059,N_11775,N_10578);
or U13060 (N_13060,N_11020,N_10678);
or U13061 (N_13061,N_11379,N_11625);
nor U13062 (N_13062,N_10886,N_11624);
nand U13063 (N_13063,N_10658,N_11097);
or U13064 (N_13064,N_11376,N_10658);
or U13065 (N_13065,N_10550,N_10889);
nand U13066 (N_13066,N_11764,N_11768);
nand U13067 (N_13067,N_11468,N_10697);
nand U13068 (N_13068,N_11634,N_11278);
xnor U13069 (N_13069,N_11356,N_10703);
nor U13070 (N_13070,N_10847,N_10542);
nand U13071 (N_13071,N_11542,N_11540);
or U13072 (N_13072,N_11381,N_11726);
nand U13073 (N_13073,N_11437,N_11376);
nor U13074 (N_13074,N_11553,N_10663);
or U13075 (N_13075,N_11850,N_11629);
and U13076 (N_13076,N_11251,N_10903);
or U13077 (N_13077,N_10767,N_10715);
or U13078 (N_13078,N_11101,N_11676);
or U13079 (N_13079,N_10986,N_11596);
and U13080 (N_13080,N_11015,N_10903);
nand U13081 (N_13081,N_11566,N_10902);
nor U13082 (N_13082,N_11829,N_10653);
nor U13083 (N_13083,N_10906,N_11187);
nor U13084 (N_13084,N_11017,N_10631);
and U13085 (N_13085,N_11202,N_11094);
nor U13086 (N_13086,N_10954,N_11286);
nand U13087 (N_13087,N_10967,N_11958);
nor U13088 (N_13088,N_10507,N_10952);
nor U13089 (N_13089,N_11356,N_10535);
or U13090 (N_13090,N_10746,N_11105);
nor U13091 (N_13091,N_11481,N_11157);
nand U13092 (N_13092,N_11019,N_11877);
or U13093 (N_13093,N_10991,N_11106);
xnor U13094 (N_13094,N_10912,N_11157);
and U13095 (N_13095,N_11807,N_10507);
nand U13096 (N_13096,N_11572,N_11653);
or U13097 (N_13097,N_11941,N_11951);
or U13098 (N_13098,N_10723,N_10558);
nand U13099 (N_13099,N_11512,N_11903);
nor U13100 (N_13100,N_10696,N_11482);
nand U13101 (N_13101,N_11345,N_10815);
nand U13102 (N_13102,N_11486,N_11956);
nor U13103 (N_13103,N_10833,N_11352);
xnor U13104 (N_13104,N_11980,N_11307);
nor U13105 (N_13105,N_11824,N_11104);
nor U13106 (N_13106,N_11249,N_10622);
and U13107 (N_13107,N_11192,N_10772);
and U13108 (N_13108,N_11343,N_10727);
nand U13109 (N_13109,N_11286,N_10610);
nor U13110 (N_13110,N_11416,N_11009);
nor U13111 (N_13111,N_10792,N_11357);
nor U13112 (N_13112,N_11075,N_11598);
and U13113 (N_13113,N_11449,N_11611);
nand U13114 (N_13114,N_11429,N_11114);
nor U13115 (N_13115,N_11824,N_11131);
nand U13116 (N_13116,N_11215,N_11776);
nand U13117 (N_13117,N_11056,N_11115);
or U13118 (N_13118,N_11921,N_10898);
xor U13119 (N_13119,N_10919,N_10640);
and U13120 (N_13120,N_10666,N_11836);
or U13121 (N_13121,N_11397,N_11911);
or U13122 (N_13122,N_11569,N_10966);
nand U13123 (N_13123,N_11784,N_11157);
nand U13124 (N_13124,N_10991,N_10624);
and U13125 (N_13125,N_11174,N_10974);
nand U13126 (N_13126,N_11308,N_11980);
nand U13127 (N_13127,N_11655,N_10533);
and U13128 (N_13128,N_11413,N_11343);
or U13129 (N_13129,N_11399,N_10609);
nor U13130 (N_13130,N_11897,N_11976);
and U13131 (N_13131,N_11948,N_11958);
nor U13132 (N_13132,N_11258,N_10891);
nand U13133 (N_13133,N_11654,N_10858);
and U13134 (N_13134,N_11682,N_11924);
xor U13135 (N_13135,N_11170,N_10784);
and U13136 (N_13136,N_11361,N_11006);
or U13137 (N_13137,N_11398,N_11553);
nand U13138 (N_13138,N_10980,N_10927);
nor U13139 (N_13139,N_11547,N_11932);
or U13140 (N_13140,N_11502,N_11664);
or U13141 (N_13141,N_11281,N_11289);
and U13142 (N_13142,N_11650,N_10898);
xnor U13143 (N_13143,N_11558,N_11203);
nand U13144 (N_13144,N_11522,N_11316);
nor U13145 (N_13145,N_10510,N_11934);
xnor U13146 (N_13146,N_11320,N_11617);
and U13147 (N_13147,N_11497,N_10959);
or U13148 (N_13148,N_11165,N_11364);
xor U13149 (N_13149,N_11545,N_11433);
xnor U13150 (N_13150,N_10730,N_11351);
and U13151 (N_13151,N_10879,N_11074);
nor U13152 (N_13152,N_11174,N_11004);
and U13153 (N_13153,N_11871,N_11433);
and U13154 (N_13154,N_11072,N_11225);
or U13155 (N_13155,N_10930,N_11700);
or U13156 (N_13156,N_11781,N_10593);
nor U13157 (N_13157,N_11674,N_10708);
and U13158 (N_13158,N_10609,N_11843);
or U13159 (N_13159,N_10806,N_11877);
nand U13160 (N_13160,N_11689,N_10927);
nand U13161 (N_13161,N_11744,N_10827);
xor U13162 (N_13162,N_11171,N_11855);
and U13163 (N_13163,N_10869,N_11477);
and U13164 (N_13164,N_11033,N_11816);
xnor U13165 (N_13165,N_10689,N_11621);
nor U13166 (N_13166,N_10586,N_11828);
nor U13167 (N_13167,N_10939,N_11791);
and U13168 (N_13168,N_11381,N_10839);
nand U13169 (N_13169,N_11864,N_10935);
nand U13170 (N_13170,N_11746,N_11111);
and U13171 (N_13171,N_10869,N_10511);
and U13172 (N_13172,N_11131,N_11315);
nor U13173 (N_13173,N_11558,N_10939);
nand U13174 (N_13174,N_11071,N_11443);
nor U13175 (N_13175,N_11289,N_11984);
and U13176 (N_13176,N_10986,N_11864);
nor U13177 (N_13177,N_11056,N_11783);
and U13178 (N_13178,N_11671,N_11972);
nand U13179 (N_13179,N_11543,N_10907);
or U13180 (N_13180,N_10653,N_11894);
nor U13181 (N_13181,N_11822,N_11143);
xnor U13182 (N_13182,N_11609,N_11387);
xnor U13183 (N_13183,N_10752,N_11332);
and U13184 (N_13184,N_11849,N_11963);
and U13185 (N_13185,N_11674,N_11986);
and U13186 (N_13186,N_11923,N_11017);
and U13187 (N_13187,N_11909,N_11653);
nor U13188 (N_13188,N_11632,N_10940);
nand U13189 (N_13189,N_10859,N_11105);
nor U13190 (N_13190,N_11740,N_11327);
nor U13191 (N_13191,N_11138,N_11270);
nor U13192 (N_13192,N_10802,N_11091);
or U13193 (N_13193,N_11620,N_11237);
nand U13194 (N_13194,N_10894,N_11281);
nand U13195 (N_13195,N_10747,N_11419);
nand U13196 (N_13196,N_11526,N_11343);
and U13197 (N_13197,N_10642,N_11588);
nor U13198 (N_13198,N_11194,N_11428);
or U13199 (N_13199,N_11196,N_11631);
nor U13200 (N_13200,N_10954,N_11941);
nor U13201 (N_13201,N_11523,N_10631);
nand U13202 (N_13202,N_11682,N_10836);
or U13203 (N_13203,N_11955,N_10547);
nand U13204 (N_13204,N_10605,N_10729);
or U13205 (N_13205,N_11657,N_10559);
nand U13206 (N_13206,N_10958,N_10847);
and U13207 (N_13207,N_11832,N_11362);
and U13208 (N_13208,N_10836,N_10859);
and U13209 (N_13209,N_11280,N_11505);
or U13210 (N_13210,N_10661,N_10649);
xor U13211 (N_13211,N_11798,N_11705);
nand U13212 (N_13212,N_11815,N_10577);
nand U13213 (N_13213,N_10941,N_11000);
or U13214 (N_13214,N_11240,N_10570);
and U13215 (N_13215,N_11102,N_11827);
xnor U13216 (N_13216,N_11731,N_10824);
nand U13217 (N_13217,N_10529,N_11454);
xnor U13218 (N_13218,N_11868,N_11779);
and U13219 (N_13219,N_11133,N_10796);
xnor U13220 (N_13220,N_11422,N_10955);
or U13221 (N_13221,N_11555,N_11976);
or U13222 (N_13222,N_11289,N_11614);
nor U13223 (N_13223,N_11568,N_11271);
or U13224 (N_13224,N_11290,N_11477);
nor U13225 (N_13225,N_10896,N_11336);
nor U13226 (N_13226,N_11885,N_11041);
nor U13227 (N_13227,N_10655,N_11061);
or U13228 (N_13228,N_11525,N_11386);
or U13229 (N_13229,N_10502,N_11163);
nor U13230 (N_13230,N_11010,N_11208);
nand U13231 (N_13231,N_11185,N_11462);
and U13232 (N_13232,N_11633,N_10791);
or U13233 (N_13233,N_11457,N_11709);
nor U13234 (N_13234,N_10974,N_10636);
or U13235 (N_13235,N_11245,N_11638);
or U13236 (N_13236,N_10780,N_10522);
nor U13237 (N_13237,N_11792,N_10939);
nor U13238 (N_13238,N_11121,N_11764);
or U13239 (N_13239,N_11554,N_10508);
nand U13240 (N_13240,N_11059,N_11461);
nor U13241 (N_13241,N_11579,N_10593);
nor U13242 (N_13242,N_10584,N_10841);
or U13243 (N_13243,N_11481,N_11631);
and U13244 (N_13244,N_11242,N_11263);
or U13245 (N_13245,N_11905,N_11693);
and U13246 (N_13246,N_11151,N_11423);
xnor U13247 (N_13247,N_10810,N_10629);
or U13248 (N_13248,N_11192,N_11346);
nand U13249 (N_13249,N_11792,N_10545);
nor U13250 (N_13250,N_11283,N_11499);
nor U13251 (N_13251,N_11752,N_11736);
nand U13252 (N_13252,N_11834,N_11870);
or U13253 (N_13253,N_11792,N_10869);
nand U13254 (N_13254,N_11602,N_10526);
nand U13255 (N_13255,N_11713,N_10756);
and U13256 (N_13256,N_11840,N_11363);
nor U13257 (N_13257,N_10930,N_10666);
or U13258 (N_13258,N_11582,N_10980);
nand U13259 (N_13259,N_11611,N_10574);
nor U13260 (N_13260,N_10880,N_11338);
xor U13261 (N_13261,N_11584,N_10501);
or U13262 (N_13262,N_11517,N_11816);
or U13263 (N_13263,N_10827,N_10951);
or U13264 (N_13264,N_10687,N_11497);
or U13265 (N_13265,N_10888,N_11044);
or U13266 (N_13266,N_11303,N_11194);
nor U13267 (N_13267,N_10962,N_10509);
nand U13268 (N_13268,N_11424,N_10501);
and U13269 (N_13269,N_11974,N_11523);
nor U13270 (N_13270,N_10980,N_11956);
nand U13271 (N_13271,N_10636,N_11107);
nor U13272 (N_13272,N_10840,N_11085);
nand U13273 (N_13273,N_11050,N_11053);
nand U13274 (N_13274,N_10700,N_10560);
nor U13275 (N_13275,N_10749,N_10887);
and U13276 (N_13276,N_11713,N_11357);
xnor U13277 (N_13277,N_11009,N_11427);
or U13278 (N_13278,N_11691,N_11488);
and U13279 (N_13279,N_11219,N_10862);
or U13280 (N_13280,N_10611,N_10504);
or U13281 (N_13281,N_11609,N_11407);
and U13282 (N_13282,N_11529,N_11501);
nor U13283 (N_13283,N_10834,N_11319);
or U13284 (N_13284,N_11856,N_11620);
or U13285 (N_13285,N_11681,N_11135);
nor U13286 (N_13286,N_11675,N_11873);
or U13287 (N_13287,N_10566,N_10701);
nor U13288 (N_13288,N_11818,N_10912);
nand U13289 (N_13289,N_11851,N_11993);
nor U13290 (N_13290,N_10920,N_10975);
nor U13291 (N_13291,N_10949,N_10540);
and U13292 (N_13292,N_11525,N_10524);
and U13293 (N_13293,N_10721,N_11156);
nand U13294 (N_13294,N_10722,N_11964);
nor U13295 (N_13295,N_11286,N_11015);
nor U13296 (N_13296,N_11894,N_10534);
or U13297 (N_13297,N_11892,N_11433);
nor U13298 (N_13298,N_11775,N_10617);
and U13299 (N_13299,N_11102,N_11161);
xor U13300 (N_13300,N_11587,N_11195);
xnor U13301 (N_13301,N_11370,N_10966);
or U13302 (N_13302,N_10815,N_10755);
and U13303 (N_13303,N_10794,N_10710);
nand U13304 (N_13304,N_10875,N_10905);
and U13305 (N_13305,N_11035,N_11257);
nand U13306 (N_13306,N_10752,N_11408);
nor U13307 (N_13307,N_11227,N_11340);
nand U13308 (N_13308,N_11014,N_11406);
nand U13309 (N_13309,N_11742,N_11839);
and U13310 (N_13310,N_11171,N_10658);
xnor U13311 (N_13311,N_10854,N_10975);
and U13312 (N_13312,N_11004,N_11142);
nand U13313 (N_13313,N_11391,N_10897);
or U13314 (N_13314,N_10995,N_11781);
or U13315 (N_13315,N_11014,N_11408);
xnor U13316 (N_13316,N_10586,N_11996);
or U13317 (N_13317,N_11572,N_11114);
nand U13318 (N_13318,N_11267,N_10594);
xnor U13319 (N_13319,N_10732,N_10612);
nor U13320 (N_13320,N_10705,N_11983);
or U13321 (N_13321,N_11031,N_10671);
and U13322 (N_13322,N_10775,N_11122);
nand U13323 (N_13323,N_11873,N_11222);
nor U13324 (N_13324,N_11594,N_11363);
nor U13325 (N_13325,N_11145,N_11227);
or U13326 (N_13326,N_10861,N_11473);
and U13327 (N_13327,N_10865,N_11176);
xor U13328 (N_13328,N_11736,N_10672);
nor U13329 (N_13329,N_11182,N_11045);
or U13330 (N_13330,N_11636,N_10701);
nor U13331 (N_13331,N_10818,N_11680);
nand U13332 (N_13332,N_10851,N_11620);
or U13333 (N_13333,N_11854,N_11432);
or U13334 (N_13334,N_10540,N_10775);
nand U13335 (N_13335,N_11308,N_11701);
nor U13336 (N_13336,N_10725,N_11450);
nor U13337 (N_13337,N_11172,N_10939);
or U13338 (N_13338,N_11474,N_10861);
and U13339 (N_13339,N_11987,N_11607);
and U13340 (N_13340,N_11415,N_11957);
xnor U13341 (N_13341,N_11973,N_10645);
or U13342 (N_13342,N_11362,N_11276);
nand U13343 (N_13343,N_11660,N_11212);
nand U13344 (N_13344,N_10750,N_11984);
or U13345 (N_13345,N_11475,N_10721);
or U13346 (N_13346,N_11358,N_11788);
or U13347 (N_13347,N_10761,N_10572);
xnor U13348 (N_13348,N_11911,N_11651);
nand U13349 (N_13349,N_10986,N_11427);
nand U13350 (N_13350,N_11556,N_10739);
nand U13351 (N_13351,N_10879,N_11481);
xor U13352 (N_13352,N_11848,N_10814);
and U13353 (N_13353,N_10744,N_10988);
xor U13354 (N_13354,N_11215,N_11515);
and U13355 (N_13355,N_11850,N_11533);
or U13356 (N_13356,N_11258,N_10747);
or U13357 (N_13357,N_10770,N_11703);
nor U13358 (N_13358,N_11171,N_11993);
nand U13359 (N_13359,N_10811,N_10733);
nand U13360 (N_13360,N_10563,N_10922);
nand U13361 (N_13361,N_11302,N_11250);
and U13362 (N_13362,N_10963,N_10912);
nor U13363 (N_13363,N_10742,N_11271);
xnor U13364 (N_13364,N_10660,N_11210);
nor U13365 (N_13365,N_11350,N_11642);
and U13366 (N_13366,N_10893,N_10614);
nor U13367 (N_13367,N_11504,N_10904);
nor U13368 (N_13368,N_11963,N_11364);
nor U13369 (N_13369,N_11170,N_11795);
xnor U13370 (N_13370,N_11330,N_11391);
or U13371 (N_13371,N_11035,N_11022);
nand U13372 (N_13372,N_10703,N_11486);
nand U13373 (N_13373,N_11148,N_11072);
nand U13374 (N_13374,N_10820,N_11923);
and U13375 (N_13375,N_11641,N_10784);
nor U13376 (N_13376,N_11777,N_11917);
or U13377 (N_13377,N_10512,N_11576);
nand U13378 (N_13378,N_11435,N_11137);
nor U13379 (N_13379,N_10546,N_11517);
or U13380 (N_13380,N_11802,N_11646);
nand U13381 (N_13381,N_10786,N_11244);
and U13382 (N_13382,N_10692,N_11880);
and U13383 (N_13383,N_11125,N_11886);
nand U13384 (N_13384,N_11443,N_10864);
and U13385 (N_13385,N_10753,N_11660);
and U13386 (N_13386,N_11030,N_10903);
nand U13387 (N_13387,N_11669,N_11693);
nor U13388 (N_13388,N_11915,N_11102);
or U13389 (N_13389,N_10739,N_11401);
nand U13390 (N_13390,N_11165,N_11538);
nor U13391 (N_13391,N_10714,N_10778);
and U13392 (N_13392,N_11966,N_11178);
nand U13393 (N_13393,N_11302,N_10958);
xor U13394 (N_13394,N_11718,N_11491);
or U13395 (N_13395,N_10779,N_11753);
or U13396 (N_13396,N_11090,N_10929);
and U13397 (N_13397,N_11489,N_10530);
xor U13398 (N_13398,N_10871,N_10967);
and U13399 (N_13399,N_11249,N_10540);
or U13400 (N_13400,N_10885,N_10578);
nor U13401 (N_13401,N_11243,N_10917);
and U13402 (N_13402,N_11575,N_10679);
nand U13403 (N_13403,N_11476,N_11916);
xnor U13404 (N_13404,N_10701,N_10532);
and U13405 (N_13405,N_11748,N_11896);
nor U13406 (N_13406,N_11457,N_11660);
and U13407 (N_13407,N_11458,N_10589);
xor U13408 (N_13408,N_11143,N_10531);
nand U13409 (N_13409,N_11690,N_11696);
and U13410 (N_13410,N_10715,N_11943);
nor U13411 (N_13411,N_11993,N_11862);
nand U13412 (N_13412,N_11396,N_11572);
nand U13413 (N_13413,N_10625,N_11848);
xor U13414 (N_13414,N_11126,N_11062);
and U13415 (N_13415,N_11480,N_11731);
nand U13416 (N_13416,N_11995,N_10721);
or U13417 (N_13417,N_10611,N_10699);
or U13418 (N_13418,N_11852,N_10836);
xnor U13419 (N_13419,N_11905,N_10650);
and U13420 (N_13420,N_11198,N_10921);
nand U13421 (N_13421,N_11427,N_10690);
nand U13422 (N_13422,N_11422,N_10591);
nor U13423 (N_13423,N_11377,N_11410);
and U13424 (N_13424,N_10887,N_10765);
or U13425 (N_13425,N_11746,N_11695);
nand U13426 (N_13426,N_11621,N_11488);
nand U13427 (N_13427,N_11907,N_10576);
or U13428 (N_13428,N_11911,N_11423);
xor U13429 (N_13429,N_10735,N_11825);
or U13430 (N_13430,N_11638,N_11556);
xor U13431 (N_13431,N_11813,N_11644);
or U13432 (N_13432,N_11138,N_11537);
or U13433 (N_13433,N_10971,N_10927);
xor U13434 (N_13434,N_11014,N_11115);
or U13435 (N_13435,N_11977,N_11013);
or U13436 (N_13436,N_11672,N_11595);
and U13437 (N_13437,N_10600,N_11906);
nor U13438 (N_13438,N_10809,N_11461);
and U13439 (N_13439,N_10551,N_10562);
nand U13440 (N_13440,N_11888,N_10956);
and U13441 (N_13441,N_11507,N_11650);
nor U13442 (N_13442,N_11481,N_10575);
nor U13443 (N_13443,N_11040,N_10649);
and U13444 (N_13444,N_10702,N_11604);
xor U13445 (N_13445,N_11167,N_10759);
and U13446 (N_13446,N_11054,N_11345);
or U13447 (N_13447,N_11288,N_11498);
or U13448 (N_13448,N_10720,N_11851);
nor U13449 (N_13449,N_11138,N_11494);
nor U13450 (N_13450,N_11572,N_10795);
xnor U13451 (N_13451,N_11516,N_11545);
and U13452 (N_13452,N_10877,N_10702);
or U13453 (N_13453,N_11804,N_10850);
nor U13454 (N_13454,N_10796,N_10838);
and U13455 (N_13455,N_11583,N_11767);
and U13456 (N_13456,N_10860,N_11065);
nand U13457 (N_13457,N_11893,N_11475);
and U13458 (N_13458,N_11134,N_11709);
or U13459 (N_13459,N_11174,N_11609);
and U13460 (N_13460,N_11032,N_11241);
nand U13461 (N_13461,N_11540,N_11892);
or U13462 (N_13462,N_10584,N_11954);
and U13463 (N_13463,N_10612,N_10718);
and U13464 (N_13464,N_10531,N_11553);
or U13465 (N_13465,N_11228,N_10945);
nand U13466 (N_13466,N_10556,N_11680);
or U13467 (N_13467,N_11173,N_11893);
nand U13468 (N_13468,N_11247,N_11010);
nand U13469 (N_13469,N_11015,N_10566);
nand U13470 (N_13470,N_11534,N_10579);
nand U13471 (N_13471,N_11614,N_11679);
or U13472 (N_13472,N_11146,N_11677);
nand U13473 (N_13473,N_11558,N_11653);
xor U13474 (N_13474,N_10743,N_10658);
or U13475 (N_13475,N_11846,N_11651);
nand U13476 (N_13476,N_11761,N_11008);
and U13477 (N_13477,N_11533,N_10826);
or U13478 (N_13478,N_11276,N_11116);
nor U13479 (N_13479,N_11674,N_11798);
and U13480 (N_13480,N_11568,N_11047);
or U13481 (N_13481,N_11703,N_10962);
nor U13482 (N_13482,N_11187,N_11163);
and U13483 (N_13483,N_11240,N_11328);
and U13484 (N_13484,N_10642,N_11344);
nor U13485 (N_13485,N_11924,N_11459);
and U13486 (N_13486,N_11109,N_11345);
xnor U13487 (N_13487,N_11239,N_11948);
nor U13488 (N_13488,N_10668,N_10638);
or U13489 (N_13489,N_11390,N_11161);
nand U13490 (N_13490,N_11772,N_11585);
or U13491 (N_13491,N_11986,N_11569);
and U13492 (N_13492,N_10997,N_10777);
nand U13493 (N_13493,N_10775,N_11788);
nor U13494 (N_13494,N_10743,N_10544);
nand U13495 (N_13495,N_11365,N_10664);
or U13496 (N_13496,N_11048,N_10645);
xnor U13497 (N_13497,N_11728,N_11768);
nor U13498 (N_13498,N_10836,N_11976);
or U13499 (N_13499,N_11443,N_11609);
nand U13500 (N_13500,N_12574,N_12632);
nand U13501 (N_13501,N_12091,N_13172);
and U13502 (N_13502,N_12039,N_12541);
xnor U13503 (N_13503,N_12411,N_12621);
xor U13504 (N_13504,N_12428,N_12085);
nor U13505 (N_13505,N_13055,N_12043);
nand U13506 (N_13506,N_12671,N_13129);
nor U13507 (N_13507,N_12740,N_12576);
xnor U13508 (N_13508,N_12603,N_12620);
and U13509 (N_13509,N_13216,N_13081);
or U13510 (N_13510,N_12993,N_12330);
or U13511 (N_13511,N_12992,N_13179);
nor U13512 (N_13512,N_12425,N_12097);
nand U13513 (N_13513,N_12797,N_12563);
nor U13514 (N_13514,N_13357,N_12329);
nand U13515 (N_13515,N_13446,N_13286);
nand U13516 (N_13516,N_12517,N_12301);
nor U13517 (N_13517,N_12659,N_13127);
and U13518 (N_13518,N_13436,N_12415);
or U13519 (N_13519,N_13365,N_13314);
and U13520 (N_13520,N_13227,N_12472);
or U13521 (N_13521,N_12610,N_12414);
nand U13522 (N_13522,N_12677,N_12887);
nor U13523 (N_13523,N_13236,N_12296);
nand U13524 (N_13524,N_12359,N_13095);
xnor U13525 (N_13525,N_13387,N_13437);
nor U13526 (N_13526,N_12124,N_12263);
or U13527 (N_13527,N_13067,N_12958);
xor U13528 (N_13528,N_12780,N_13298);
or U13529 (N_13529,N_12573,N_13377);
or U13530 (N_13530,N_13197,N_12736);
xnor U13531 (N_13531,N_12836,N_13145);
and U13532 (N_13532,N_13428,N_13186);
or U13533 (N_13533,N_12936,N_12783);
and U13534 (N_13534,N_12223,N_12073);
nor U13535 (N_13535,N_12109,N_12021);
nor U13536 (N_13536,N_12034,N_13287);
and U13537 (N_13537,N_12712,N_12844);
nor U13538 (N_13538,N_12834,N_13169);
nor U13539 (N_13539,N_12969,N_13176);
or U13540 (N_13540,N_12549,N_12130);
and U13541 (N_13541,N_13394,N_12737);
nor U13542 (N_13542,N_12633,N_12370);
nand U13543 (N_13543,N_13209,N_12930);
or U13544 (N_13544,N_13331,N_13320);
and U13545 (N_13545,N_12427,N_12278);
and U13546 (N_13546,N_12470,N_12644);
and U13547 (N_13547,N_12165,N_13049);
and U13548 (N_13548,N_12688,N_12842);
nand U13549 (N_13549,N_13430,N_12041);
nor U13550 (N_13550,N_12618,N_12848);
nand U13551 (N_13551,N_12657,N_12469);
and U13552 (N_13552,N_12817,N_13375);
nand U13553 (N_13553,N_13392,N_12260);
nand U13554 (N_13554,N_12285,N_12434);
nor U13555 (N_13555,N_12976,N_13107);
nand U13556 (N_13556,N_12920,N_13166);
or U13557 (N_13557,N_12599,N_12652);
or U13558 (N_13558,N_12042,N_13251);
nand U13559 (N_13559,N_12116,N_12353);
nor U13560 (N_13560,N_12303,N_12932);
or U13561 (N_13561,N_12024,N_12485);
xor U13562 (N_13562,N_12382,N_13143);
and U13563 (N_13563,N_12525,N_12261);
and U13564 (N_13564,N_13250,N_12514);
or U13565 (N_13565,N_12935,N_12372);
nor U13566 (N_13566,N_13241,N_12964);
nand U13567 (N_13567,N_12600,N_12283);
and U13568 (N_13568,N_12539,N_12536);
and U13569 (N_13569,N_13473,N_12735);
or U13570 (N_13570,N_12955,N_13259);
xnor U13571 (N_13571,N_12203,N_12271);
and U13572 (N_13572,N_13489,N_12210);
nand U13573 (N_13573,N_12134,N_12457);
and U13574 (N_13574,N_12018,N_13461);
nand U13575 (N_13575,N_12937,N_12369);
nand U13576 (N_13576,N_12860,N_12674);
nand U13577 (N_13577,N_12592,N_12533);
or U13578 (N_13578,N_12365,N_13496);
nor U13579 (N_13579,N_12154,N_12083);
nor U13580 (N_13580,N_13078,N_12529);
nand U13581 (N_13581,N_13327,N_13367);
or U13582 (N_13582,N_12702,N_12367);
and U13583 (N_13583,N_13344,N_13455);
and U13584 (N_13584,N_13256,N_12785);
xnor U13585 (N_13585,N_12497,N_12550);
nor U13586 (N_13586,N_12527,N_12123);
xnor U13587 (N_13587,N_12653,N_12241);
nor U13588 (N_13588,N_12647,N_12172);
nand U13589 (N_13589,N_13041,N_12381);
nor U13590 (N_13590,N_12136,N_12654);
nor U13591 (N_13591,N_12581,N_12884);
nor U13592 (N_13592,N_12145,N_12254);
nor U13593 (N_13593,N_13062,N_13244);
nand U13594 (N_13594,N_13371,N_13408);
and U13595 (N_13595,N_12128,N_13016);
nor U13596 (N_13596,N_13221,N_13118);
nor U13597 (N_13597,N_12507,N_13383);
nor U13598 (N_13598,N_12392,N_12997);
nand U13599 (N_13599,N_12755,N_12243);
or U13600 (N_13600,N_12886,N_13499);
nand U13601 (N_13601,N_12905,N_12888);
or U13602 (N_13602,N_13417,N_13283);
and U13603 (N_13603,N_12462,N_13029);
or U13604 (N_13604,N_12008,N_12929);
xnor U13605 (N_13605,N_12175,N_12733);
and U13606 (N_13606,N_12751,N_12690);
xor U13607 (N_13607,N_12163,N_12919);
nand U13608 (N_13608,N_13388,N_12569);
or U13609 (N_13609,N_12456,N_12294);
nand U13610 (N_13610,N_12629,N_13312);
nand U13611 (N_13611,N_12790,N_13152);
nor U13612 (N_13612,N_13103,N_12894);
nand U13613 (N_13613,N_12302,N_12126);
and U13614 (N_13614,N_12814,N_12962);
or U13615 (N_13615,N_13120,N_12227);
xor U13616 (N_13616,N_12917,N_12342);
or U13617 (N_13617,N_12501,N_13249);
or U13618 (N_13618,N_13155,N_13402);
and U13619 (N_13619,N_13463,N_12177);
nand U13620 (N_13620,N_13316,N_12351);
or U13621 (N_13621,N_12761,N_13201);
and U13622 (N_13622,N_12255,N_12849);
nand U13623 (N_13623,N_12200,N_12763);
nand U13624 (N_13624,N_12173,N_12720);
or U13625 (N_13625,N_12987,N_12216);
or U13626 (N_13626,N_12762,N_13454);
nand U13627 (N_13627,N_12194,N_13459);
and U13628 (N_13628,N_12412,N_12631);
nor U13629 (N_13629,N_12845,N_12960);
xor U13630 (N_13630,N_13262,N_12323);
and U13631 (N_13631,N_13258,N_13360);
and U13632 (N_13632,N_12511,N_12634);
nand U13633 (N_13633,N_13082,N_12304);
xnor U13634 (N_13634,N_13278,N_12193);
nor U13635 (N_13635,N_12312,N_13114);
nand U13636 (N_13636,N_12240,N_13228);
nor U13637 (N_13637,N_12284,N_12403);
nor U13638 (N_13638,N_13140,N_12057);
nand U13639 (N_13639,N_13247,N_12945);
nand U13640 (N_13640,N_13126,N_12608);
or U13641 (N_13641,N_12448,N_12521);
nand U13642 (N_13642,N_12524,N_13279);
or U13643 (N_13643,N_13415,N_12038);
nor U13644 (N_13644,N_12515,N_12277);
or U13645 (N_13645,N_12114,N_12874);
nand U13646 (N_13646,N_12025,N_12378);
or U13647 (N_13647,N_13181,N_13348);
or U13648 (N_13648,N_13215,N_13024);
nor U13649 (N_13649,N_12309,N_12584);
and U13650 (N_13650,N_12075,N_12858);
and U13651 (N_13651,N_13384,N_12899);
nand U13652 (N_13652,N_12396,N_12979);
nor U13653 (N_13653,N_12379,N_12878);
nor U13654 (N_13654,N_12204,N_12129);
nor U13655 (N_13655,N_12951,N_12292);
xnor U13656 (N_13656,N_12744,N_12575);
nor U13657 (N_13657,N_13273,N_13341);
and U13658 (N_13658,N_12120,N_13260);
or U13659 (N_13659,N_12387,N_13465);
nand U13660 (N_13660,N_13191,N_12221);
and U13661 (N_13661,N_12107,N_12914);
nand U13662 (N_13662,N_13486,N_12244);
nand U13663 (N_13663,N_13094,N_13013);
nor U13664 (N_13664,N_13476,N_12809);
xnor U13665 (N_13665,N_12236,N_12272);
nand U13666 (N_13666,N_12693,N_12326);
nand U13667 (N_13667,N_13347,N_12161);
or U13668 (N_13668,N_12670,N_13170);
and U13669 (N_13669,N_12832,N_13019);
and U13670 (N_13670,N_12101,N_13219);
nand U13671 (N_13671,N_13231,N_12746);
or U13672 (N_13672,N_13291,N_13440);
or U13673 (N_13673,N_12642,N_13196);
nand U13674 (N_13674,N_12486,N_12374);
xnor U13675 (N_13675,N_12625,N_12532);
and U13676 (N_13676,N_13009,N_12007);
nand U13677 (N_13677,N_13115,N_13335);
xor U13678 (N_13678,N_12417,N_12139);
or U13679 (N_13679,N_12125,N_12696);
or U13680 (N_13680,N_12667,N_12321);
nand U13681 (N_13681,N_12698,N_12155);
and U13682 (N_13682,N_13426,N_12703);
nor U13683 (N_13683,N_12835,N_12416);
and U13684 (N_13684,N_13400,N_13000);
xor U13685 (N_13685,N_12508,N_12896);
nand U13686 (N_13686,N_12251,N_13077);
or U13687 (N_13687,N_13192,N_12553);
and U13688 (N_13688,N_12289,N_13039);
nand U13689 (N_13689,N_12561,N_13222);
nand U13690 (N_13690,N_12559,N_12466);
nand U13691 (N_13691,N_12168,N_12582);
or U13692 (N_13692,N_12691,N_12646);
or U13693 (N_13693,N_13033,N_12557);
nor U13694 (N_13694,N_12178,N_12577);
and U13695 (N_13695,N_13492,N_12348);
or U13696 (N_13696,N_12731,N_12053);
xor U13697 (N_13697,N_12622,N_12767);
xor U13698 (N_13698,N_13272,N_12020);
and U13699 (N_13699,N_13178,N_13484);
or U13700 (N_13700,N_12764,N_13407);
nor U13701 (N_13701,N_12605,N_12186);
or U13702 (N_13702,N_12217,N_12407);
and U13703 (N_13703,N_12601,N_12266);
or U13704 (N_13704,N_12055,N_13467);
and U13705 (N_13705,N_12829,N_12921);
nand U13706 (N_13706,N_12355,N_13480);
and U13707 (N_13707,N_12482,N_12866);
nor U13708 (N_13708,N_12808,N_13482);
nor U13709 (N_13709,N_13306,N_12461);
or U13710 (N_13710,N_12555,N_12686);
nand U13711 (N_13711,N_13281,N_13004);
or U13712 (N_13712,N_12721,N_13157);
xnor U13713 (N_13713,N_12291,N_12117);
nand U13714 (N_13714,N_12941,N_12115);
or U13715 (N_13715,N_13416,N_13211);
nand U13716 (N_13716,N_12804,N_12389);
or U13717 (N_13717,N_13401,N_12707);
nor U13718 (N_13718,N_13253,N_13205);
nor U13719 (N_13719,N_12287,N_12395);
xor U13720 (N_13720,N_12910,N_12548);
or U13721 (N_13721,N_12813,N_13297);
nor U13722 (N_13722,N_12383,N_12138);
and U13723 (N_13723,N_12946,N_13443);
nor U13724 (N_13724,N_12617,N_13106);
nand U13725 (N_13725,N_12401,N_12830);
nor U13726 (N_13726,N_12071,N_13132);
nor U13727 (N_13727,N_13261,N_12509);
nor U13728 (N_13728,N_13254,N_13300);
xor U13729 (N_13729,N_12588,N_12554);
or U13730 (N_13730,N_13410,N_13310);
nor U13731 (N_13731,N_12870,N_12726);
and U13732 (N_13732,N_13154,N_12897);
nor U13733 (N_13733,N_12788,N_12841);
nand U13734 (N_13734,N_12350,N_12856);
nand U13735 (N_13735,N_12789,N_12019);
nand U13736 (N_13736,N_12597,N_12347);
and U13737 (N_13737,N_12257,N_12052);
or U13738 (N_13738,N_13425,N_12708);
or U13739 (N_13739,N_12170,N_12093);
xnor U13740 (N_13740,N_12441,N_12999);
and U13741 (N_13741,N_12049,N_12096);
xor U13742 (N_13742,N_12880,N_12787);
xor U13743 (N_13743,N_13223,N_12716);
or U13744 (N_13744,N_12158,N_12766);
and U13745 (N_13745,N_12637,N_12528);
nand U13746 (N_13746,N_13105,N_13042);
and U13747 (N_13747,N_13488,N_12916);
nand U13748 (N_13748,N_12220,N_12567);
nor U13749 (N_13749,N_13399,N_12754);
and U13750 (N_13750,N_12400,N_12794);
or U13751 (N_13751,N_13030,N_13137);
nand U13752 (N_13752,N_13195,N_13146);
or U13753 (N_13753,N_12824,N_13475);
and U13754 (N_13754,N_12076,N_12742);
nor U13755 (N_13755,N_13006,N_12939);
nand U13756 (N_13756,N_13074,N_12331);
nand U13757 (N_13757,N_12059,N_12628);
nor U13758 (N_13758,N_13429,N_12229);
xnor U13759 (N_13759,N_13269,N_12784);
nand U13760 (N_13760,N_13046,N_12424);
nor U13761 (N_13761,N_13060,N_12853);
or U13762 (N_13762,N_13063,N_13018);
and U13763 (N_13763,N_12885,N_12013);
nor U13764 (N_13764,N_12973,N_13175);
nor U13765 (N_13765,N_13217,N_12812);
and U13766 (N_13766,N_13449,N_12638);
or U13767 (N_13767,N_12118,N_13023);
and U13768 (N_13768,N_12922,N_12393);
nor U13769 (N_13769,N_13161,N_12782);
and U13770 (N_13770,N_13056,N_13128);
or U13771 (N_13771,N_13321,N_12732);
and U13772 (N_13772,N_12868,N_13433);
nor U13773 (N_13773,N_13020,N_13037);
and U13774 (N_13774,N_12171,N_13136);
nand U13775 (N_13775,N_13149,N_12942);
or U13776 (N_13776,N_13025,N_12966);
xor U13777 (N_13777,N_12239,N_12643);
or U13778 (N_13778,N_12974,N_12913);
nand U13779 (N_13779,N_12003,N_12336);
nor U13780 (N_13780,N_12094,N_13342);
and U13781 (N_13781,N_13343,N_12310);
nor U13782 (N_13782,N_12526,N_12893);
nor U13783 (N_13783,N_12440,N_13255);
xor U13784 (N_13784,N_12664,N_12743);
or U13785 (N_13785,N_12806,N_13150);
nand U13786 (N_13786,N_13069,N_12730);
nor U13787 (N_13787,N_12237,N_12859);
nand U13788 (N_13788,N_13317,N_12778);
nor U13789 (N_13789,N_13450,N_12196);
nand U13790 (N_13790,N_13393,N_13193);
nor U13791 (N_13791,N_12564,N_12104);
nor U13792 (N_13792,N_13379,N_12062);
nand U13793 (N_13793,N_12361,N_13307);
nor U13794 (N_13794,N_12458,N_12869);
and U13795 (N_13795,N_12169,N_13481);
nor U13796 (N_13796,N_12218,N_13374);
and U13797 (N_13797,N_13418,N_12673);
or U13798 (N_13798,N_13116,N_12623);
nand U13799 (N_13799,N_13057,N_12028);
and U13800 (N_13800,N_12591,N_13498);
xnor U13801 (N_13801,N_13304,N_13294);
xor U13802 (N_13802,N_12847,N_12965);
nor U13803 (N_13803,N_13160,N_12089);
or U13804 (N_13804,N_13366,N_13280);
nand U13805 (N_13805,N_12680,N_12727);
nor U13806 (N_13806,N_13288,N_12252);
nor U13807 (N_13807,N_12571,N_12040);
and U13808 (N_13808,N_12538,N_13212);
nor U13809 (N_13809,N_12818,N_12478);
nand U13810 (N_13810,N_13447,N_13035);
and U13811 (N_13811,N_12433,N_12197);
and U13812 (N_13812,N_12322,N_13048);
nor U13813 (N_13813,N_13293,N_12645);
nor U13814 (N_13814,N_13303,N_12516);
and U13815 (N_13815,N_13403,N_12102);
and U13816 (N_13816,N_12045,N_12611);
nor U13817 (N_13817,N_12319,N_12402);
nand U13818 (N_13818,N_12235,N_12700);
nor U13819 (N_13819,N_12820,N_12607);
nor U13820 (N_13820,N_12971,N_12248);
or U13821 (N_13821,N_12384,N_12500);
or U13822 (N_13822,N_12530,N_13071);
nand U13823 (N_13823,N_13124,N_13438);
or U13824 (N_13824,N_12443,N_12772);
and U13825 (N_13825,N_12810,N_13015);
nand U13826 (N_13826,N_12898,N_12014);
nand U13827 (N_13827,N_12706,N_12224);
and U13828 (N_13828,N_12775,N_12774);
nand U13829 (N_13829,N_12488,N_12816);
or U13830 (N_13830,N_13412,N_12222);
and U13831 (N_13831,N_12092,N_12662);
or U13832 (N_13832,N_12430,N_12495);
nor U13833 (N_13833,N_12906,N_13479);
and U13834 (N_13834,N_13117,N_12668);
or U13835 (N_13835,N_13066,N_12795);
nand U13836 (N_13836,N_13458,N_12182);
and U13837 (N_13837,N_13292,N_13245);
nand U13838 (N_13838,N_12314,N_12655);
xor U13839 (N_13839,N_13065,N_12658);
and U13840 (N_13840,N_12952,N_12146);
nor U13841 (N_13841,N_12811,N_13174);
and U13842 (N_13842,N_12035,N_12327);
nor U13843 (N_13843,N_12205,N_12349);
and U13844 (N_13844,N_12565,N_12069);
and U13845 (N_13845,N_13010,N_13100);
nor U13846 (N_13846,N_12245,N_12022);
nor U13847 (N_13847,N_12212,N_13084);
nor U13848 (N_13848,N_12988,N_13411);
nand U13849 (N_13849,N_12998,N_12475);
and U13850 (N_13850,N_13182,N_12892);
or U13851 (N_13851,N_12449,N_12980);
xnor U13852 (N_13852,N_13495,N_13336);
nand U13853 (N_13853,N_12846,N_12915);
or U13854 (N_13854,N_12149,N_12436);
nand U13855 (N_13855,N_12311,N_12724);
nor U13856 (N_13856,N_12699,N_12468);
or U13857 (N_13857,N_13134,N_12595);
xor U13858 (N_13858,N_12077,N_12641);
and U13859 (N_13859,N_12131,N_12981);
nand U13860 (N_13860,N_12972,N_12745);
nor U13861 (N_13861,N_13086,N_12523);
or U13862 (N_13862,N_12975,N_13239);
xnor U13863 (N_13863,N_12479,N_12079);
nor U13864 (N_13864,N_12288,N_13026);
nor U13865 (N_13865,N_13003,N_13434);
nand U13866 (N_13866,N_13096,N_12883);
or U13867 (N_13867,N_12465,N_12385);
xor U13868 (N_13868,N_12474,N_12406);
or U13869 (N_13869,N_12346,N_12450);
nor U13870 (N_13870,N_12070,N_12800);
nor U13871 (N_13871,N_12545,N_12048);
or U13872 (N_13872,N_12982,N_13271);
or U13873 (N_13873,N_12029,N_12873);
or U13874 (N_13874,N_12967,N_12044);
or U13875 (N_13875,N_12086,N_12923);
nand U13876 (N_13876,N_12332,N_12150);
or U13877 (N_13877,N_12851,N_12843);
or U13878 (N_13878,N_12300,N_12924);
or U13879 (N_13879,N_12211,N_12144);
or U13880 (N_13880,N_12318,N_13237);
xor U13881 (N_13881,N_12306,N_12748);
and U13882 (N_13882,N_13469,N_13319);
and U13883 (N_13883,N_12650,N_12802);
and U13884 (N_13884,N_12308,N_13268);
and U13885 (N_13885,N_12959,N_12606);
and U13886 (N_13886,N_12183,N_12159);
or U13887 (N_13887,N_12535,N_12000);
nand U13888 (N_13888,N_12589,N_13072);
and U13889 (N_13889,N_12678,N_12734);
and U13890 (N_13890,N_13102,N_12861);
nand U13891 (N_13891,N_13011,N_12598);
or U13892 (N_13892,N_13131,N_13194);
nor U13893 (N_13893,N_12017,N_12943);
nand U13894 (N_13894,N_12325,N_12487);
and U13895 (N_13895,N_12164,N_12391);
nand U13896 (N_13896,N_13439,N_13470);
or U13897 (N_13897,N_12704,N_13098);
or U13898 (N_13898,N_12586,N_12345);
or U13899 (N_13899,N_12410,N_13462);
or U13900 (N_13900,N_12438,N_12963);
or U13901 (N_13901,N_13159,N_13104);
xor U13902 (N_13902,N_12030,N_12320);
nor U13903 (N_13903,N_12174,N_13460);
or U13904 (N_13904,N_12911,N_13121);
nand U13905 (N_13905,N_13092,N_12009);
nor U13906 (N_13906,N_12047,N_13032);
nor U13907 (N_13907,N_12825,N_13008);
and U13908 (N_13908,N_13097,N_12881);
nor U13909 (N_13909,N_12119,N_13151);
nor U13910 (N_13910,N_12256,N_12750);
nor U13911 (N_13911,N_12463,N_12467);
and U13912 (N_13912,N_12759,N_12837);
nand U13913 (N_13913,N_13246,N_13266);
xnor U13914 (N_13914,N_12219,N_13276);
nand U13915 (N_13915,N_12953,N_12135);
and U13916 (N_13916,N_12950,N_12518);
nand U13917 (N_13917,N_12335,N_12640);
xor U13918 (N_13918,N_12356,N_13133);
or U13919 (N_13919,N_13180,N_13432);
and U13920 (N_13920,N_12232,N_12604);
nand U13921 (N_13921,N_13419,N_13075);
nand U13922 (N_13922,N_12088,N_12376);
nor U13923 (N_13923,N_12012,N_12828);
nand U13924 (N_13924,N_12895,N_12213);
nand U13925 (N_13925,N_13238,N_12684);
nor U13926 (N_13926,N_12099,N_13183);
nor U13927 (N_13927,N_12675,N_12713);
xnor U13928 (N_13928,N_12738,N_12033);
xnor U13929 (N_13929,N_13373,N_12275);
and U13930 (N_13930,N_13409,N_12187);
nor U13931 (N_13931,N_13378,N_13177);
nor U13932 (N_13932,N_12792,N_13210);
and U13933 (N_13933,N_12293,N_12421);
nor U13934 (N_13934,N_13189,N_12111);
nand U13935 (N_13935,N_13452,N_13220);
and U13936 (N_13936,N_13315,N_12143);
nor U13937 (N_13937,N_12334,N_12160);
xnor U13938 (N_13938,N_12050,N_13309);
or U13939 (N_13939,N_12231,N_12580);
or U13940 (N_13940,N_12253,N_12908);
nand U13941 (N_13941,N_12739,N_12333);
or U13942 (N_13942,N_13034,N_12409);
xnor U13943 (N_13943,N_12520,N_13352);
nand U13944 (N_13944,N_13285,N_12619);
nor U13945 (N_13945,N_13125,N_12585);
or U13946 (N_13946,N_12815,N_12770);
nand U13947 (N_13947,N_13349,N_13028);
nor U13948 (N_13948,N_12689,N_12961);
nand U13949 (N_13949,N_12281,N_13345);
and U13950 (N_13950,N_13040,N_12926);
nor U13951 (N_13951,N_12907,N_12872);
nand U13952 (N_13952,N_13295,N_12380);
xor U13953 (N_13953,N_13188,N_13017);
xnor U13954 (N_13954,N_13248,N_12016);
nor U13955 (N_13955,N_12429,N_13386);
or U13956 (N_13956,N_12725,N_12863);
and U13957 (N_13957,N_12666,N_12499);
and U13958 (N_13958,N_13204,N_12133);
or U13959 (N_13959,N_13144,N_13167);
and U13960 (N_13960,N_12390,N_13005);
nor U13961 (N_13961,N_13362,N_12397);
and U13962 (N_13962,N_13138,N_12026);
nor U13963 (N_13963,N_12343,N_12371);
and U13964 (N_13964,N_13141,N_13334);
or U13965 (N_13965,N_13089,N_13301);
or U13966 (N_13966,N_12840,N_12191);
nand U13967 (N_13967,N_13240,N_13083);
nor U13968 (N_13968,N_12799,N_12572);
and U13969 (N_13969,N_13308,N_12705);
and U13970 (N_13970,N_12460,N_12153);
and U13971 (N_13971,N_12781,N_12510);
or U13972 (N_13972,N_12862,N_13206);
or U13973 (N_13973,N_13045,N_13444);
xor U13974 (N_13974,N_13485,N_12912);
xor U13975 (N_13975,N_13275,N_13299);
or U13976 (N_13976,N_12295,N_12238);
nand U13977 (N_13977,N_12386,N_13477);
and U13978 (N_13978,N_12167,N_12566);
or U13979 (N_13979,N_12082,N_12206);
nor U13980 (N_13980,N_13333,N_12776);
nor U13981 (N_13981,N_12354,N_13421);
and U13982 (N_13982,N_13274,N_12192);
nor U13983 (N_13983,N_13311,N_12230);
xnor U13984 (N_13984,N_12519,N_12676);
and U13985 (N_13985,N_12270,N_13226);
and U13986 (N_13986,N_13364,N_12656);
and U13987 (N_13987,N_12865,N_12624);
and U13988 (N_13988,N_13381,N_13318);
nand U13989 (N_13989,N_12728,N_12749);
nor U13990 (N_13990,N_12627,N_12080);
and U13991 (N_13991,N_12105,N_12269);
nor U13992 (N_13992,N_12340,N_13346);
or U13993 (N_13993,N_12717,N_13202);
and U13994 (N_13994,N_12398,N_13478);
nand U13995 (N_13995,N_12771,N_13265);
and U13996 (N_13996,N_13340,N_12822);
or U13997 (N_13997,N_12362,N_12685);
and U13998 (N_13998,N_12188,N_12831);
and U13999 (N_13999,N_12968,N_13232);
and U14000 (N_14000,N_12977,N_12259);
and U14001 (N_14001,N_12454,N_12990);
or U14002 (N_14002,N_13058,N_12723);
nand U14003 (N_14003,N_12938,N_12803);
or U14004 (N_14004,N_12452,N_12328);
nand U14005 (N_14005,N_12084,N_13351);
or U14006 (N_14006,N_13323,N_12665);
or U14007 (N_14007,N_12758,N_13187);
nand U14008 (N_14008,N_13277,N_12209);
or U14009 (N_14009,N_12635,N_13064);
and U14010 (N_14010,N_12011,N_12768);
nor U14011 (N_14011,N_12337,N_12453);
nor U14012 (N_14012,N_13491,N_12991);
nor U14013 (N_14013,N_12364,N_12819);
and U14014 (N_14014,N_12857,N_12985);
nor U14015 (N_14015,N_13218,N_12298);
and U14016 (N_14016,N_12805,N_12630);
nor U14017 (N_14017,N_13332,N_13090);
or U14018 (N_14018,N_12729,N_12481);
and U14019 (N_14019,N_13445,N_12442);
nor U14020 (N_14020,N_12127,N_12001);
or U14021 (N_14021,N_12447,N_12064);
or U14022 (N_14022,N_13038,N_12201);
or U14023 (N_14023,N_13036,N_12722);
nor U14024 (N_14024,N_13184,N_12357);
nor U14025 (N_14025,N_13200,N_12989);
and U14026 (N_14026,N_12875,N_12451);
nand U14027 (N_14027,N_13313,N_13326);
nand U14028 (N_14028,N_12801,N_12491);
nor U14029 (N_14029,N_12697,N_13158);
nand U14030 (N_14030,N_12476,N_12512);
or U14031 (N_14031,N_13404,N_13397);
and U14032 (N_14032,N_12464,N_12274);
and U14033 (N_14033,N_12484,N_12185);
nand U14034 (N_14034,N_13267,N_12583);
nand U14035 (N_14035,N_12531,N_13153);
nor U14036 (N_14036,N_13471,N_13087);
nor U14037 (N_14037,N_13431,N_12940);
nor U14038 (N_14038,N_13472,N_12081);
and U14039 (N_14039,N_12002,N_13050);
nand U14040 (N_14040,N_12852,N_12546);
xnor U14041 (N_14041,N_12909,N_12683);
or U14042 (N_14042,N_13171,N_12681);
and U14043 (N_14043,N_12032,N_12552);
nor U14044 (N_14044,N_12338,N_12399);
or U14045 (N_14045,N_12826,N_12854);
and U14046 (N_14046,N_12694,N_12276);
xnor U14047 (N_14047,N_12791,N_12986);
or U14048 (N_14048,N_12877,N_12663);
xor U14049 (N_14049,N_12996,N_12543);
or U14050 (N_14050,N_12983,N_13199);
and U14051 (N_14051,N_12714,N_12423);
or U14052 (N_14052,N_12358,N_13466);
nor U14053 (N_14053,N_12228,N_12756);
and U14054 (N_14054,N_12375,N_13422);
and U14055 (N_14055,N_12777,N_12636);
and U14056 (N_14056,N_13079,N_12360);
and U14057 (N_14057,N_12394,N_13165);
and U14058 (N_14058,N_12570,N_12918);
or U14059 (N_14059,N_12268,N_12366);
nand U14060 (N_14060,N_12015,N_12498);
nor U14061 (N_14061,N_13494,N_12418);
and U14062 (N_14062,N_12547,N_13474);
and U14063 (N_14063,N_12956,N_13355);
or U14064 (N_14064,N_13405,N_13483);
or U14065 (N_14065,N_12198,N_13270);
and U14066 (N_14066,N_13361,N_13229);
nor U14067 (N_14067,N_12793,N_12151);
and U14068 (N_14068,N_12181,N_12184);
nor U14069 (N_14069,N_12513,N_13414);
nor U14070 (N_14070,N_13243,N_12054);
or U14071 (N_14071,N_13356,N_13091);
or U14072 (N_14072,N_13073,N_12544);
or U14073 (N_14073,N_12928,N_12307);
nand U14074 (N_14074,N_12065,N_13198);
or U14075 (N_14075,N_12503,N_12855);
nand U14076 (N_14076,N_13061,N_12010);
or U14077 (N_14077,N_12432,N_12578);
nand U14078 (N_14078,N_12058,N_12890);
or U14079 (N_14079,N_12542,N_12280);
xnor U14080 (N_14080,N_12821,N_12947);
nand U14081 (N_14081,N_13101,N_13339);
and U14082 (N_14082,N_12901,N_12879);
or U14083 (N_14083,N_12587,N_12265);
or U14084 (N_14084,N_13328,N_13370);
nand U14085 (N_14085,N_13368,N_12534);
and U14086 (N_14086,N_13139,N_12651);
nor U14087 (N_14087,N_12156,N_12970);
nor U14088 (N_14088,N_12027,N_12090);
and U14089 (N_14089,N_12954,N_12148);
nand U14090 (N_14090,N_13113,N_12339);
or U14091 (N_14091,N_12649,N_12108);
nand U14092 (N_14092,N_13148,N_13208);
nor U14093 (N_14093,N_13305,N_13001);
xnor U14094 (N_14094,N_12098,N_13085);
or U14095 (N_14095,N_13325,N_13289);
nand U14096 (N_14096,N_12141,N_12413);
nor U14097 (N_14097,N_13156,N_12214);
nand U14098 (N_14098,N_12695,N_13135);
nor U14099 (N_14099,N_13027,N_12445);
nor U14100 (N_14100,N_12046,N_13213);
xnor U14101 (N_14101,N_12494,N_13427);
nand U14102 (N_14102,N_12602,N_12103);
nor U14103 (N_14103,N_12246,N_13406);
or U14104 (N_14104,N_12121,N_12037);
or U14105 (N_14105,N_12437,N_12556);
or U14106 (N_14106,N_12426,N_12299);
and U14107 (N_14107,N_12142,N_12408);
and U14108 (N_14108,N_12439,N_12639);
nand U14109 (N_14109,N_13391,N_12247);
xor U14110 (N_14110,N_12373,N_12687);
xor U14111 (N_14111,N_13456,N_12839);
nor U14112 (N_14112,N_12612,N_12506);
xor U14113 (N_14113,N_13322,N_13119);
nor U14114 (N_14114,N_12850,N_13442);
nand U14115 (N_14115,N_12233,N_12036);
or U14116 (N_14116,N_13376,N_12051);
or U14117 (N_14117,N_13413,N_12579);
or U14118 (N_14118,N_13490,N_12900);
and U14119 (N_14119,N_12492,N_13441);
nand U14120 (N_14120,N_12226,N_13354);
or U14121 (N_14121,N_13163,N_13052);
nand U14122 (N_14122,N_12477,N_12444);
nand U14123 (N_14123,N_12422,N_12242);
xnor U14124 (N_14124,N_13257,N_12072);
xor U14125 (N_14125,N_12994,N_13168);
and U14126 (N_14126,N_12388,N_12368);
nor U14127 (N_14127,N_12823,N_13396);
or U14128 (N_14128,N_13225,N_12669);
and U14129 (N_14129,N_12189,N_12068);
or U14130 (N_14130,N_13337,N_12558);
or U14131 (N_14131,N_12827,N_12264);
and U14132 (N_14132,N_12005,N_12833);
nor U14133 (N_14133,N_12316,N_13264);
or U14134 (N_14134,N_12060,N_12066);
nand U14135 (N_14135,N_12202,N_12949);
and U14136 (N_14136,N_12313,N_12480);
nor U14137 (N_14137,N_13284,N_13021);
nand U14138 (N_14138,N_12435,N_12023);
or U14139 (N_14139,N_12207,N_12773);
xor U14140 (N_14140,N_13338,N_12902);
nand U14141 (N_14141,N_13324,N_12190);
or U14142 (N_14142,N_12147,N_13088);
nor U14143 (N_14143,N_13173,N_12157);
nand U14144 (N_14144,N_13302,N_12769);
nand U14145 (N_14145,N_12838,N_12615);
and U14146 (N_14146,N_12927,N_13350);
and U14147 (N_14147,N_12590,N_13385);
nor U14148 (N_14148,N_13031,N_12709);
xor U14149 (N_14149,N_13420,N_12286);
and U14150 (N_14150,N_13012,N_12341);
or U14151 (N_14151,N_12290,N_13380);
nor U14152 (N_14152,N_12661,N_13207);
nand U14153 (N_14153,N_12798,N_13099);
or U14154 (N_14154,N_12106,N_12882);
nand U14155 (N_14155,N_12137,N_12765);
nor U14156 (N_14156,N_12648,N_12344);
nor U14157 (N_14157,N_12262,N_12864);
and U14158 (N_14158,N_13059,N_13224);
nor U14159 (N_14159,N_12305,N_13359);
or U14160 (N_14160,N_13329,N_12891);
nand U14161 (N_14161,N_12063,N_12672);
or U14162 (N_14162,N_12679,N_12199);
xnor U14163 (N_14163,N_13464,N_13109);
or U14164 (N_14164,N_12682,N_12490);
and U14165 (N_14165,N_12903,N_12719);
nor U14166 (N_14166,N_13468,N_12540);
nor U14167 (N_14167,N_12493,N_13369);
nand U14168 (N_14168,N_12455,N_12944);
and U14169 (N_14169,N_13235,N_12250);
nand U14170 (N_14170,N_12537,N_12660);
and U14171 (N_14171,N_12074,N_13185);
nor U14172 (N_14172,N_12234,N_12249);
nand U14173 (N_14173,N_13363,N_13123);
nor U14174 (N_14174,N_12752,N_12282);
and U14175 (N_14175,N_12225,N_12419);
and U14176 (N_14176,N_13203,N_12715);
nand U14177 (N_14177,N_12934,N_12180);
or U14178 (N_14178,N_13448,N_12176);
nor U14179 (N_14179,N_13070,N_12166);
nor U14180 (N_14180,N_13353,N_12522);
or U14181 (N_14181,N_12004,N_12113);
nand U14182 (N_14182,N_13130,N_12995);
and U14183 (N_14183,N_12087,N_12504);
nand U14184 (N_14184,N_12273,N_13054);
and U14185 (N_14185,N_12446,N_12140);
xor U14186 (N_14186,N_12110,N_13389);
and U14187 (N_14187,N_12747,N_12377);
and U14188 (N_14188,N_13053,N_12267);
and U14189 (N_14189,N_12195,N_12984);
xor U14190 (N_14190,N_12258,N_12718);
or U14191 (N_14191,N_13122,N_12867);
and U14192 (N_14192,N_12710,N_13330);
and U14193 (N_14193,N_13395,N_13043);
or U14194 (N_14194,N_12179,N_13457);
nor U14195 (N_14195,N_12122,N_12100);
or U14196 (N_14196,N_12889,N_12701);
or U14197 (N_14197,N_13358,N_13162);
nand U14198 (N_14198,N_13047,N_12796);
or U14199 (N_14199,N_12473,N_12505);
nor U14200 (N_14200,N_12904,N_13390);
and U14201 (N_14201,N_13487,N_12324);
nand U14202 (N_14202,N_13382,N_12056);
or U14203 (N_14203,N_12562,N_13076);
and U14204 (N_14204,N_12162,N_12948);
and U14205 (N_14205,N_12626,N_13242);
or U14206 (N_14206,N_12483,N_12095);
nor U14207 (N_14207,N_12420,N_13451);
and U14208 (N_14208,N_12760,N_13423);
and U14209 (N_14209,N_12978,N_12779);
nor U14210 (N_14210,N_12741,N_13110);
and U14211 (N_14211,N_12933,N_12613);
nand U14212 (N_14212,N_12405,N_12757);
nor U14213 (N_14213,N_13080,N_13398);
and U14214 (N_14214,N_12317,N_12297);
nor U14215 (N_14215,N_12594,N_13230);
and U14216 (N_14216,N_12067,N_12496);
nor U14217 (N_14217,N_12786,N_13164);
xnor U14218 (N_14218,N_13252,N_12404);
nand U14219 (N_14219,N_12471,N_13044);
and U14220 (N_14220,N_12596,N_13453);
nand U14221 (N_14221,N_12459,N_13002);
nand U14222 (N_14222,N_13290,N_13282);
nand U14223 (N_14223,N_12711,N_12279);
nor U14224 (N_14224,N_12502,N_12957);
nand U14225 (N_14225,N_12614,N_12551);
xnor U14226 (N_14226,N_12006,N_13435);
and U14227 (N_14227,N_12352,N_12609);
or U14228 (N_14228,N_12215,N_13022);
nor U14229 (N_14229,N_12031,N_13296);
nor U14230 (N_14230,N_12132,N_13372);
or U14231 (N_14231,N_12807,N_12593);
nand U14232 (N_14232,N_12753,N_13147);
or U14233 (N_14233,N_13112,N_12112);
and U14234 (N_14234,N_13007,N_12431);
xor U14235 (N_14235,N_12871,N_12152);
and U14236 (N_14236,N_12925,N_13068);
or U14237 (N_14237,N_13263,N_13111);
and U14238 (N_14238,N_13214,N_13424);
or U14239 (N_14239,N_12315,N_12363);
or U14240 (N_14240,N_12931,N_12078);
nor U14241 (N_14241,N_13497,N_13051);
nor U14242 (N_14242,N_12876,N_13093);
nand U14243 (N_14243,N_12208,N_13190);
and U14244 (N_14244,N_13233,N_12568);
nand U14245 (N_14245,N_12616,N_12489);
and U14246 (N_14246,N_12560,N_13234);
or U14247 (N_14247,N_13014,N_12061);
nor U14248 (N_14248,N_13493,N_13108);
xnor U14249 (N_14249,N_13142,N_12692);
or U14250 (N_14250,N_13199,N_12835);
nand U14251 (N_14251,N_12999,N_13307);
xnor U14252 (N_14252,N_12926,N_13085);
or U14253 (N_14253,N_12729,N_12311);
nand U14254 (N_14254,N_12895,N_13032);
or U14255 (N_14255,N_12479,N_13487);
xnor U14256 (N_14256,N_12956,N_12791);
or U14257 (N_14257,N_13236,N_12922);
nand U14258 (N_14258,N_12004,N_12578);
nor U14259 (N_14259,N_12480,N_12061);
nor U14260 (N_14260,N_12877,N_12517);
nand U14261 (N_14261,N_12881,N_13309);
or U14262 (N_14262,N_13370,N_13099);
nor U14263 (N_14263,N_13340,N_13060);
or U14264 (N_14264,N_12856,N_13472);
nand U14265 (N_14265,N_12384,N_12228);
nand U14266 (N_14266,N_12484,N_12610);
or U14267 (N_14267,N_13409,N_12819);
nor U14268 (N_14268,N_13075,N_12132);
nor U14269 (N_14269,N_12078,N_12928);
and U14270 (N_14270,N_13196,N_12760);
nand U14271 (N_14271,N_13006,N_12620);
or U14272 (N_14272,N_12315,N_13402);
xor U14273 (N_14273,N_12787,N_13149);
xnor U14274 (N_14274,N_12195,N_12877);
or U14275 (N_14275,N_12651,N_12078);
and U14276 (N_14276,N_12279,N_13350);
and U14277 (N_14277,N_12561,N_12887);
xnor U14278 (N_14278,N_12666,N_12573);
nand U14279 (N_14279,N_12072,N_13148);
and U14280 (N_14280,N_13181,N_12177);
nand U14281 (N_14281,N_12081,N_12817);
nand U14282 (N_14282,N_12600,N_12094);
and U14283 (N_14283,N_12050,N_13490);
or U14284 (N_14284,N_12811,N_12287);
nand U14285 (N_14285,N_13113,N_13267);
and U14286 (N_14286,N_12213,N_12835);
or U14287 (N_14287,N_12281,N_12762);
nand U14288 (N_14288,N_13294,N_13295);
and U14289 (N_14289,N_12647,N_12512);
and U14290 (N_14290,N_13098,N_12389);
nand U14291 (N_14291,N_12514,N_12923);
or U14292 (N_14292,N_13008,N_12866);
and U14293 (N_14293,N_12146,N_13038);
and U14294 (N_14294,N_13257,N_12595);
or U14295 (N_14295,N_12846,N_12408);
nand U14296 (N_14296,N_12771,N_12674);
nand U14297 (N_14297,N_13441,N_12331);
nor U14298 (N_14298,N_12753,N_12033);
nand U14299 (N_14299,N_12559,N_13308);
or U14300 (N_14300,N_12103,N_12878);
and U14301 (N_14301,N_12498,N_13279);
or U14302 (N_14302,N_12305,N_13024);
nand U14303 (N_14303,N_12185,N_13273);
nor U14304 (N_14304,N_12289,N_12895);
nand U14305 (N_14305,N_13142,N_13003);
and U14306 (N_14306,N_13134,N_12204);
nor U14307 (N_14307,N_13067,N_12521);
xnor U14308 (N_14308,N_12805,N_12167);
or U14309 (N_14309,N_12412,N_13087);
nor U14310 (N_14310,N_12110,N_12896);
nor U14311 (N_14311,N_12304,N_12895);
nor U14312 (N_14312,N_12302,N_12735);
nor U14313 (N_14313,N_13411,N_12982);
and U14314 (N_14314,N_12105,N_12628);
or U14315 (N_14315,N_12994,N_13259);
nor U14316 (N_14316,N_12214,N_12863);
or U14317 (N_14317,N_12823,N_12371);
nor U14318 (N_14318,N_12318,N_12143);
and U14319 (N_14319,N_12246,N_13423);
or U14320 (N_14320,N_13449,N_12128);
nor U14321 (N_14321,N_12006,N_12913);
nor U14322 (N_14322,N_12668,N_12685);
or U14323 (N_14323,N_12204,N_12390);
nand U14324 (N_14324,N_12019,N_12752);
or U14325 (N_14325,N_12171,N_12740);
nand U14326 (N_14326,N_12732,N_12611);
nor U14327 (N_14327,N_12382,N_12325);
and U14328 (N_14328,N_12268,N_13261);
nor U14329 (N_14329,N_12365,N_12915);
nand U14330 (N_14330,N_13425,N_12760);
and U14331 (N_14331,N_12007,N_12255);
nand U14332 (N_14332,N_12889,N_12859);
and U14333 (N_14333,N_12622,N_13228);
nor U14334 (N_14334,N_12517,N_12530);
and U14335 (N_14335,N_12289,N_13479);
or U14336 (N_14336,N_13060,N_12692);
and U14337 (N_14337,N_12980,N_13496);
nand U14338 (N_14338,N_12936,N_12398);
nor U14339 (N_14339,N_13047,N_13479);
nand U14340 (N_14340,N_13330,N_12740);
or U14341 (N_14341,N_12006,N_13194);
nand U14342 (N_14342,N_12757,N_13339);
nor U14343 (N_14343,N_12921,N_12996);
nand U14344 (N_14344,N_12239,N_13414);
or U14345 (N_14345,N_12113,N_12336);
nor U14346 (N_14346,N_12190,N_12966);
or U14347 (N_14347,N_13268,N_13042);
or U14348 (N_14348,N_12666,N_12143);
nand U14349 (N_14349,N_13335,N_12625);
or U14350 (N_14350,N_13283,N_12162);
or U14351 (N_14351,N_12011,N_13029);
or U14352 (N_14352,N_13129,N_12966);
nand U14353 (N_14353,N_13143,N_12623);
nor U14354 (N_14354,N_13066,N_12977);
or U14355 (N_14355,N_13086,N_13334);
nor U14356 (N_14356,N_12739,N_13036);
or U14357 (N_14357,N_12003,N_12975);
nor U14358 (N_14358,N_12900,N_13116);
nor U14359 (N_14359,N_12864,N_13443);
or U14360 (N_14360,N_12253,N_13148);
and U14361 (N_14361,N_12693,N_12178);
nand U14362 (N_14362,N_12708,N_12705);
or U14363 (N_14363,N_13496,N_12022);
and U14364 (N_14364,N_12711,N_13133);
nor U14365 (N_14365,N_13028,N_13232);
nand U14366 (N_14366,N_12351,N_13318);
or U14367 (N_14367,N_13251,N_13466);
and U14368 (N_14368,N_12772,N_12795);
nand U14369 (N_14369,N_12484,N_12467);
or U14370 (N_14370,N_13168,N_13098);
nand U14371 (N_14371,N_12781,N_13221);
xor U14372 (N_14372,N_13435,N_13192);
nand U14373 (N_14373,N_12746,N_13484);
and U14374 (N_14374,N_12289,N_12243);
or U14375 (N_14375,N_12373,N_12089);
and U14376 (N_14376,N_12153,N_13408);
nand U14377 (N_14377,N_12622,N_12983);
and U14378 (N_14378,N_12240,N_12774);
and U14379 (N_14379,N_13344,N_13272);
nand U14380 (N_14380,N_12123,N_13105);
or U14381 (N_14381,N_13245,N_12267);
and U14382 (N_14382,N_13415,N_12050);
nand U14383 (N_14383,N_13353,N_12453);
nand U14384 (N_14384,N_13491,N_12057);
nor U14385 (N_14385,N_13001,N_12753);
and U14386 (N_14386,N_12268,N_12091);
nor U14387 (N_14387,N_12804,N_12973);
nor U14388 (N_14388,N_12551,N_13357);
and U14389 (N_14389,N_12411,N_13016);
nand U14390 (N_14390,N_13448,N_13131);
and U14391 (N_14391,N_12824,N_12254);
xor U14392 (N_14392,N_12136,N_12338);
nor U14393 (N_14393,N_12330,N_13353);
or U14394 (N_14394,N_12666,N_12575);
or U14395 (N_14395,N_12340,N_13261);
nor U14396 (N_14396,N_12181,N_12863);
nor U14397 (N_14397,N_13138,N_12038);
or U14398 (N_14398,N_12698,N_12879);
and U14399 (N_14399,N_12043,N_12983);
nor U14400 (N_14400,N_12192,N_13112);
nand U14401 (N_14401,N_12030,N_12445);
and U14402 (N_14402,N_13111,N_12813);
and U14403 (N_14403,N_12419,N_12281);
nand U14404 (N_14404,N_12663,N_12713);
nor U14405 (N_14405,N_12070,N_13011);
or U14406 (N_14406,N_13395,N_12999);
or U14407 (N_14407,N_12986,N_12053);
nor U14408 (N_14408,N_12609,N_13009);
or U14409 (N_14409,N_12023,N_12474);
xor U14410 (N_14410,N_13255,N_12550);
nor U14411 (N_14411,N_12964,N_12751);
and U14412 (N_14412,N_13414,N_12133);
nand U14413 (N_14413,N_13042,N_13390);
or U14414 (N_14414,N_13028,N_13024);
nor U14415 (N_14415,N_13106,N_12206);
nand U14416 (N_14416,N_12080,N_13310);
nor U14417 (N_14417,N_12322,N_13034);
xor U14418 (N_14418,N_12520,N_13347);
nand U14419 (N_14419,N_12591,N_13182);
and U14420 (N_14420,N_13174,N_12925);
and U14421 (N_14421,N_12463,N_12308);
and U14422 (N_14422,N_12763,N_13154);
nand U14423 (N_14423,N_12657,N_13169);
or U14424 (N_14424,N_13010,N_13353);
and U14425 (N_14425,N_12581,N_12260);
and U14426 (N_14426,N_12222,N_13384);
nand U14427 (N_14427,N_13484,N_12072);
or U14428 (N_14428,N_12177,N_13464);
and U14429 (N_14429,N_12264,N_13220);
nand U14430 (N_14430,N_12010,N_12070);
or U14431 (N_14431,N_12429,N_12090);
nand U14432 (N_14432,N_12259,N_13462);
nand U14433 (N_14433,N_12319,N_13446);
and U14434 (N_14434,N_12444,N_13150);
nand U14435 (N_14435,N_13014,N_13098);
nor U14436 (N_14436,N_13257,N_12866);
and U14437 (N_14437,N_12786,N_12513);
or U14438 (N_14438,N_12583,N_12790);
nor U14439 (N_14439,N_12423,N_12086);
nand U14440 (N_14440,N_12199,N_12650);
xnor U14441 (N_14441,N_12751,N_12162);
or U14442 (N_14442,N_12805,N_13267);
nor U14443 (N_14443,N_12680,N_12122);
or U14444 (N_14444,N_12192,N_12134);
nand U14445 (N_14445,N_13423,N_13376);
nand U14446 (N_14446,N_13203,N_12894);
xnor U14447 (N_14447,N_13409,N_13444);
nand U14448 (N_14448,N_13386,N_13235);
nor U14449 (N_14449,N_12354,N_12909);
and U14450 (N_14450,N_13058,N_12514);
nor U14451 (N_14451,N_12308,N_13460);
nor U14452 (N_14452,N_12461,N_13296);
or U14453 (N_14453,N_13454,N_12718);
xor U14454 (N_14454,N_13267,N_12942);
nand U14455 (N_14455,N_13209,N_12521);
nand U14456 (N_14456,N_13334,N_12881);
and U14457 (N_14457,N_13177,N_13417);
or U14458 (N_14458,N_12671,N_12052);
nor U14459 (N_14459,N_13343,N_13221);
and U14460 (N_14460,N_12276,N_12894);
nor U14461 (N_14461,N_12497,N_12678);
or U14462 (N_14462,N_13341,N_12908);
xnor U14463 (N_14463,N_12783,N_12903);
and U14464 (N_14464,N_12786,N_12369);
or U14465 (N_14465,N_12992,N_12994);
and U14466 (N_14466,N_12826,N_13473);
xnor U14467 (N_14467,N_12797,N_13036);
nor U14468 (N_14468,N_12296,N_12601);
and U14469 (N_14469,N_13312,N_13073);
nor U14470 (N_14470,N_13351,N_12962);
nand U14471 (N_14471,N_13465,N_13385);
nand U14472 (N_14472,N_12048,N_12611);
or U14473 (N_14473,N_12296,N_12779);
nand U14474 (N_14474,N_12543,N_13245);
xor U14475 (N_14475,N_13148,N_12365);
nand U14476 (N_14476,N_12658,N_13346);
nand U14477 (N_14477,N_12438,N_13102);
and U14478 (N_14478,N_12009,N_12088);
or U14479 (N_14479,N_12293,N_13426);
nand U14480 (N_14480,N_13216,N_12814);
and U14481 (N_14481,N_12705,N_12224);
nand U14482 (N_14482,N_13081,N_12998);
or U14483 (N_14483,N_12090,N_13485);
nor U14484 (N_14484,N_13076,N_12444);
nor U14485 (N_14485,N_12634,N_12400);
nor U14486 (N_14486,N_12832,N_13290);
and U14487 (N_14487,N_12388,N_13330);
and U14488 (N_14488,N_13466,N_12377);
or U14489 (N_14489,N_12949,N_12180);
or U14490 (N_14490,N_12214,N_12539);
and U14491 (N_14491,N_13098,N_12358);
or U14492 (N_14492,N_12729,N_12157);
nor U14493 (N_14493,N_12589,N_12502);
or U14494 (N_14494,N_13265,N_12575);
nand U14495 (N_14495,N_12851,N_12786);
nand U14496 (N_14496,N_12983,N_12982);
nand U14497 (N_14497,N_13122,N_12329);
and U14498 (N_14498,N_12654,N_13298);
and U14499 (N_14499,N_13031,N_13446);
nor U14500 (N_14500,N_12049,N_12346);
and U14501 (N_14501,N_13171,N_12745);
or U14502 (N_14502,N_12641,N_13330);
nand U14503 (N_14503,N_12677,N_12102);
or U14504 (N_14504,N_13101,N_12976);
nand U14505 (N_14505,N_12878,N_12058);
or U14506 (N_14506,N_12707,N_12081);
and U14507 (N_14507,N_12134,N_12003);
nand U14508 (N_14508,N_13497,N_12101);
nor U14509 (N_14509,N_13484,N_12790);
and U14510 (N_14510,N_13343,N_12525);
nor U14511 (N_14511,N_12206,N_13267);
or U14512 (N_14512,N_12014,N_13186);
and U14513 (N_14513,N_13248,N_13277);
and U14514 (N_14514,N_13406,N_13465);
or U14515 (N_14515,N_12285,N_12342);
xnor U14516 (N_14516,N_13352,N_13299);
or U14517 (N_14517,N_12112,N_12566);
nor U14518 (N_14518,N_12810,N_12774);
nand U14519 (N_14519,N_12654,N_12371);
nor U14520 (N_14520,N_13079,N_12390);
and U14521 (N_14521,N_12413,N_12936);
and U14522 (N_14522,N_13431,N_13133);
nor U14523 (N_14523,N_12514,N_12703);
nand U14524 (N_14524,N_12621,N_13232);
and U14525 (N_14525,N_12240,N_12451);
or U14526 (N_14526,N_13207,N_12627);
and U14527 (N_14527,N_13270,N_12946);
or U14528 (N_14528,N_12287,N_12636);
nand U14529 (N_14529,N_12190,N_12430);
nor U14530 (N_14530,N_12154,N_13127);
nand U14531 (N_14531,N_13120,N_12986);
or U14532 (N_14532,N_12544,N_12228);
nand U14533 (N_14533,N_12339,N_12164);
nand U14534 (N_14534,N_12139,N_12359);
or U14535 (N_14535,N_12480,N_13179);
and U14536 (N_14536,N_12085,N_12163);
and U14537 (N_14537,N_12846,N_12590);
or U14538 (N_14538,N_13421,N_13468);
nand U14539 (N_14539,N_13122,N_13418);
and U14540 (N_14540,N_13437,N_12824);
nand U14541 (N_14541,N_12007,N_13249);
or U14542 (N_14542,N_13044,N_12054);
nor U14543 (N_14543,N_13054,N_12734);
and U14544 (N_14544,N_13424,N_12444);
nand U14545 (N_14545,N_13365,N_13138);
nand U14546 (N_14546,N_12969,N_12093);
xor U14547 (N_14547,N_12560,N_13332);
nand U14548 (N_14548,N_12087,N_12197);
and U14549 (N_14549,N_13226,N_12795);
and U14550 (N_14550,N_12545,N_13191);
nor U14551 (N_14551,N_12700,N_13112);
nor U14552 (N_14552,N_12250,N_13276);
nor U14553 (N_14553,N_13409,N_13125);
nor U14554 (N_14554,N_13149,N_12850);
and U14555 (N_14555,N_12984,N_12688);
and U14556 (N_14556,N_12377,N_12461);
and U14557 (N_14557,N_12219,N_12734);
nor U14558 (N_14558,N_13211,N_12353);
and U14559 (N_14559,N_13400,N_12110);
nand U14560 (N_14560,N_13256,N_12857);
xor U14561 (N_14561,N_12597,N_12315);
nand U14562 (N_14562,N_12478,N_13451);
or U14563 (N_14563,N_12214,N_12840);
nor U14564 (N_14564,N_13066,N_12918);
nand U14565 (N_14565,N_12922,N_13385);
nor U14566 (N_14566,N_13187,N_12781);
or U14567 (N_14567,N_12647,N_12283);
and U14568 (N_14568,N_12219,N_12201);
and U14569 (N_14569,N_13412,N_12670);
nand U14570 (N_14570,N_13335,N_13263);
nor U14571 (N_14571,N_12065,N_12435);
or U14572 (N_14572,N_13275,N_12307);
xor U14573 (N_14573,N_12833,N_13389);
or U14574 (N_14574,N_12154,N_13439);
nor U14575 (N_14575,N_12408,N_13153);
and U14576 (N_14576,N_12254,N_12208);
nor U14577 (N_14577,N_13087,N_12766);
nor U14578 (N_14578,N_12869,N_13189);
nand U14579 (N_14579,N_12131,N_12314);
nand U14580 (N_14580,N_13383,N_12779);
nand U14581 (N_14581,N_12805,N_13046);
nor U14582 (N_14582,N_12300,N_12563);
nand U14583 (N_14583,N_13296,N_12972);
and U14584 (N_14584,N_13466,N_12015);
xnor U14585 (N_14585,N_13306,N_12632);
or U14586 (N_14586,N_12172,N_12970);
xor U14587 (N_14587,N_12908,N_13437);
or U14588 (N_14588,N_13454,N_12964);
nand U14589 (N_14589,N_12148,N_12089);
and U14590 (N_14590,N_12027,N_12466);
nand U14591 (N_14591,N_12521,N_12733);
or U14592 (N_14592,N_12127,N_12600);
or U14593 (N_14593,N_12480,N_12114);
or U14594 (N_14594,N_12188,N_12384);
and U14595 (N_14595,N_12413,N_12103);
and U14596 (N_14596,N_13329,N_13025);
and U14597 (N_14597,N_12132,N_13345);
nor U14598 (N_14598,N_12444,N_12745);
or U14599 (N_14599,N_12271,N_12733);
or U14600 (N_14600,N_12642,N_12879);
nor U14601 (N_14601,N_12937,N_13399);
nand U14602 (N_14602,N_13388,N_13450);
nand U14603 (N_14603,N_13244,N_12838);
nand U14604 (N_14604,N_12883,N_12202);
or U14605 (N_14605,N_12638,N_12083);
nand U14606 (N_14606,N_12530,N_13157);
nand U14607 (N_14607,N_12552,N_12807);
and U14608 (N_14608,N_12741,N_12268);
or U14609 (N_14609,N_12076,N_12373);
nor U14610 (N_14610,N_12543,N_12170);
nor U14611 (N_14611,N_12035,N_12107);
nand U14612 (N_14612,N_12566,N_12341);
or U14613 (N_14613,N_12490,N_12684);
or U14614 (N_14614,N_12200,N_13161);
xor U14615 (N_14615,N_12238,N_12155);
and U14616 (N_14616,N_13265,N_13104);
nand U14617 (N_14617,N_12463,N_12281);
or U14618 (N_14618,N_12276,N_13104);
or U14619 (N_14619,N_12764,N_12016);
or U14620 (N_14620,N_12455,N_12755);
and U14621 (N_14621,N_12869,N_12884);
nand U14622 (N_14622,N_12691,N_12192);
or U14623 (N_14623,N_12898,N_12178);
xnor U14624 (N_14624,N_13171,N_13347);
or U14625 (N_14625,N_12661,N_13072);
and U14626 (N_14626,N_13289,N_12555);
or U14627 (N_14627,N_12006,N_12516);
or U14628 (N_14628,N_12603,N_13158);
and U14629 (N_14629,N_13395,N_12095);
and U14630 (N_14630,N_13080,N_12453);
and U14631 (N_14631,N_12989,N_12728);
or U14632 (N_14632,N_12851,N_12740);
nand U14633 (N_14633,N_12027,N_13086);
nand U14634 (N_14634,N_12947,N_13259);
nor U14635 (N_14635,N_13389,N_12715);
or U14636 (N_14636,N_13135,N_12320);
and U14637 (N_14637,N_12987,N_13150);
or U14638 (N_14638,N_12523,N_13227);
or U14639 (N_14639,N_12695,N_12921);
and U14640 (N_14640,N_13468,N_12925);
nand U14641 (N_14641,N_12222,N_13382);
nor U14642 (N_14642,N_13355,N_12709);
nor U14643 (N_14643,N_13475,N_12943);
nand U14644 (N_14644,N_13360,N_12824);
xnor U14645 (N_14645,N_12510,N_12359);
or U14646 (N_14646,N_12654,N_12513);
nand U14647 (N_14647,N_12960,N_12106);
xor U14648 (N_14648,N_12328,N_12556);
or U14649 (N_14649,N_13380,N_12793);
and U14650 (N_14650,N_12317,N_12774);
or U14651 (N_14651,N_12135,N_12096);
or U14652 (N_14652,N_12985,N_12910);
nand U14653 (N_14653,N_12374,N_12888);
and U14654 (N_14654,N_12965,N_12303);
nand U14655 (N_14655,N_12338,N_12571);
nor U14656 (N_14656,N_12815,N_13178);
or U14657 (N_14657,N_13379,N_12711);
and U14658 (N_14658,N_12719,N_12260);
and U14659 (N_14659,N_12036,N_13184);
xor U14660 (N_14660,N_12403,N_12377);
nor U14661 (N_14661,N_12582,N_13284);
and U14662 (N_14662,N_13201,N_13466);
and U14663 (N_14663,N_13353,N_13364);
xnor U14664 (N_14664,N_12382,N_13051);
nand U14665 (N_14665,N_13404,N_12163);
nand U14666 (N_14666,N_12773,N_12144);
xor U14667 (N_14667,N_12234,N_13447);
nor U14668 (N_14668,N_12146,N_13021);
xor U14669 (N_14669,N_12920,N_12799);
or U14670 (N_14670,N_12421,N_12803);
nand U14671 (N_14671,N_12397,N_12048);
and U14672 (N_14672,N_12959,N_12282);
nor U14673 (N_14673,N_13485,N_13430);
nand U14674 (N_14674,N_12126,N_12993);
and U14675 (N_14675,N_13357,N_12084);
nor U14676 (N_14676,N_12618,N_13450);
xor U14677 (N_14677,N_13169,N_12710);
nand U14678 (N_14678,N_13389,N_13378);
nand U14679 (N_14679,N_12122,N_12269);
or U14680 (N_14680,N_13439,N_12913);
xor U14681 (N_14681,N_13185,N_12725);
or U14682 (N_14682,N_12023,N_13297);
nand U14683 (N_14683,N_12549,N_13481);
nor U14684 (N_14684,N_12237,N_12185);
nor U14685 (N_14685,N_12008,N_12181);
nand U14686 (N_14686,N_12681,N_12937);
xnor U14687 (N_14687,N_12881,N_12330);
and U14688 (N_14688,N_13310,N_13459);
nand U14689 (N_14689,N_13228,N_13071);
nor U14690 (N_14690,N_12448,N_13488);
and U14691 (N_14691,N_12030,N_12818);
nor U14692 (N_14692,N_12677,N_12225);
nor U14693 (N_14693,N_12079,N_13480);
or U14694 (N_14694,N_12781,N_12856);
nand U14695 (N_14695,N_13318,N_12925);
and U14696 (N_14696,N_12684,N_13300);
nor U14697 (N_14697,N_12738,N_13405);
and U14698 (N_14698,N_12998,N_12652);
or U14699 (N_14699,N_12603,N_12496);
nand U14700 (N_14700,N_13222,N_12544);
or U14701 (N_14701,N_13304,N_12040);
nor U14702 (N_14702,N_13474,N_13150);
and U14703 (N_14703,N_12981,N_12102);
or U14704 (N_14704,N_12052,N_12542);
xnor U14705 (N_14705,N_13495,N_12583);
nand U14706 (N_14706,N_13410,N_13266);
xnor U14707 (N_14707,N_13323,N_13459);
nor U14708 (N_14708,N_12290,N_12746);
or U14709 (N_14709,N_13121,N_12202);
and U14710 (N_14710,N_12169,N_12180);
and U14711 (N_14711,N_12935,N_12922);
nand U14712 (N_14712,N_13411,N_12779);
and U14713 (N_14713,N_13235,N_12219);
and U14714 (N_14714,N_12613,N_12626);
and U14715 (N_14715,N_13358,N_12118);
nor U14716 (N_14716,N_12570,N_13423);
nand U14717 (N_14717,N_13028,N_12600);
xnor U14718 (N_14718,N_12482,N_13201);
nand U14719 (N_14719,N_13083,N_12943);
or U14720 (N_14720,N_12217,N_13471);
nor U14721 (N_14721,N_12400,N_12573);
nor U14722 (N_14722,N_12280,N_13324);
nand U14723 (N_14723,N_13311,N_13247);
or U14724 (N_14724,N_13395,N_12792);
nand U14725 (N_14725,N_12227,N_12973);
nand U14726 (N_14726,N_12974,N_12132);
nand U14727 (N_14727,N_12850,N_13392);
nor U14728 (N_14728,N_12620,N_12333);
nand U14729 (N_14729,N_12767,N_13154);
xnor U14730 (N_14730,N_12675,N_12084);
and U14731 (N_14731,N_13406,N_12018);
and U14732 (N_14732,N_12056,N_13459);
nor U14733 (N_14733,N_12077,N_12555);
nor U14734 (N_14734,N_12465,N_12155);
nor U14735 (N_14735,N_12244,N_12818);
and U14736 (N_14736,N_13259,N_12257);
or U14737 (N_14737,N_12660,N_13307);
nor U14738 (N_14738,N_13490,N_12364);
nand U14739 (N_14739,N_13162,N_13468);
or U14740 (N_14740,N_13427,N_13452);
nand U14741 (N_14741,N_12969,N_13156);
nor U14742 (N_14742,N_12378,N_12443);
nor U14743 (N_14743,N_12396,N_12370);
nor U14744 (N_14744,N_12312,N_12779);
or U14745 (N_14745,N_13346,N_12359);
or U14746 (N_14746,N_12257,N_12423);
or U14747 (N_14747,N_12369,N_12313);
and U14748 (N_14748,N_12727,N_13326);
nand U14749 (N_14749,N_13143,N_12547);
and U14750 (N_14750,N_12477,N_13137);
and U14751 (N_14751,N_12678,N_13218);
or U14752 (N_14752,N_12187,N_13281);
nor U14753 (N_14753,N_12984,N_13280);
nand U14754 (N_14754,N_12112,N_12897);
nand U14755 (N_14755,N_13484,N_13479);
nor U14756 (N_14756,N_12798,N_13088);
xor U14757 (N_14757,N_12015,N_12943);
or U14758 (N_14758,N_12418,N_12959);
nor U14759 (N_14759,N_13055,N_12970);
xor U14760 (N_14760,N_12598,N_12539);
and U14761 (N_14761,N_13425,N_12698);
nor U14762 (N_14762,N_12028,N_13278);
or U14763 (N_14763,N_13253,N_13459);
nor U14764 (N_14764,N_13002,N_12515);
nor U14765 (N_14765,N_12445,N_12691);
nand U14766 (N_14766,N_12973,N_13127);
and U14767 (N_14767,N_12212,N_12032);
or U14768 (N_14768,N_12683,N_13006);
xor U14769 (N_14769,N_13384,N_12177);
or U14770 (N_14770,N_12204,N_12601);
nor U14771 (N_14771,N_12466,N_12422);
and U14772 (N_14772,N_12609,N_12688);
and U14773 (N_14773,N_12714,N_12846);
nand U14774 (N_14774,N_13091,N_12309);
nor U14775 (N_14775,N_12479,N_12881);
and U14776 (N_14776,N_12367,N_12406);
nor U14777 (N_14777,N_13389,N_12770);
and U14778 (N_14778,N_12756,N_12490);
nand U14779 (N_14779,N_13071,N_12449);
or U14780 (N_14780,N_12425,N_13333);
nand U14781 (N_14781,N_12483,N_13279);
and U14782 (N_14782,N_13368,N_13272);
nand U14783 (N_14783,N_13405,N_12573);
and U14784 (N_14784,N_12446,N_12898);
nand U14785 (N_14785,N_12974,N_12542);
and U14786 (N_14786,N_12631,N_12809);
nand U14787 (N_14787,N_13259,N_12972);
or U14788 (N_14788,N_13037,N_12636);
and U14789 (N_14789,N_12941,N_13361);
or U14790 (N_14790,N_13215,N_12674);
nand U14791 (N_14791,N_12193,N_12859);
and U14792 (N_14792,N_12928,N_12304);
nand U14793 (N_14793,N_13072,N_12145);
nand U14794 (N_14794,N_12878,N_12098);
or U14795 (N_14795,N_13356,N_12567);
and U14796 (N_14796,N_13062,N_12589);
or U14797 (N_14797,N_12060,N_13485);
or U14798 (N_14798,N_12251,N_12808);
or U14799 (N_14799,N_12094,N_13353);
nor U14800 (N_14800,N_12899,N_13282);
nor U14801 (N_14801,N_12603,N_12756);
nor U14802 (N_14802,N_12068,N_13048);
nand U14803 (N_14803,N_12598,N_12004);
nor U14804 (N_14804,N_13344,N_12765);
nor U14805 (N_14805,N_12039,N_12263);
and U14806 (N_14806,N_13010,N_12458);
nand U14807 (N_14807,N_12936,N_13441);
and U14808 (N_14808,N_12247,N_13246);
or U14809 (N_14809,N_12758,N_12805);
or U14810 (N_14810,N_12650,N_12764);
and U14811 (N_14811,N_12700,N_12566);
and U14812 (N_14812,N_12038,N_12579);
and U14813 (N_14813,N_12462,N_12031);
nand U14814 (N_14814,N_12001,N_13182);
nor U14815 (N_14815,N_13445,N_12376);
nand U14816 (N_14816,N_13355,N_12436);
and U14817 (N_14817,N_12536,N_12001);
nor U14818 (N_14818,N_13464,N_12954);
and U14819 (N_14819,N_12911,N_12060);
nor U14820 (N_14820,N_13423,N_12492);
and U14821 (N_14821,N_12348,N_12724);
or U14822 (N_14822,N_13136,N_13349);
nor U14823 (N_14823,N_12955,N_13460);
and U14824 (N_14824,N_12113,N_13425);
or U14825 (N_14825,N_12579,N_12685);
nor U14826 (N_14826,N_12928,N_12836);
nand U14827 (N_14827,N_12747,N_13311);
or U14828 (N_14828,N_13221,N_12466);
nand U14829 (N_14829,N_12424,N_13291);
nand U14830 (N_14830,N_13152,N_12038);
xnor U14831 (N_14831,N_13467,N_12332);
nor U14832 (N_14832,N_12738,N_12983);
xor U14833 (N_14833,N_13043,N_13241);
and U14834 (N_14834,N_12425,N_12993);
and U14835 (N_14835,N_12334,N_12384);
nand U14836 (N_14836,N_12593,N_12113);
or U14837 (N_14837,N_12675,N_12527);
and U14838 (N_14838,N_12460,N_12439);
or U14839 (N_14839,N_12942,N_12142);
nor U14840 (N_14840,N_12987,N_13307);
or U14841 (N_14841,N_12755,N_12101);
xnor U14842 (N_14842,N_13024,N_13092);
nor U14843 (N_14843,N_13155,N_12125);
nor U14844 (N_14844,N_12070,N_12463);
or U14845 (N_14845,N_13186,N_12119);
and U14846 (N_14846,N_12810,N_12840);
nand U14847 (N_14847,N_13258,N_12302);
or U14848 (N_14848,N_12336,N_12122);
and U14849 (N_14849,N_12250,N_12044);
and U14850 (N_14850,N_12675,N_12162);
and U14851 (N_14851,N_12722,N_13080);
or U14852 (N_14852,N_13413,N_12647);
nand U14853 (N_14853,N_12612,N_13230);
nand U14854 (N_14854,N_12417,N_12797);
nand U14855 (N_14855,N_13373,N_12849);
nor U14856 (N_14856,N_12245,N_13300);
or U14857 (N_14857,N_13451,N_13260);
xnor U14858 (N_14858,N_12889,N_12087);
or U14859 (N_14859,N_12126,N_12966);
nor U14860 (N_14860,N_13228,N_12288);
or U14861 (N_14861,N_12632,N_12174);
or U14862 (N_14862,N_12271,N_12391);
nor U14863 (N_14863,N_12554,N_12400);
or U14864 (N_14864,N_12902,N_13250);
xor U14865 (N_14865,N_13217,N_13184);
nand U14866 (N_14866,N_12661,N_13485);
nand U14867 (N_14867,N_12462,N_12335);
nor U14868 (N_14868,N_12977,N_12261);
nor U14869 (N_14869,N_13190,N_12885);
and U14870 (N_14870,N_12170,N_12076);
nand U14871 (N_14871,N_12799,N_12241);
or U14872 (N_14872,N_13352,N_12988);
nor U14873 (N_14873,N_12900,N_13370);
or U14874 (N_14874,N_12653,N_13402);
nor U14875 (N_14875,N_12386,N_12130);
and U14876 (N_14876,N_13440,N_13479);
nand U14877 (N_14877,N_12104,N_13435);
nand U14878 (N_14878,N_13008,N_12014);
or U14879 (N_14879,N_12713,N_12104);
nor U14880 (N_14880,N_13376,N_12222);
or U14881 (N_14881,N_13488,N_12755);
nand U14882 (N_14882,N_12421,N_12938);
nand U14883 (N_14883,N_13340,N_12440);
nand U14884 (N_14884,N_13129,N_13442);
and U14885 (N_14885,N_13030,N_12787);
nor U14886 (N_14886,N_12444,N_13163);
and U14887 (N_14887,N_13491,N_13336);
nor U14888 (N_14888,N_12318,N_12866);
and U14889 (N_14889,N_12970,N_12848);
xnor U14890 (N_14890,N_12052,N_13419);
nor U14891 (N_14891,N_12770,N_12776);
nand U14892 (N_14892,N_13051,N_12560);
and U14893 (N_14893,N_12695,N_13314);
nor U14894 (N_14894,N_13207,N_13001);
or U14895 (N_14895,N_13390,N_12984);
nor U14896 (N_14896,N_13100,N_12763);
or U14897 (N_14897,N_12921,N_13280);
nor U14898 (N_14898,N_12917,N_13163);
nor U14899 (N_14899,N_12012,N_12111);
and U14900 (N_14900,N_13126,N_12740);
nor U14901 (N_14901,N_13187,N_12194);
nor U14902 (N_14902,N_12985,N_12770);
nor U14903 (N_14903,N_12598,N_13393);
nand U14904 (N_14904,N_12013,N_13434);
nand U14905 (N_14905,N_12523,N_12861);
and U14906 (N_14906,N_12780,N_13196);
nor U14907 (N_14907,N_12729,N_12475);
nand U14908 (N_14908,N_12897,N_12245);
and U14909 (N_14909,N_12021,N_13111);
and U14910 (N_14910,N_12836,N_13492);
xor U14911 (N_14911,N_12811,N_13290);
xor U14912 (N_14912,N_12400,N_12356);
and U14913 (N_14913,N_12130,N_12780);
or U14914 (N_14914,N_13071,N_13483);
nor U14915 (N_14915,N_13224,N_13440);
and U14916 (N_14916,N_12680,N_12088);
or U14917 (N_14917,N_12978,N_13276);
nand U14918 (N_14918,N_13021,N_12406);
and U14919 (N_14919,N_12604,N_12138);
and U14920 (N_14920,N_13050,N_12302);
and U14921 (N_14921,N_12360,N_13433);
nand U14922 (N_14922,N_13362,N_12821);
nor U14923 (N_14923,N_12107,N_12116);
and U14924 (N_14924,N_12596,N_12254);
nand U14925 (N_14925,N_12084,N_12428);
and U14926 (N_14926,N_13292,N_12048);
or U14927 (N_14927,N_12888,N_12026);
or U14928 (N_14928,N_12608,N_12648);
or U14929 (N_14929,N_13161,N_13193);
xor U14930 (N_14930,N_12950,N_12887);
nor U14931 (N_14931,N_13239,N_13297);
or U14932 (N_14932,N_12888,N_12304);
and U14933 (N_14933,N_12976,N_13440);
xor U14934 (N_14934,N_12632,N_12633);
and U14935 (N_14935,N_12538,N_12840);
or U14936 (N_14936,N_12872,N_12216);
and U14937 (N_14937,N_13175,N_12044);
and U14938 (N_14938,N_13457,N_12563);
nand U14939 (N_14939,N_13257,N_13253);
or U14940 (N_14940,N_12311,N_13300);
or U14941 (N_14941,N_13087,N_12620);
nand U14942 (N_14942,N_12907,N_13138);
nand U14943 (N_14943,N_12695,N_12555);
nand U14944 (N_14944,N_13417,N_13210);
nand U14945 (N_14945,N_12132,N_12230);
nand U14946 (N_14946,N_12163,N_12648);
nand U14947 (N_14947,N_12154,N_12178);
or U14948 (N_14948,N_12284,N_12046);
and U14949 (N_14949,N_13373,N_13258);
or U14950 (N_14950,N_13337,N_12923);
and U14951 (N_14951,N_13042,N_12962);
and U14952 (N_14952,N_12379,N_13115);
xor U14953 (N_14953,N_12338,N_13469);
nand U14954 (N_14954,N_12649,N_12947);
nand U14955 (N_14955,N_12073,N_12854);
or U14956 (N_14956,N_13409,N_12822);
and U14957 (N_14957,N_13375,N_12279);
nand U14958 (N_14958,N_13462,N_12589);
xnor U14959 (N_14959,N_12318,N_12490);
nor U14960 (N_14960,N_12291,N_12196);
nor U14961 (N_14961,N_12295,N_12848);
nor U14962 (N_14962,N_12693,N_13434);
nand U14963 (N_14963,N_13128,N_13235);
nor U14964 (N_14964,N_13318,N_12803);
nor U14965 (N_14965,N_13291,N_12069);
or U14966 (N_14966,N_12315,N_12239);
nor U14967 (N_14967,N_12981,N_12231);
nand U14968 (N_14968,N_13253,N_13126);
and U14969 (N_14969,N_12571,N_12329);
and U14970 (N_14970,N_12492,N_13450);
xor U14971 (N_14971,N_13083,N_13385);
or U14972 (N_14972,N_12062,N_12673);
or U14973 (N_14973,N_12927,N_13128);
nand U14974 (N_14974,N_12767,N_12905);
and U14975 (N_14975,N_12078,N_12915);
nand U14976 (N_14976,N_12266,N_12097);
or U14977 (N_14977,N_12441,N_13480);
or U14978 (N_14978,N_12717,N_13265);
and U14979 (N_14979,N_12855,N_12261);
and U14980 (N_14980,N_12628,N_13408);
nand U14981 (N_14981,N_12073,N_13494);
or U14982 (N_14982,N_12459,N_12763);
nor U14983 (N_14983,N_12817,N_12384);
nand U14984 (N_14984,N_12547,N_13432);
or U14985 (N_14985,N_12543,N_12563);
and U14986 (N_14986,N_12515,N_12622);
and U14987 (N_14987,N_12934,N_12986);
and U14988 (N_14988,N_12409,N_12954);
nor U14989 (N_14989,N_12053,N_12694);
and U14990 (N_14990,N_12577,N_13078);
and U14991 (N_14991,N_12962,N_13403);
xnor U14992 (N_14992,N_12162,N_12907);
or U14993 (N_14993,N_13290,N_13143);
and U14994 (N_14994,N_13451,N_13150);
nor U14995 (N_14995,N_12757,N_12067);
or U14996 (N_14996,N_12285,N_13053);
nand U14997 (N_14997,N_13283,N_12634);
or U14998 (N_14998,N_13353,N_13083);
or U14999 (N_14999,N_13419,N_12359);
nand UO_0 (O_0,N_14103,N_13514);
or UO_1 (O_1,N_14313,N_14271);
nand UO_2 (O_2,N_13710,N_14736);
nor UO_3 (O_3,N_14635,N_13510);
nor UO_4 (O_4,N_14906,N_14037);
or UO_5 (O_5,N_14807,N_14865);
nor UO_6 (O_6,N_14938,N_13521);
xnor UO_7 (O_7,N_13727,N_14274);
nand UO_8 (O_8,N_13706,N_14999);
nor UO_9 (O_9,N_14073,N_14318);
or UO_10 (O_10,N_14117,N_14132);
and UO_11 (O_11,N_14230,N_14581);
or UO_12 (O_12,N_14102,N_13925);
and UO_13 (O_13,N_14530,N_13627);
or UO_14 (O_14,N_14489,N_13705);
nand UO_15 (O_15,N_14410,N_14256);
xor UO_16 (O_16,N_14605,N_14754);
nand UO_17 (O_17,N_13550,N_13578);
nand UO_18 (O_18,N_14782,N_14088);
and UO_19 (O_19,N_13532,N_14294);
nand UO_20 (O_20,N_13573,N_13622);
nor UO_21 (O_21,N_14401,N_13780);
nand UO_22 (O_22,N_14761,N_14273);
and UO_23 (O_23,N_13701,N_14882);
nand UO_24 (O_24,N_14971,N_13534);
nor UO_25 (O_25,N_14074,N_13614);
nor UO_26 (O_26,N_13676,N_14645);
and UO_27 (O_27,N_14300,N_14476);
nand UO_28 (O_28,N_13940,N_13507);
and UO_29 (O_29,N_14198,N_13672);
or UO_30 (O_30,N_14549,N_13973);
and UO_31 (O_31,N_14362,N_13669);
nand UO_32 (O_32,N_13610,N_14125);
and UO_33 (O_33,N_14408,N_14657);
nor UO_34 (O_34,N_14900,N_14350);
nand UO_35 (O_35,N_13520,N_14773);
nor UO_36 (O_36,N_13792,N_14707);
nor UO_37 (O_37,N_13751,N_13882);
nand UO_38 (O_38,N_14646,N_14332);
or UO_39 (O_39,N_14629,N_14021);
and UO_40 (O_40,N_14881,N_14502);
nand UO_41 (O_41,N_14799,N_14993);
or UO_42 (O_42,N_14994,N_14421);
nand UO_43 (O_43,N_14015,N_13778);
or UO_44 (O_44,N_14991,N_13665);
or UO_45 (O_45,N_14439,N_14741);
and UO_46 (O_46,N_14298,N_13768);
nor UO_47 (O_47,N_13581,N_13749);
and UO_48 (O_48,N_14086,N_13640);
nor UO_49 (O_49,N_14727,N_13860);
nor UO_50 (O_50,N_14365,N_14837);
nor UO_51 (O_51,N_13855,N_14307);
or UO_52 (O_52,N_14783,N_13781);
nor UO_53 (O_53,N_14340,N_13689);
nor UO_54 (O_54,N_14995,N_14469);
nand UO_55 (O_55,N_13828,N_13591);
nor UO_56 (O_56,N_13530,N_14739);
nor UO_57 (O_57,N_14732,N_13686);
nor UO_58 (O_58,N_14317,N_14978);
and UO_59 (O_59,N_14441,N_14396);
and UO_60 (O_60,N_13722,N_14763);
and UO_61 (O_61,N_13808,N_14575);
nand UO_62 (O_62,N_14705,N_14531);
nor UO_63 (O_63,N_14291,N_14311);
nand UO_64 (O_64,N_14893,N_14243);
nand UO_65 (O_65,N_14455,N_14566);
or UO_66 (O_66,N_14323,N_14212);
nand UO_67 (O_67,N_14608,N_14505);
nand UO_68 (O_68,N_14159,N_14180);
nand UO_69 (O_69,N_14861,N_14829);
and UO_70 (O_70,N_14589,N_14173);
nor UO_71 (O_71,N_13791,N_14599);
or UO_72 (O_72,N_14265,N_13753);
nor UO_73 (O_73,N_14637,N_13841);
nand UO_74 (O_74,N_13880,N_14299);
or UO_75 (O_75,N_14831,N_14095);
or UO_76 (O_76,N_14667,N_13859);
nand UO_77 (O_77,N_14329,N_13731);
nor UO_78 (O_78,N_14746,N_13748);
nor UO_79 (O_79,N_14022,N_14417);
nand UO_80 (O_80,N_14819,N_14992);
nand UO_81 (O_81,N_13766,N_14312);
or UO_82 (O_82,N_14536,N_13823);
xnor UO_83 (O_83,N_14208,N_13592);
nor UO_84 (O_84,N_13699,N_14945);
nor UO_85 (O_85,N_14356,N_13545);
nor UO_86 (O_86,N_14220,N_14399);
or UO_87 (O_87,N_13990,N_14172);
nand UO_88 (O_88,N_14302,N_14116);
nand UO_89 (O_89,N_13746,N_13715);
nand UO_90 (O_90,N_14135,N_14528);
nand UO_91 (O_91,N_14868,N_14885);
or UO_92 (O_92,N_13915,N_14810);
and UO_93 (O_93,N_14050,N_13836);
nor UO_94 (O_94,N_14260,N_14656);
xnor UO_95 (O_95,N_14788,N_13936);
or UO_96 (O_96,N_14390,N_14328);
nand UO_97 (O_97,N_13683,N_14263);
nor UO_98 (O_98,N_14579,N_14440);
nor UO_99 (O_99,N_13975,N_13724);
nand UO_100 (O_100,N_14631,N_13502);
nor UO_101 (O_101,N_14745,N_14703);
nor UO_102 (O_102,N_13713,N_14675);
nand UO_103 (O_103,N_13541,N_14150);
and UO_104 (O_104,N_13922,N_14163);
xor UO_105 (O_105,N_14368,N_13908);
nor UO_106 (O_106,N_13795,N_13786);
xor UO_107 (O_107,N_14493,N_14169);
nor UO_108 (O_108,N_14008,N_14688);
or UO_109 (O_109,N_13759,N_14082);
or UO_110 (O_110,N_14310,N_14982);
nor UO_111 (O_111,N_14934,N_13983);
nand UO_112 (O_112,N_14834,N_14716);
nor UO_113 (O_113,N_14085,N_14084);
nor UO_114 (O_114,N_14553,N_14551);
nor UO_115 (O_115,N_14935,N_14331);
or UO_116 (O_116,N_14238,N_14953);
nor UO_117 (O_117,N_14869,N_14130);
nor UO_118 (O_118,N_13552,N_13666);
nor UO_119 (O_119,N_14529,N_14558);
and UO_120 (O_120,N_14899,N_13889);
or UO_121 (O_121,N_14278,N_14002);
nand UO_122 (O_122,N_14738,N_14341);
and UO_123 (O_123,N_14149,N_14471);
and UO_124 (O_124,N_14812,N_14460);
or UO_125 (O_125,N_14098,N_13943);
nor UO_126 (O_126,N_14563,N_14670);
nand UO_127 (O_127,N_13799,N_13692);
nor UO_128 (O_128,N_14853,N_13803);
and UO_129 (O_129,N_14509,N_14508);
or UO_130 (O_130,N_13667,N_14973);
and UO_131 (O_131,N_14916,N_14927);
nor UO_132 (O_132,N_13989,N_14977);
or UO_133 (O_133,N_14519,N_14758);
nand UO_134 (O_134,N_13829,N_14663);
and UO_135 (O_135,N_14627,N_14178);
nor UO_136 (O_136,N_14932,N_14018);
and UO_137 (O_137,N_14980,N_14028);
and UO_138 (O_138,N_14570,N_14137);
nor UO_139 (O_139,N_13916,N_13721);
nand UO_140 (O_140,N_14557,N_14501);
or UO_141 (O_141,N_13593,N_14388);
nor UO_142 (O_142,N_13533,N_13563);
nor UO_143 (O_143,N_14258,N_14513);
and UO_144 (O_144,N_14308,N_13760);
nand UO_145 (O_145,N_14418,N_14025);
or UO_146 (O_146,N_14147,N_14956);
or UO_147 (O_147,N_14846,N_13688);
or UO_148 (O_148,N_14468,N_14001);
nand UO_149 (O_149,N_14730,N_14464);
nand UO_150 (O_150,N_14045,N_14912);
and UO_151 (O_151,N_13577,N_14040);
and UO_152 (O_152,N_14038,N_14621);
or UO_153 (O_153,N_14063,N_14897);
or UO_154 (O_154,N_14016,N_14611);
nor UO_155 (O_155,N_14940,N_13546);
nand UO_156 (O_156,N_14620,N_13694);
nor UO_157 (O_157,N_13862,N_14643);
nor UO_158 (O_158,N_13637,N_13516);
nand UO_159 (O_159,N_13921,N_13540);
and UO_160 (O_160,N_13785,N_14477);
nor UO_161 (O_161,N_13805,N_14983);
nor UO_162 (O_162,N_13772,N_14062);
or UO_163 (O_163,N_14106,N_13905);
nor UO_164 (O_164,N_14357,N_13594);
or UO_165 (O_165,N_14077,N_13639);
or UO_166 (O_166,N_14474,N_14032);
xnor UO_167 (O_167,N_14626,N_14111);
nor UO_168 (O_168,N_14504,N_13767);
or UO_169 (O_169,N_13528,N_13869);
xnor UO_170 (O_170,N_13500,N_14600);
nor UO_171 (O_171,N_14876,N_13548);
nand UO_172 (O_172,N_14862,N_14110);
or UO_173 (O_173,N_14237,N_14515);
xor UO_174 (O_174,N_13868,N_13896);
or UO_175 (O_175,N_13560,N_13604);
nand UO_176 (O_176,N_14339,N_14959);
nor UO_177 (O_177,N_13717,N_14485);
and UO_178 (O_178,N_14197,N_13503);
and UO_179 (O_179,N_14510,N_13582);
xnor UO_180 (O_180,N_14400,N_13765);
nor UO_181 (O_181,N_13652,N_14583);
and UO_182 (O_182,N_14261,N_14547);
and UO_183 (O_183,N_14520,N_13903);
and UO_184 (O_184,N_14438,N_14607);
or UO_185 (O_185,N_13920,N_13709);
xor UO_186 (O_186,N_13616,N_14889);
nor UO_187 (O_187,N_14780,N_13901);
or UO_188 (O_188,N_14457,N_13719);
nand UO_189 (O_189,N_14975,N_13917);
nor UO_190 (O_190,N_14678,N_14684);
nand UO_191 (O_191,N_14347,N_14898);
nand UO_192 (O_192,N_14053,N_13877);
or UO_193 (O_193,N_14363,N_14950);
xor UO_194 (O_194,N_14142,N_14448);
nand UO_195 (O_195,N_14896,N_14458);
and UO_196 (O_196,N_14434,N_14380);
nor UO_197 (O_197,N_14718,N_14488);
and UO_198 (O_198,N_14453,N_14473);
nor UO_199 (O_199,N_14686,N_14673);
or UO_200 (O_200,N_14721,N_14955);
and UO_201 (O_201,N_14914,N_14944);
and UO_202 (O_202,N_13586,N_13956);
nand UO_203 (O_203,N_13935,N_14917);
or UO_204 (O_204,N_14574,N_13583);
nand UO_205 (O_205,N_13807,N_14949);
nor UO_206 (O_206,N_13991,N_14648);
and UO_207 (O_207,N_14521,N_14597);
nor UO_208 (O_208,N_13924,N_14036);
or UO_209 (O_209,N_14427,N_13579);
and UO_210 (O_210,N_13839,N_14321);
or UO_211 (O_211,N_14348,N_14630);
and UO_212 (O_212,N_14422,N_14541);
nand UO_213 (O_213,N_14165,N_13512);
or UO_214 (O_214,N_14280,N_13865);
or UO_215 (O_215,N_14405,N_13661);
nor UO_216 (O_216,N_14268,N_14568);
nor UO_217 (O_217,N_14466,N_14325);
and UO_218 (O_218,N_14925,N_13815);
and UO_219 (O_219,N_14090,N_14151);
or UO_220 (O_220,N_14552,N_13971);
nand UO_221 (O_221,N_14289,N_14497);
xnor UO_222 (O_222,N_14722,N_14929);
nor UO_223 (O_223,N_14787,N_14481);
and UO_224 (O_224,N_14044,N_14004);
nand UO_225 (O_225,N_13720,N_13911);
nor UO_226 (O_226,N_14478,N_14437);
or UO_227 (O_227,N_14801,N_14123);
and UO_228 (O_228,N_14857,N_13707);
nor UO_229 (O_229,N_13575,N_13726);
nand UO_230 (O_230,N_14930,N_13831);
and UO_231 (O_231,N_14561,N_13523);
nand UO_232 (O_232,N_14470,N_14669);
nand UO_233 (O_233,N_13856,N_14998);
nand UO_234 (O_234,N_14207,N_13526);
and UO_235 (O_235,N_14231,N_13623);
xor UO_236 (O_236,N_14890,N_14604);
or UO_237 (O_237,N_14072,N_13811);
and UO_238 (O_238,N_14849,N_13761);
nor UO_239 (O_239,N_14818,N_14591);
nand UO_240 (O_240,N_14815,N_14511);
or UO_241 (O_241,N_14776,N_13634);
and UO_242 (O_242,N_14447,N_14742);
nand UO_243 (O_243,N_13564,N_14239);
and UO_244 (O_244,N_13966,N_13848);
or UO_245 (O_245,N_13544,N_13810);
and UO_246 (O_246,N_14413,N_13660);
and UO_247 (O_247,N_13553,N_14548);
or UO_248 (O_248,N_14426,N_13984);
xor UO_249 (O_249,N_14203,N_14115);
nand UO_250 (O_250,N_13702,N_14910);
and UO_251 (O_251,N_14623,N_13685);
xor UO_252 (O_252,N_13601,N_14322);
and UO_253 (O_253,N_14692,N_14976);
nand UO_254 (O_254,N_14080,N_13904);
nand UO_255 (O_255,N_14726,N_13944);
nor UO_256 (O_256,N_14218,N_13976);
or UO_257 (O_257,N_14676,N_13574);
nor UO_258 (O_258,N_14392,N_14498);
or UO_259 (O_259,N_13913,N_14247);
nor UO_260 (O_260,N_14624,N_14847);
or UO_261 (O_261,N_14217,N_14257);
nor UO_262 (O_262,N_13888,N_13840);
nand UO_263 (O_263,N_14068,N_14695);
nor UO_264 (O_264,N_13597,N_14951);
and UO_265 (O_265,N_13682,N_14297);
and UO_266 (O_266,N_14097,N_14444);
and UO_267 (O_267,N_14704,N_14565);
or UO_268 (O_268,N_13513,N_14790);
nor UO_269 (O_269,N_14379,N_14381);
nand UO_270 (O_270,N_13504,N_13568);
nor UO_271 (O_271,N_14843,N_13754);
or UO_272 (O_272,N_13609,N_13764);
and UO_273 (O_273,N_14734,N_14200);
xnor UO_274 (O_274,N_14720,N_14567);
xnor UO_275 (O_275,N_14587,N_14223);
xor UO_276 (O_276,N_13942,N_14324);
and UO_277 (O_277,N_14352,N_14369);
nand UO_278 (O_278,N_14592,N_14006);
xnor UO_279 (O_279,N_13511,N_14081);
nand UO_280 (O_280,N_14586,N_14333);
xor UO_281 (O_281,N_13654,N_14985);
and UO_282 (O_282,N_13775,N_14887);
or UO_283 (O_283,N_14717,N_13851);
nand UO_284 (O_284,N_14618,N_14747);
or UO_285 (O_285,N_14672,N_14997);
and UO_286 (O_286,N_14759,N_14967);
or UO_287 (O_287,N_14491,N_14644);
nor UO_288 (O_288,N_14824,N_14941);
or UO_289 (O_289,N_13804,N_14281);
and UO_290 (O_290,N_13657,N_13641);
and UO_291 (O_291,N_13835,N_14811);
and UO_292 (O_292,N_13946,N_13978);
nand UO_293 (O_293,N_13628,N_13812);
nor UO_294 (O_294,N_14306,N_14674);
nand UO_295 (O_295,N_14507,N_14010);
nand UO_296 (O_296,N_14778,N_14866);
or UO_297 (O_297,N_13571,N_14495);
xor UO_298 (O_298,N_14984,N_14728);
nor UO_299 (O_299,N_13950,N_14245);
xnor UO_300 (O_300,N_14556,N_14284);
or UO_301 (O_301,N_14228,N_14420);
nor UO_302 (O_302,N_14714,N_13501);
nand UO_303 (O_303,N_14192,N_14710);
or UO_304 (O_304,N_13662,N_14139);
and UO_305 (O_305,N_13849,N_13830);
and UO_306 (O_306,N_13963,N_14083);
or UO_307 (O_307,N_13518,N_14595);
nor UO_308 (O_308,N_13827,N_14685);
or UO_309 (O_309,N_14639,N_13615);
nor UO_310 (O_310,N_14562,N_14823);
xnor UO_311 (O_311,N_14743,N_14346);
or UO_312 (O_312,N_14019,N_14908);
nand UO_313 (O_313,N_13525,N_14706);
nand UO_314 (O_314,N_13678,N_13870);
and UO_315 (O_315,N_14054,N_14781);
nand UO_316 (O_316,N_13633,N_13557);
or UO_317 (O_317,N_14891,N_14057);
nor UO_318 (O_318,N_14170,N_13826);
nand UO_319 (O_319,N_14128,N_14250);
nor UO_320 (O_320,N_14569,N_13598);
nor UO_321 (O_321,N_14414,N_13802);
nand UO_322 (O_322,N_13535,N_14406);
nand UO_323 (O_323,N_13522,N_14537);
xor UO_324 (O_324,N_14156,N_14349);
nand UO_325 (O_325,N_14839,N_14337);
nand UO_326 (O_326,N_14576,N_14282);
nor UO_327 (O_327,N_14065,N_13996);
xnor UO_328 (O_328,N_14355,N_13987);
nand UO_329 (O_329,N_14184,N_14248);
nor UO_330 (O_330,N_13673,N_14118);
or UO_331 (O_331,N_14958,N_13900);
nand UO_332 (O_332,N_14012,N_13910);
nand UO_333 (O_333,N_14462,N_13517);
or UO_334 (O_334,N_13524,N_13818);
nor UO_335 (O_335,N_14193,N_14026);
or UO_336 (O_336,N_14385,N_14093);
xnor UO_337 (O_337,N_14628,N_13938);
or UO_338 (O_338,N_14366,N_14735);
nand UO_339 (O_339,N_13585,N_14708);
or UO_340 (O_340,N_13789,N_14969);
nand UO_341 (O_341,N_14484,N_14677);
or UO_342 (O_342,N_13612,N_14603);
nor UO_343 (O_343,N_14211,N_14602);
nor UO_344 (O_344,N_13825,N_14194);
nand UO_345 (O_345,N_14397,N_14451);
or UO_346 (O_346,N_14622,N_14101);
or UO_347 (O_347,N_14126,N_14870);
nor UO_348 (O_348,N_13816,N_13611);
or UO_349 (O_349,N_13708,N_14848);
or UO_350 (O_350,N_14240,N_13626);
nand UO_351 (O_351,N_14749,N_14968);
and UO_352 (O_352,N_13543,N_14543);
xnor UO_353 (O_353,N_14027,N_14506);
and UO_354 (O_354,N_13605,N_13923);
and UO_355 (O_355,N_14697,N_13930);
nand UO_356 (O_356,N_14729,N_14176);
nor UO_357 (O_357,N_13620,N_14965);
nor UO_358 (O_358,N_13907,N_14475);
nand UO_359 (O_359,N_14430,N_14907);
or UO_360 (O_360,N_14472,N_14533);
and UO_361 (O_361,N_13926,N_13677);
nand UO_362 (O_362,N_13890,N_14024);
nor UO_363 (O_363,N_13948,N_13613);
or UO_364 (O_364,N_14540,N_13584);
or UO_365 (O_365,N_13695,N_14903);
or UO_366 (O_366,N_14059,N_14031);
and UO_367 (O_367,N_14376,N_14109);
or UO_368 (O_368,N_13668,N_14058);
and UO_369 (O_369,N_13788,N_14601);
and UO_370 (O_370,N_13687,N_14652);
nor UO_371 (O_371,N_14305,N_14227);
or UO_372 (O_372,N_14500,N_13927);
nor UO_373 (O_373,N_13596,N_14168);
nand UO_374 (O_374,N_13947,N_14793);
nand UO_375 (O_375,N_14161,N_14435);
or UO_376 (O_376,N_14445,N_14241);
or UO_377 (O_377,N_14724,N_13755);
xnor UO_378 (O_378,N_14796,N_13798);
or UO_379 (O_379,N_14658,N_14092);
or UO_380 (O_380,N_13580,N_13783);
xor UO_381 (O_381,N_14210,N_13853);
xnor UO_382 (O_382,N_13891,N_13663);
nor UO_383 (O_383,N_14309,N_13843);
nand UO_384 (O_384,N_14814,N_13842);
and UO_385 (O_385,N_14559,N_14989);
nor UO_386 (O_386,N_13819,N_13752);
nand UO_387 (O_387,N_14661,N_14372);
nand UO_388 (O_388,N_14859,N_14875);
nor UO_389 (O_389,N_13964,N_14377);
nor UO_390 (O_390,N_13995,N_14087);
or UO_391 (O_391,N_14588,N_14554);
nand UO_392 (O_392,N_13732,N_13821);
and UO_393 (O_393,N_13602,N_14733);
nand UO_394 (O_394,N_14785,N_13797);
or UO_395 (O_395,N_14146,N_13897);
or UO_396 (O_396,N_14723,N_13680);
nor UO_397 (O_397,N_13737,N_14610);
nor UO_398 (O_398,N_14696,N_14404);
nor UO_399 (O_399,N_13993,N_14817);
and UO_400 (O_400,N_14216,N_13834);
or UO_401 (O_401,N_14232,N_14872);
xor UO_402 (O_402,N_14415,N_14590);
and UO_403 (O_403,N_14199,N_14775);
and UO_404 (O_404,N_13833,N_14391);
and UO_405 (O_405,N_14972,N_13632);
nor UO_406 (O_406,N_14517,N_14594);
nor UO_407 (O_407,N_14338,N_14113);
nor UO_408 (O_408,N_13728,N_14880);
and UO_409 (O_409,N_14598,N_13782);
nor UO_410 (O_410,N_14030,N_14617);
nor UO_411 (O_411,N_13556,N_14725);
nor UO_412 (O_412,N_14236,N_14664);
xor UO_413 (O_413,N_14525,N_14632);
nor UO_414 (O_414,N_14345,N_14371);
and UO_415 (O_415,N_13902,N_13675);
or UO_416 (O_416,N_14616,N_14296);
nand UO_417 (O_417,N_13527,N_13967);
nand UO_418 (O_418,N_13625,N_14252);
nor UO_419 (O_419,N_14845,N_14655);
or UO_420 (O_420,N_14094,N_14546);
nand UO_421 (O_421,N_13887,N_14167);
and UO_422 (O_422,N_14343,N_14316);
nand UO_423 (O_423,N_13595,N_14071);
and UO_424 (O_424,N_14361,N_14099);
or UO_425 (O_425,N_14091,N_14014);
nor UO_426 (O_426,N_13893,N_13779);
or UO_427 (O_427,N_14432,N_13739);
nand UO_428 (O_428,N_13861,N_14039);
nand UO_429 (O_429,N_14662,N_14544);
nand UO_430 (O_430,N_13992,N_14974);
or UO_431 (O_431,N_14964,N_13740);
nand UO_432 (O_432,N_13847,N_14269);
and UO_433 (O_433,N_14804,N_13969);
nand UO_434 (O_434,N_14936,N_13776);
or UO_435 (O_435,N_14480,N_14336);
or UO_436 (O_436,N_13959,N_13957);
nand UO_437 (O_437,N_13636,N_14879);
or UO_438 (O_438,N_14593,N_14836);
nand UO_439 (O_439,N_14572,N_13820);
nand UO_440 (O_440,N_14794,N_14181);
or UO_441 (O_441,N_14023,N_13747);
nor UO_442 (O_442,N_14942,N_14564);
xnor UO_443 (O_443,N_14254,N_14262);
nor UO_444 (O_444,N_13505,N_13554);
nand UO_445 (O_445,N_14619,N_13757);
nand UO_446 (O_446,N_14690,N_13806);
nand UO_447 (O_447,N_13972,N_13857);
or UO_448 (O_448,N_14049,N_14948);
and UO_449 (O_449,N_14206,N_14699);
nand UO_450 (O_450,N_14774,N_14416);
nor UO_451 (O_451,N_13651,N_14651);
or UO_452 (O_452,N_14826,N_14806);
nand UO_453 (O_453,N_13941,N_14383);
nand UO_454 (O_454,N_14042,N_14808);
nor UO_455 (O_455,N_13712,N_13958);
and UO_456 (O_456,N_14979,N_14850);
and UO_457 (O_457,N_14000,N_13743);
and UO_458 (O_458,N_14913,N_14764);
and UO_459 (O_459,N_14145,N_14768);
nor UO_460 (O_460,N_14403,N_14789);
nor UO_461 (O_461,N_14246,N_14452);
or UO_462 (O_462,N_14459,N_14527);
nand UO_463 (O_463,N_13734,N_13558);
and UO_464 (O_464,N_14209,N_14076);
xnor UO_465 (O_465,N_13960,N_14479);
or UO_466 (O_466,N_14996,N_13872);
or UO_467 (O_467,N_13599,N_14205);
or UO_468 (O_468,N_14104,N_14911);
and UO_469 (O_469,N_14679,N_14360);
xor UO_470 (O_470,N_13933,N_14535);
nand UO_471 (O_471,N_14795,N_14330);
nor UO_472 (O_472,N_14121,N_14382);
or UO_473 (O_473,N_14108,N_14202);
nand UO_474 (O_474,N_13638,N_14970);
xor UO_475 (O_475,N_13875,N_14858);
and UO_476 (O_476,N_14744,N_14467);
nor UO_477 (O_477,N_14926,N_13617);
or UO_478 (O_478,N_14538,N_14671);
nor UO_479 (O_479,N_13733,N_13697);
and UO_480 (O_480,N_14251,N_14204);
or UO_481 (O_481,N_14359,N_14855);
nand UO_482 (O_482,N_13515,N_14921);
and UO_483 (O_483,N_14303,N_14190);
nor UO_484 (O_484,N_13871,N_14020);
nor UO_485 (O_485,N_13878,N_14048);
or UO_486 (O_486,N_13852,N_14825);
or UO_487 (O_487,N_14625,N_14373);
nand UO_488 (O_488,N_14353,N_14143);
nor UO_489 (O_489,N_14140,N_13691);
nand UO_490 (O_490,N_14902,N_13790);
and UO_491 (O_491,N_13693,N_14195);
nor UO_492 (O_492,N_14830,N_13945);
nor UO_493 (O_493,N_13994,N_14089);
or UO_494 (O_494,N_14096,N_13932);
nand UO_495 (O_495,N_14433,N_13906);
nand UO_496 (O_496,N_14275,N_14542);
nand UO_497 (O_497,N_14319,N_13777);
and UO_498 (O_498,N_14351,N_14183);
and UO_499 (O_499,N_13837,N_14918);
and UO_500 (O_500,N_14221,N_14335);
xnor UO_501 (O_501,N_13895,N_13814);
nand UO_502 (O_502,N_14805,N_14043);
nor UO_503 (O_503,N_14047,N_14187);
or UO_504 (O_504,N_14878,N_14841);
xnor UO_505 (O_505,N_14526,N_14107);
and UO_506 (O_506,N_13537,N_14411);
and UO_507 (O_507,N_14755,N_13645);
and UO_508 (O_508,N_14443,N_14753);
xnor UO_509 (O_509,N_14532,N_13809);
nor UO_510 (O_510,N_14842,N_14124);
and UO_511 (O_511,N_14119,N_13542);
nand UO_512 (O_512,N_14874,N_13787);
nor UO_513 (O_513,N_14487,N_14803);
and UO_514 (O_514,N_13674,N_14585);
and UO_515 (O_515,N_13867,N_13624);
nor UO_516 (O_516,N_14387,N_14863);
and UO_517 (O_517,N_14512,N_14370);
and UO_518 (O_518,N_14144,N_14833);
or UO_519 (O_519,N_14152,N_13784);
xor UO_520 (O_520,N_14395,N_13817);
or UO_521 (O_521,N_14719,N_14266);
and UO_522 (O_522,N_14642,N_14154);
nand UO_523 (O_523,N_13649,N_13770);
nand UO_524 (O_524,N_13650,N_14694);
xor UO_525 (O_525,N_14920,N_14293);
and UO_526 (O_526,N_13569,N_14659);
and UO_527 (O_527,N_14270,N_13773);
nand UO_528 (O_528,N_14253,N_13763);
nor UO_529 (O_529,N_13619,N_14055);
and UO_530 (O_530,N_14713,N_13529);
nor UO_531 (O_531,N_13643,N_14954);
nor UO_532 (O_532,N_13653,N_13876);
and UO_533 (O_533,N_14003,N_14374);
or UO_534 (O_534,N_14272,N_14005);
or UO_535 (O_535,N_13647,N_14577);
or UO_536 (O_536,N_14384,N_14687);
or UO_537 (O_537,N_13985,N_13801);
or UO_538 (O_538,N_14981,N_13863);
nand UO_539 (O_539,N_13912,N_14636);
nand UO_540 (O_540,N_14582,N_13725);
nand UO_541 (O_541,N_14769,N_13696);
nand UO_542 (O_542,N_14946,N_14524);
xor UO_543 (O_543,N_14682,N_14215);
or UO_544 (O_544,N_14514,N_13587);
and UO_545 (O_545,N_14813,N_14584);
and UO_546 (O_546,N_13899,N_14233);
and UO_547 (O_547,N_14182,N_14737);
and UO_548 (O_548,N_14762,N_13745);
xnor UO_549 (O_549,N_14409,N_13588);
nor UO_550 (O_550,N_13536,N_14490);
nand UO_551 (O_551,N_14450,N_14650);
or UO_552 (O_552,N_13562,N_13738);
or UO_553 (O_553,N_14786,N_14665);
nor UO_554 (O_554,N_13793,N_13549);
nand UO_555 (O_555,N_14402,N_14522);
or UO_556 (O_556,N_14518,N_14573);
nand UO_557 (O_557,N_14276,N_13873);
nor UO_558 (O_558,N_14820,N_14419);
xor UO_559 (O_559,N_14680,N_14756);
xor UO_560 (O_560,N_14301,N_13886);
xnor UO_561 (O_561,N_14295,N_13965);
or UO_562 (O_562,N_13970,N_13729);
and UO_563 (O_563,N_13703,N_14691);
nor UO_564 (O_564,N_14011,N_14354);
nor UO_565 (O_565,N_14244,N_14449);
nand UO_566 (O_566,N_14066,N_13714);
or UO_567 (O_567,N_14342,N_14131);
nor UO_568 (O_568,N_13919,N_13723);
nand UO_569 (O_569,N_14171,N_13845);
nand UO_570 (O_570,N_13898,N_14873);
nor UO_571 (O_571,N_14185,N_13730);
nand UO_572 (O_572,N_14832,N_14456);
nand UO_573 (O_573,N_14766,N_13644);
xor UO_574 (O_574,N_14653,N_14386);
nor UO_575 (O_575,N_14784,N_14496);
or UO_576 (O_576,N_14668,N_14041);
nand UO_577 (O_577,N_14134,N_13671);
nand UO_578 (O_578,N_13735,N_14314);
nor UO_579 (O_579,N_14864,N_13664);
or UO_580 (O_580,N_13813,N_14436);
nor UO_581 (O_581,N_14867,N_14809);
and UO_582 (O_582,N_13832,N_14122);
or UO_583 (O_583,N_14539,N_13659);
nor UO_584 (O_584,N_13980,N_14499);
and UO_585 (O_585,N_13551,N_13999);
nand UO_586 (O_586,N_13929,N_14904);
xnor UO_587 (O_587,N_14698,N_14064);
xnor UO_588 (O_588,N_13909,N_14943);
nor UO_589 (O_589,N_14700,N_14133);
or UO_590 (O_590,N_14571,N_14153);
and UO_591 (O_591,N_14545,N_14860);
and UO_592 (O_592,N_13988,N_14007);
nor UO_593 (O_593,N_13629,N_14013);
nand UO_594 (O_594,N_13968,N_14654);
nor UO_595 (O_595,N_14127,N_14844);
nand UO_596 (O_596,N_14894,N_14919);
and UO_597 (O_597,N_13952,N_14960);
xor UO_598 (O_598,N_14075,N_13931);
nor UO_599 (O_599,N_14425,N_14196);
nand UO_600 (O_600,N_14884,N_14398);
and UO_601 (O_601,N_14986,N_14229);
nor UO_602 (O_602,N_14748,N_14334);
or UO_603 (O_603,N_13974,N_13934);
xor UO_604 (O_604,N_14923,N_14952);
xnor UO_605 (O_605,N_14905,N_13631);
xnor UO_606 (O_606,N_13892,N_13914);
nand UO_607 (O_607,N_13954,N_14828);
or UO_608 (O_608,N_14871,N_14389);
nor UO_609 (O_609,N_14693,N_14155);
nor UO_610 (O_610,N_13822,N_14492);
nand UO_611 (O_611,N_14056,N_13506);
nor UO_612 (O_612,N_14213,N_14615);
nor UO_613 (O_613,N_13698,N_13606);
xnor UO_614 (O_614,N_14765,N_14606);
and UO_615 (O_615,N_13796,N_14174);
nor UO_616 (O_616,N_13570,N_14214);
nor UO_617 (O_617,N_14711,N_13979);
or UO_618 (O_618,N_14550,N_14883);
and UO_619 (O_619,N_13572,N_14259);
or UO_620 (O_620,N_13736,N_14962);
and UO_621 (O_621,N_14612,N_13590);
xor UO_622 (O_622,N_14375,N_14394);
or UO_623 (O_623,N_14856,N_14990);
nor UO_624 (O_624,N_13603,N_14740);
xor UO_625 (O_625,N_14578,N_14234);
and UO_626 (O_626,N_14290,N_13949);
nor UO_627 (O_627,N_14105,N_14226);
and UO_628 (O_628,N_13607,N_14060);
or UO_629 (O_629,N_13561,N_13918);
nor UO_630 (O_630,N_13928,N_14315);
or UO_631 (O_631,N_14407,N_14798);
nand UO_632 (O_632,N_14660,N_14800);
nand UO_633 (O_633,N_14320,N_14364);
nor UO_634 (O_634,N_14580,N_14757);
nand UO_635 (O_635,N_13742,N_13937);
or UO_636 (O_636,N_14029,N_13681);
or UO_637 (O_637,N_14947,N_13750);
or UO_638 (O_638,N_14560,N_14750);
or UO_639 (O_639,N_14067,N_14177);
or UO_640 (O_640,N_14160,N_14367);
and UO_641 (O_641,N_14327,N_14523);
nand UO_642 (O_642,N_14429,N_14264);
or UO_643 (O_643,N_14933,N_14428);
nor UO_644 (O_644,N_14486,N_14797);
nor UO_645 (O_645,N_14751,N_14821);
nor UO_646 (O_646,N_13700,N_14017);
and UO_647 (O_647,N_14052,N_14596);
xnor UO_648 (O_648,N_14638,N_13850);
or UO_649 (O_649,N_14431,N_14423);
nand UO_650 (O_650,N_14702,N_13716);
or UO_651 (O_651,N_13854,N_14070);
and UO_652 (O_652,N_14640,N_14516);
nand UO_653 (O_653,N_14888,N_14442);
nor UO_654 (O_654,N_14802,N_13670);
and UO_655 (O_655,N_13771,N_13684);
and UO_656 (O_656,N_14033,N_14249);
or UO_657 (O_657,N_14100,N_14358);
nand UO_658 (O_658,N_13576,N_14148);
xnor UO_659 (O_659,N_14069,N_14463);
nor UO_660 (O_660,N_13646,N_14191);
nand UO_661 (O_661,N_14957,N_14009);
and UO_662 (O_662,N_14683,N_14634);
nor UO_663 (O_663,N_13794,N_13883);
nor UO_664 (O_664,N_14393,N_14219);
nor UO_665 (O_665,N_13800,N_13621);
nor UO_666 (O_666,N_14061,N_14827);
and UO_667 (O_667,N_14483,N_14963);
and UO_668 (O_668,N_13565,N_14129);
or UO_669 (O_669,N_13756,N_14141);
nand UO_670 (O_670,N_14175,N_14854);
nand UO_671 (O_671,N_13953,N_14966);
nand UO_672 (O_672,N_14901,N_14136);
nor UO_673 (O_673,N_13961,N_14378);
nor UO_674 (O_674,N_13986,N_14835);
nand UO_675 (O_675,N_14731,N_14852);
or UO_676 (O_676,N_14816,N_13718);
or UO_677 (O_677,N_14461,N_13656);
xor UO_678 (O_678,N_13858,N_14112);
nor UO_679 (O_679,N_14689,N_14166);
nor UO_680 (O_680,N_14701,N_14051);
or UO_681 (O_681,N_13509,N_14189);
or UO_682 (O_682,N_14779,N_13589);
nor UO_683 (O_683,N_13874,N_13655);
and UO_684 (O_684,N_13951,N_14482);
xor UO_685 (O_685,N_13866,N_14712);
and UO_686 (O_686,N_14928,N_13838);
and UO_687 (O_687,N_14162,N_13600);
or UO_688 (O_688,N_14222,N_13962);
nand UO_689 (O_689,N_13955,N_14915);
xor UO_690 (O_690,N_14851,N_14225);
xnor UO_691 (O_691,N_14503,N_14078);
xnor UO_692 (O_692,N_14715,N_14292);
and UO_693 (O_693,N_14034,N_13894);
nor UO_694 (O_694,N_13998,N_13538);
or UO_695 (O_695,N_14681,N_14709);
and UO_696 (O_696,N_13881,N_13758);
xor UO_697 (O_697,N_13555,N_14188);
nor UO_698 (O_698,N_13679,N_14424);
nor UO_699 (O_699,N_13885,N_13658);
or UO_700 (O_700,N_14201,N_13690);
and UO_701 (O_701,N_14158,N_14288);
or UO_702 (O_702,N_14922,N_13547);
xor UO_703 (O_703,N_14924,N_13567);
nand UO_704 (O_704,N_13774,N_13508);
nor UO_705 (O_705,N_14412,N_14840);
or UO_706 (O_706,N_13762,N_13741);
or UO_707 (O_707,N_14283,N_14792);
and UO_708 (O_708,N_14242,N_14609);
nand UO_709 (O_709,N_14344,N_14649);
nand UO_710 (O_710,N_14120,N_14079);
nand UO_711 (O_711,N_13630,N_13864);
and UO_712 (O_712,N_14186,N_13884);
nor UO_713 (O_713,N_14877,N_13559);
xor UO_714 (O_714,N_14285,N_14822);
or UO_715 (O_715,N_14647,N_14224);
and UO_716 (O_716,N_14138,N_14035);
or UO_717 (O_717,N_14895,N_13982);
and UO_718 (O_718,N_14279,N_14454);
nor UO_719 (O_719,N_13744,N_13846);
and UO_720 (O_720,N_13566,N_13939);
and UO_721 (O_721,N_14446,N_14752);
or UO_722 (O_722,N_14939,N_13824);
nand UO_723 (O_723,N_14760,N_14287);
nand UO_724 (O_724,N_14937,N_14931);
or UO_725 (O_725,N_13635,N_14613);
nor UO_726 (O_726,N_14465,N_14886);
nand UO_727 (O_727,N_14909,N_14791);
nand UO_728 (O_728,N_13977,N_13519);
nand UO_729 (O_729,N_14770,N_13608);
and UO_730 (O_730,N_14772,N_14164);
nor UO_731 (O_731,N_13539,N_14179);
and UO_732 (O_732,N_13531,N_14555);
nor UO_733 (O_733,N_14534,N_14235);
nor UO_734 (O_734,N_13618,N_14046);
nor UO_735 (O_735,N_14838,N_14961);
and UO_736 (O_736,N_14114,N_13648);
nor UO_737 (O_737,N_14771,N_14777);
and UO_738 (O_738,N_13844,N_14326);
nand UO_739 (O_739,N_14304,N_14267);
nor UO_740 (O_740,N_14157,N_14767);
and UO_741 (O_741,N_14641,N_13981);
and UO_742 (O_742,N_14987,N_13879);
xor UO_743 (O_743,N_13642,N_13997);
nor UO_744 (O_744,N_13769,N_14633);
or UO_745 (O_745,N_13711,N_14255);
or UO_746 (O_746,N_14494,N_14614);
nor UO_747 (O_747,N_14988,N_14666);
nor UO_748 (O_748,N_14277,N_14892);
and UO_749 (O_749,N_14286,N_13704);
and UO_750 (O_750,N_14606,N_13919);
or UO_751 (O_751,N_14029,N_14365);
nand UO_752 (O_752,N_13662,N_13905);
nand UO_753 (O_753,N_14909,N_14420);
and UO_754 (O_754,N_14347,N_14742);
or UO_755 (O_755,N_14960,N_13609);
nor UO_756 (O_756,N_14237,N_13530);
nand UO_757 (O_757,N_14946,N_14135);
nand UO_758 (O_758,N_14200,N_13849);
nand UO_759 (O_759,N_14599,N_14461);
and UO_760 (O_760,N_14935,N_14126);
and UO_761 (O_761,N_13548,N_13811);
and UO_762 (O_762,N_13864,N_14892);
nand UO_763 (O_763,N_14430,N_14511);
or UO_764 (O_764,N_14433,N_13676);
or UO_765 (O_765,N_13772,N_13608);
and UO_766 (O_766,N_14404,N_13551);
or UO_767 (O_767,N_13835,N_14724);
xor UO_768 (O_768,N_13627,N_14941);
and UO_769 (O_769,N_13759,N_13528);
or UO_770 (O_770,N_14045,N_14561);
nand UO_771 (O_771,N_13714,N_13738);
nor UO_772 (O_772,N_14432,N_13773);
or UO_773 (O_773,N_13529,N_14722);
nand UO_774 (O_774,N_13570,N_14875);
and UO_775 (O_775,N_14629,N_14576);
nand UO_776 (O_776,N_14127,N_14910);
or UO_777 (O_777,N_13845,N_14727);
nor UO_778 (O_778,N_14815,N_14451);
or UO_779 (O_779,N_13877,N_14597);
and UO_780 (O_780,N_14376,N_13630);
nand UO_781 (O_781,N_14470,N_14916);
xnor UO_782 (O_782,N_14487,N_13779);
nand UO_783 (O_783,N_13866,N_14524);
and UO_784 (O_784,N_13820,N_14392);
xnor UO_785 (O_785,N_14957,N_14264);
or UO_786 (O_786,N_14002,N_13930);
or UO_787 (O_787,N_14391,N_13644);
nor UO_788 (O_788,N_14593,N_13975);
nor UO_789 (O_789,N_13512,N_14552);
nor UO_790 (O_790,N_14131,N_14867);
nand UO_791 (O_791,N_14817,N_14813);
and UO_792 (O_792,N_14849,N_13639);
or UO_793 (O_793,N_14408,N_13531);
and UO_794 (O_794,N_14473,N_13585);
and UO_795 (O_795,N_13610,N_14887);
nor UO_796 (O_796,N_13755,N_13954);
and UO_797 (O_797,N_14071,N_14172);
and UO_798 (O_798,N_14869,N_14995);
or UO_799 (O_799,N_14875,N_14487);
or UO_800 (O_800,N_13728,N_14866);
nand UO_801 (O_801,N_14257,N_14383);
or UO_802 (O_802,N_14709,N_14568);
and UO_803 (O_803,N_13672,N_14543);
nand UO_804 (O_804,N_14623,N_14989);
or UO_805 (O_805,N_14843,N_14511);
or UO_806 (O_806,N_13906,N_13597);
xnor UO_807 (O_807,N_14756,N_13866);
nor UO_808 (O_808,N_13898,N_14396);
and UO_809 (O_809,N_14842,N_13804);
and UO_810 (O_810,N_13648,N_14058);
and UO_811 (O_811,N_14041,N_14538);
or UO_812 (O_812,N_14022,N_14259);
or UO_813 (O_813,N_14523,N_14266);
or UO_814 (O_814,N_13690,N_14518);
or UO_815 (O_815,N_13965,N_14727);
nand UO_816 (O_816,N_13768,N_13884);
or UO_817 (O_817,N_13731,N_13647);
nand UO_818 (O_818,N_14729,N_14523);
nor UO_819 (O_819,N_14153,N_13996);
nor UO_820 (O_820,N_13987,N_14783);
and UO_821 (O_821,N_14835,N_14635);
or UO_822 (O_822,N_13911,N_14616);
nor UO_823 (O_823,N_14354,N_13596);
nor UO_824 (O_824,N_14187,N_13533);
nand UO_825 (O_825,N_13789,N_13984);
and UO_826 (O_826,N_14379,N_14468);
or UO_827 (O_827,N_13675,N_14528);
nand UO_828 (O_828,N_14021,N_14149);
xnor UO_829 (O_829,N_14167,N_14445);
nand UO_830 (O_830,N_14708,N_14835);
and UO_831 (O_831,N_14299,N_13580);
or UO_832 (O_832,N_13523,N_14414);
nand UO_833 (O_833,N_14704,N_14195);
nand UO_834 (O_834,N_14810,N_13720);
and UO_835 (O_835,N_14012,N_14042);
nor UO_836 (O_836,N_14545,N_14829);
nand UO_837 (O_837,N_14499,N_13620);
and UO_838 (O_838,N_14564,N_14123);
nor UO_839 (O_839,N_13740,N_14260);
or UO_840 (O_840,N_14629,N_14157);
nand UO_841 (O_841,N_14627,N_14976);
nor UO_842 (O_842,N_13564,N_13996);
nand UO_843 (O_843,N_14933,N_14426);
nor UO_844 (O_844,N_13644,N_13895);
xnor UO_845 (O_845,N_14394,N_14697);
and UO_846 (O_846,N_13937,N_13954);
nor UO_847 (O_847,N_14176,N_14410);
and UO_848 (O_848,N_14716,N_14253);
or UO_849 (O_849,N_13578,N_14659);
nand UO_850 (O_850,N_14110,N_13782);
or UO_851 (O_851,N_14687,N_13928);
nor UO_852 (O_852,N_14245,N_13641);
xnor UO_853 (O_853,N_14242,N_14501);
and UO_854 (O_854,N_13638,N_14346);
xor UO_855 (O_855,N_14868,N_13828);
and UO_856 (O_856,N_14828,N_14136);
nand UO_857 (O_857,N_14307,N_13813);
or UO_858 (O_858,N_13548,N_14535);
or UO_859 (O_859,N_14100,N_13818);
nor UO_860 (O_860,N_13890,N_14474);
or UO_861 (O_861,N_13953,N_13836);
nor UO_862 (O_862,N_13830,N_14348);
or UO_863 (O_863,N_14003,N_13751);
nand UO_864 (O_864,N_14234,N_14973);
nand UO_865 (O_865,N_13634,N_14413);
nand UO_866 (O_866,N_14059,N_14154);
nor UO_867 (O_867,N_14213,N_13716);
and UO_868 (O_868,N_14902,N_13817);
and UO_869 (O_869,N_14744,N_14820);
nor UO_870 (O_870,N_14616,N_14716);
xnor UO_871 (O_871,N_14540,N_13858);
xor UO_872 (O_872,N_13814,N_14067);
nand UO_873 (O_873,N_13843,N_14315);
or UO_874 (O_874,N_14564,N_14525);
or UO_875 (O_875,N_14189,N_13639);
or UO_876 (O_876,N_13955,N_13662);
or UO_877 (O_877,N_14891,N_14955);
xor UO_878 (O_878,N_13935,N_14099);
xor UO_879 (O_879,N_14253,N_14981);
xor UO_880 (O_880,N_13953,N_14211);
and UO_881 (O_881,N_14345,N_13973);
or UO_882 (O_882,N_13937,N_14473);
nor UO_883 (O_883,N_13981,N_14670);
or UO_884 (O_884,N_14809,N_14877);
or UO_885 (O_885,N_13949,N_13883);
or UO_886 (O_886,N_14271,N_14283);
nor UO_887 (O_887,N_14745,N_14063);
nor UO_888 (O_888,N_14600,N_14148);
or UO_889 (O_889,N_13512,N_13591);
or UO_890 (O_890,N_13621,N_13760);
or UO_891 (O_891,N_13602,N_13990);
nor UO_892 (O_892,N_14270,N_14495);
nand UO_893 (O_893,N_14561,N_13941);
or UO_894 (O_894,N_14643,N_14453);
or UO_895 (O_895,N_14726,N_14479);
nor UO_896 (O_896,N_13724,N_13749);
and UO_897 (O_897,N_14478,N_14206);
or UO_898 (O_898,N_14256,N_13865);
nor UO_899 (O_899,N_14169,N_14123);
and UO_900 (O_900,N_13982,N_14199);
and UO_901 (O_901,N_14663,N_14064);
nand UO_902 (O_902,N_14966,N_14071);
nor UO_903 (O_903,N_13616,N_14212);
and UO_904 (O_904,N_14035,N_14638);
and UO_905 (O_905,N_14586,N_14620);
and UO_906 (O_906,N_14438,N_14094);
or UO_907 (O_907,N_13505,N_13541);
and UO_908 (O_908,N_14730,N_14256);
nand UO_909 (O_909,N_14251,N_13969);
nand UO_910 (O_910,N_14142,N_14359);
nor UO_911 (O_911,N_13553,N_13796);
or UO_912 (O_912,N_13994,N_14011);
nor UO_913 (O_913,N_14607,N_13805);
nor UO_914 (O_914,N_14539,N_13569);
and UO_915 (O_915,N_14177,N_13796);
nand UO_916 (O_916,N_14406,N_13941);
nor UO_917 (O_917,N_14409,N_13670);
and UO_918 (O_918,N_14632,N_14421);
and UO_919 (O_919,N_13993,N_14588);
and UO_920 (O_920,N_13678,N_13962);
or UO_921 (O_921,N_14798,N_14064);
xor UO_922 (O_922,N_14819,N_14773);
nor UO_923 (O_923,N_14509,N_14278);
xor UO_924 (O_924,N_14544,N_13621);
nor UO_925 (O_925,N_13727,N_14453);
nor UO_926 (O_926,N_14894,N_13670);
xnor UO_927 (O_927,N_13962,N_13612);
and UO_928 (O_928,N_14477,N_13960);
or UO_929 (O_929,N_13612,N_14071);
nand UO_930 (O_930,N_14700,N_13515);
and UO_931 (O_931,N_14527,N_14189);
xor UO_932 (O_932,N_13799,N_14903);
nor UO_933 (O_933,N_13906,N_13644);
and UO_934 (O_934,N_14170,N_14479);
and UO_935 (O_935,N_13592,N_14397);
and UO_936 (O_936,N_13712,N_13804);
and UO_937 (O_937,N_14927,N_14594);
and UO_938 (O_938,N_14991,N_13720);
or UO_939 (O_939,N_13978,N_14453);
nor UO_940 (O_940,N_14710,N_14347);
nor UO_941 (O_941,N_13964,N_14878);
xor UO_942 (O_942,N_14418,N_13616);
nor UO_943 (O_943,N_14055,N_13784);
xor UO_944 (O_944,N_14443,N_14457);
nand UO_945 (O_945,N_14337,N_14170);
nor UO_946 (O_946,N_13645,N_13547);
nand UO_947 (O_947,N_14589,N_13565);
nor UO_948 (O_948,N_13664,N_14758);
nor UO_949 (O_949,N_13771,N_14146);
and UO_950 (O_950,N_14629,N_14046);
nor UO_951 (O_951,N_14688,N_13547);
or UO_952 (O_952,N_13705,N_13918);
and UO_953 (O_953,N_14846,N_13905);
nor UO_954 (O_954,N_14990,N_14726);
and UO_955 (O_955,N_13887,N_14466);
or UO_956 (O_956,N_14744,N_14733);
and UO_957 (O_957,N_14774,N_14397);
or UO_958 (O_958,N_14427,N_14041);
nor UO_959 (O_959,N_14021,N_13594);
and UO_960 (O_960,N_14730,N_14887);
and UO_961 (O_961,N_13590,N_14212);
nand UO_962 (O_962,N_14368,N_13790);
nor UO_963 (O_963,N_13670,N_14389);
and UO_964 (O_964,N_14571,N_14882);
nor UO_965 (O_965,N_14953,N_13964);
or UO_966 (O_966,N_14092,N_14308);
or UO_967 (O_967,N_14619,N_14004);
nand UO_968 (O_968,N_14052,N_14680);
and UO_969 (O_969,N_14352,N_14785);
nor UO_970 (O_970,N_14944,N_14649);
nor UO_971 (O_971,N_14617,N_13530);
or UO_972 (O_972,N_14547,N_14895);
nor UO_973 (O_973,N_14481,N_13605);
nand UO_974 (O_974,N_14695,N_13586);
xnor UO_975 (O_975,N_14667,N_14421);
nand UO_976 (O_976,N_14308,N_13603);
and UO_977 (O_977,N_14655,N_13861);
and UO_978 (O_978,N_14939,N_14699);
and UO_979 (O_979,N_14113,N_14711);
xnor UO_980 (O_980,N_13686,N_14418);
xor UO_981 (O_981,N_14147,N_13854);
nand UO_982 (O_982,N_13777,N_14336);
or UO_983 (O_983,N_13511,N_14591);
xnor UO_984 (O_984,N_14507,N_14114);
or UO_985 (O_985,N_14385,N_14495);
nand UO_986 (O_986,N_13869,N_13876);
nand UO_987 (O_987,N_13615,N_14558);
nor UO_988 (O_988,N_14253,N_13662);
or UO_989 (O_989,N_13625,N_14942);
or UO_990 (O_990,N_14337,N_14594);
or UO_991 (O_991,N_14773,N_14085);
and UO_992 (O_992,N_14754,N_14159);
and UO_993 (O_993,N_14363,N_14673);
or UO_994 (O_994,N_14298,N_14322);
nor UO_995 (O_995,N_13517,N_13892);
nor UO_996 (O_996,N_13523,N_13991);
nand UO_997 (O_997,N_14539,N_14943);
nand UO_998 (O_998,N_13644,N_14969);
nand UO_999 (O_999,N_14418,N_14738);
xor UO_1000 (O_1000,N_13995,N_13985);
nor UO_1001 (O_1001,N_14168,N_14184);
nor UO_1002 (O_1002,N_14682,N_13674);
nor UO_1003 (O_1003,N_13592,N_14429);
nand UO_1004 (O_1004,N_14835,N_14887);
nor UO_1005 (O_1005,N_14521,N_14931);
and UO_1006 (O_1006,N_14220,N_14442);
nor UO_1007 (O_1007,N_14291,N_14437);
nand UO_1008 (O_1008,N_14510,N_14214);
nor UO_1009 (O_1009,N_14690,N_14622);
nand UO_1010 (O_1010,N_14430,N_14866);
xnor UO_1011 (O_1011,N_14015,N_14952);
nand UO_1012 (O_1012,N_14134,N_14240);
nand UO_1013 (O_1013,N_13879,N_14983);
and UO_1014 (O_1014,N_13651,N_13574);
nand UO_1015 (O_1015,N_13651,N_14177);
nand UO_1016 (O_1016,N_14111,N_14463);
or UO_1017 (O_1017,N_13800,N_14723);
nor UO_1018 (O_1018,N_14593,N_14429);
xnor UO_1019 (O_1019,N_14671,N_14283);
and UO_1020 (O_1020,N_14013,N_14698);
nand UO_1021 (O_1021,N_14812,N_14636);
and UO_1022 (O_1022,N_14556,N_14083);
and UO_1023 (O_1023,N_14188,N_13720);
xnor UO_1024 (O_1024,N_14505,N_14245);
nand UO_1025 (O_1025,N_14878,N_13867);
and UO_1026 (O_1026,N_14974,N_14585);
or UO_1027 (O_1027,N_13712,N_13600);
xnor UO_1028 (O_1028,N_14265,N_13719);
nand UO_1029 (O_1029,N_14281,N_13687);
nor UO_1030 (O_1030,N_13607,N_14156);
nor UO_1031 (O_1031,N_13632,N_14448);
nand UO_1032 (O_1032,N_13760,N_14405);
xnor UO_1033 (O_1033,N_14745,N_13776);
xnor UO_1034 (O_1034,N_13975,N_14741);
or UO_1035 (O_1035,N_14032,N_14552);
and UO_1036 (O_1036,N_14201,N_14596);
or UO_1037 (O_1037,N_14573,N_14763);
nor UO_1038 (O_1038,N_14359,N_13762);
xnor UO_1039 (O_1039,N_14368,N_13711);
and UO_1040 (O_1040,N_14557,N_14350);
nor UO_1041 (O_1041,N_13527,N_14289);
nor UO_1042 (O_1042,N_14361,N_14355);
nand UO_1043 (O_1043,N_13861,N_14103);
nor UO_1044 (O_1044,N_13594,N_14615);
nand UO_1045 (O_1045,N_14349,N_14450);
nand UO_1046 (O_1046,N_13643,N_13871);
nand UO_1047 (O_1047,N_14193,N_14230);
nand UO_1048 (O_1048,N_14720,N_14305);
nand UO_1049 (O_1049,N_14227,N_14450);
nor UO_1050 (O_1050,N_13811,N_14418);
nor UO_1051 (O_1051,N_13910,N_14920);
xor UO_1052 (O_1052,N_14303,N_14171);
and UO_1053 (O_1053,N_14045,N_13600);
or UO_1054 (O_1054,N_14419,N_14825);
nand UO_1055 (O_1055,N_14032,N_13728);
and UO_1056 (O_1056,N_14524,N_14858);
and UO_1057 (O_1057,N_14750,N_14428);
and UO_1058 (O_1058,N_14118,N_14539);
nand UO_1059 (O_1059,N_13509,N_13908);
or UO_1060 (O_1060,N_14853,N_14055);
and UO_1061 (O_1061,N_14505,N_13610);
xor UO_1062 (O_1062,N_14765,N_14007);
nand UO_1063 (O_1063,N_14118,N_13655);
nor UO_1064 (O_1064,N_14560,N_13935);
nand UO_1065 (O_1065,N_14524,N_14761);
nor UO_1066 (O_1066,N_14584,N_13912);
or UO_1067 (O_1067,N_14178,N_13780);
and UO_1068 (O_1068,N_14766,N_13975);
nand UO_1069 (O_1069,N_14172,N_14058);
nor UO_1070 (O_1070,N_14985,N_14269);
xor UO_1071 (O_1071,N_14949,N_14186);
nor UO_1072 (O_1072,N_14022,N_14056);
or UO_1073 (O_1073,N_13776,N_13566);
or UO_1074 (O_1074,N_14217,N_13911);
nor UO_1075 (O_1075,N_14765,N_13511);
nor UO_1076 (O_1076,N_14840,N_14941);
nand UO_1077 (O_1077,N_14258,N_14559);
or UO_1078 (O_1078,N_14368,N_14968);
nor UO_1079 (O_1079,N_14392,N_13673);
nand UO_1080 (O_1080,N_13766,N_14802);
or UO_1081 (O_1081,N_14730,N_14115);
nor UO_1082 (O_1082,N_13902,N_13684);
nor UO_1083 (O_1083,N_13574,N_14310);
nor UO_1084 (O_1084,N_14317,N_13920);
nor UO_1085 (O_1085,N_14758,N_13823);
nor UO_1086 (O_1086,N_13718,N_13662);
nand UO_1087 (O_1087,N_13514,N_13734);
nor UO_1088 (O_1088,N_14988,N_14078);
and UO_1089 (O_1089,N_14554,N_14172);
and UO_1090 (O_1090,N_13599,N_13982);
xor UO_1091 (O_1091,N_13745,N_14961);
and UO_1092 (O_1092,N_14417,N_14221);
nor UO_1093 (O_1093,N_14381,N_13735);
or UO_1094 (O_1094,N_14748,N_13888);
or UO_1095 (O_1095,N_13907,N_14809);
nor UO_1096 (O_1096,N_13959,N_14965);
nor UO_1097 (O_1097,N_13690,N_14321);
nor UO_1098 (O_1098,N_14490,N_14350);
or UO_1099 (O_1099,N_14325,N_14551);
and UO_1100 (O_1100,N_14844,N_14955);
or UO_1101 (O_1101,N_14564,N_14487);
and UO_1102 (O_1102,N_14678,N_14304);
nor UO_1103 (O_1103,N_14406,N_13832);
or UO_1104 (O_1104,N_14647,N_13582);
nor UO_1105 (O_1105,N_14083,N_13574);
nand UO_1106 (O_1106,N_14395,N_14714);
and UO_1107 (O_1107,N_14502,N_13840);
and UO_1108 (O_1108,N_14159,N_13555);
and UO_1109 (O_1109,N_13634,N_13771);
and UO_1110 (O_1110,N_14473,N_13786);
and UO_1111 (O_1111,N_14991,N_13986);
nand UO_1112 (O_1112,N_13682,N_13942);
or UO_1113 (O_1113,N_13736,N_13638);
nor UO_1114 (O_1114,N_14587,N_14891);
nor UO_1115 (O_1115,N_14758,N_14165);
nor UO_1116 (O_1116,N_14554,N_14700);
nand UO_1117 (O_1117,N_14542,N_14117);
or UO_1118 (O_1118,N_14809,N_13607);
nand UO_1119 (O_1119,N_14313,N_14715);
nor UO_1120 (O_1120,N_14225,N_13507);
or UO_1121 (O_1121,N_14129,N_14668);
nand UO_1122 (O_1122,N_13586,N_14206);
and UO_1123 (O_1123,N_14183,N_14762);
xnor UO_1124 (O_1124,N_14152,N_14708);
nor UO_1125 (O_1125,N_14564,N_14584);
nand UO_1126 (O_1126,N_14289,N_14223);
or UO_1127 (O_1127,N_13638,N_14532);
or UO_1128 (O_1128,N_14005,N_14765);
or UO_1129 (O_1129,N_13596,N_14193);
nor UO_1130 (O_1130,N_14410,N_14295);
nand UO_1131 (O_1131,N_13841,N_14340);
or UO_1132 (O_1132,N_14613,N_14815);
nor UO_1133 (O_1133,N_13603,N_14971);
and UO_1134 (O_1134,N_14673,N_14084);
nand UO_1135 (O_1135,N_14003,N_14663);
or UO_1136 (O_1136,N_14240,N_13796);
xor UO_1137 (O_1137,N_14414,N_14009);
nand UO_1138 (O_1138,N_14008,N_13698);
and UO_1139 (O_1139,N_13606,N_14348);
nand UO_1140 (O_1140,N_13969,N_13917);
or UO_1141 (O_1141,N_14181,N_13513);
and UO_1142 (O_1142,N_14088,N_14892);
nor UO_1143 (O_1143,N_14074,N_13695);
and UO_1144 (O_1144,N_14694,N_13540);
or UO_1145 (O_1145,N_14483,N_14845);
nand UO_1146 (O_1146,N_14194,N_13844);
nand UO_1147 (O_1147,N_14692,N_14062);
nor UO_1148 (O_1148,N_14817,N_14195);
or UO_1149 (O_1149,N_14049,N_14097);
xnor UO_1150 (O_1150,N_13834,N_14361);
nand UO_1151 (O_1151,N_14955,N_14251);
or UO_1152 (O_1152,N_14022,N_13575);
and UO_1153 (O_1153,N_14240,N_13833);
or UO_1154 (O_1154,N_13753,N_13647);
and UO_1155 (O_1155,N_14948,N_14878);
nor UO_1156 (O_1156,N_14781,N_14333);
or UO_1157 (O_1157,N_13811,N_13601);
and UO_1158 (O_1158,N_13914,N_13581);
and UO_1159 (O_1159,N_13820,N_13805);
or UO_1160 (O_1160,N_14628,N_14442);
nor UO_1161 (O_1161,N_14823,N_13824);
nand UO_1162 (O_1162,N_14202,N_14714);
and UO_1163 (O_1163,N_14045,N_14456);
or UO_1164 (O_1164,N_14963,N_13573);
or UO_1165 (O_1165,N_14714,N_14577);
or UO_1166 (O_1166,N_14845,N_13917);
and UO_1167 (O_1167,N_14333,N_13847);
nor UO_1168 (O_1168,N_14460,N_14709);
and UO_1169 (O_1169,N_14599,N_14646);
nand UO_1170 (O_1170,N_14006,N_14570);
nand UO_1171 (O_1171,N_14860,N_13677);
or UO_1172 (O_1172,N_13501,N_13718);
or UO_1173 (O_1173,N_14261,N_14675);
or UO_1174 (O_1174,N_14218,N_14884);
nand UO_1175 (O_1175,N_13831,N_14611);
or UO_1176 (O_1176,N_14885,N_14125);
nor UO_1177 (O_1177,N_13548,N_13893);
and UO_1178 (O_1178,N_14741,N_13774);
xor UO_1179 (O_1179,N_13922,N_14126);
nand UO_1180 (O_1180,N_13719,N_14743);
nand UO_1181 (O_1181,N_14242,N_14037);
or UO_1182 (O_1182,N_13830,N_13521);
and UO_1183 (O_1183,N_13593,N_14965);
nor UO_1184 (O_1184,N_14977,N_14238);
nor UO_1185 (O_1185,N_14964,N_14298);
nor UO_1186 (O_1186,N_14290,N_14092);
nand UO_1187 (O_1187,N_14301,N_14154);
or UO_1188 (O_1188,N_14250,N_14144);
nor UO_1189 (O_1189,N_14190,N_14729);
xnor UO_1190 (O_1190,N_13651,N_13924);
xor UO_1191 (O_1191,N_14879,N_14126);
and UO_1192 (O_1192,N_13847,N_14007);
and UO_1193 (O_1193,N_14731,N_13510);
or UO_1194 (O_1194,N_13897,N_14207);
nand UO_1195 (O_1195,N_14920,N_13623);
nand UO_1196 (O_1196,N_14668,N_14037);
nor UO_1197 (O_1197,N_14943,N_14828);
nor UO_1198 (O_1198,N_14618,N_13902);
nor UO_1199 (O_1199,N_14363,N_14116);
or UO_1200 (O_1200,N_13582,N_13855);
xor UO_1201 (O_1201,N_13825,N_13851);
or UO_1202 (O_1202,N_14986,N_13599);
or UO_1203 (O_1203,N_14903,N_14849);
nor UO_1204 (O_1204,N_13705,N_14610);
xnor UO_1205 (O_1205,N_14828,N_14225);
nor UO_1206 (O_1206,N_14338,N_14374);
and UO_1207 (O_1207,N_14339,N_14461);
nor UO_1208 (O_1208,N_14660,N_13792);
or UO_1209 (O_1209,N_13555,N_13544);
xor UO_1210 (O_1210,N_14352,N_13562);
and UO_1211 (O_1211,N_13920,N_13690);
and UO_1212 (O_1212,N_14373,N_14525);
or UO_1213 (O_1213,N_13954,N_14050);
and UO_1214 (O_1214,N_13727,N_13827);
nand UO_1215 (O_1215,N_14638,N_14702);
nand UO_1216 (O_1216,N_13989,N_13812);
and UO_1217 (O_1217,N_14732,N_13584);
and UO_1218 (O_1218,N_14812,N_13510);
or UO_1219 (O_1219,N_13809,N_14123);
xnor UO_1220 (O_1220,N_14549,N_13915);
nand UO_1221 (O_1221,N_13781,N_14604);
nor UO_1222 (O_1222,N_14835,N_14184);
nor UO_1223 (O_1223,N_13770,N_14057);
nor UO_1224 (O_1224,N_14100,N_14351);
or UO_1225 (O_1225,N_14456,N_14167);
nor UO_1226 (O_1226,N_14881,N_14897);
nand UO_1227 (O_1227,N_14695,N_13657);
xor UO_1228 (O_1228,N_13813,N_14097);
or UO_1229 (O_1229,N_14815,N_14081);
and UO_1230 (O_1230,N_14581,N_14154);
nor UO_1231 (O_1231,N_14110,N_13524);
nand UO_1232 (O_1232,N_14843,N_14190);
nor UO_1233 (O_1233,N_14236,N_14973);
nor UO_1234 (O_1234,N_13964,N_13591);
xnor UO_1235 (O_1235,N_14853,N_13591);
nand UO_1236 (O_1236,N_13611,N_14117);
nor UO_1237 (O_1237,N_14522,N_13978);
nand UO_1238 (O_1238,N_13608,N_13642);
and UO_1239 (O_1239,N_13589,N_14654);
nor UO_1240 (O_1240,N_14097,N_13782);
nand UO_1241 (O_1241,N_14598,N_13690);
and UO_1242 (O_1242,N_14024,N_14450);
and UO_1243 (O_1243,N_14020,N_13691);
nand UO_1244 (O_1244,N_14288,N_14533);
nand UO_1245 (O_1245,N_13807,N_13643);
or UO_1246 (O_1246,N_14927,N_14017);
or UO_1247 (O_1247,N_14158,N_14570);
and UO_1248 (O_1248,N_14606,N_14616);
nor UO_1249 (O_1249,N_14999,N_14036);
or UO_1250 (O_1250,N_14225,N_14834);
nand UO_1251 (O_1251,N_14133,N_13686);
nand UO_1252 (O_1252,N_14194,N_13542);
or UO_1253 (O_1253,N_14121,N_14844);
nand UO_1254 (O_1254,N_13792,N_14535);
xnor UO_1255 (O_1255,N_13872,N_14196);
and UO_1256 (O_1256,N_14966,N_13603);
nor UO_1257 (O_1257,N_14686,N_14656);
nor UO_1258 (O_1258,N_13802,N_14577);
nor UO_1259 (O_1259,N_13925,N_14385);
nand UO_1260 (O_1260,N_13876,N_14889);
nand UO_1261 (O_1261,N_14384,N_14117);
nor UO_1262 (O_1262,N_14776,N_14028);
and UO_1263 (O_1263,N_13746,N_14972);
nor UO_1264 (O_1264,N_14357,N_14851);
xnor UO_1265 (O_1265,N_13528,N_13983);
or UO_1266 (O_1266,N_14693,N_14950);
and UO_1267 (O_1267,N_14562,N_13656);
and UO_1268 (O_1268,N_13691,N_13781);
nand UO_1269 (O_1269,N_14400,N_14140);
nor UO_1270 (O_1270,N_14251,N_13839);
nand UO_1271 (O_1271,N_13521,N_14132);
nor UO_1272 (O_1272,N_14389,N_14189);
nand UO_1273 (O_1273,N_14674,N_14288);
nor UO_1274 (O_1274,N_13884,N_13987);
or UO_1275 (O_1275,N_14233,N_13623);
xnor UO_1276 (O_1276,N_13783,N_13665);
nand UO_1277 (O_1277,N_13650,N_14679);
nand UO_1278 (O_1278,N_14126,N_14924);
nor UO_1279 (O_1279,N_13855,N_13675);
or UO_1280 (O_1280,N_14253,N_13838);
or UO_1281 (O_1281,N_14330,N_14517);
nor UO_1282 (O_1282,N_13914,N_13568);
nor UO_1283 (O_1283,N_13673,N_14542);
and UO_1284 (O_1284,N_14812,N_14913);
nand UO_1285 (O_1285,N_13884,N_13928);
xor UO_1286 (O_1286,N_14186,N_14182);
or UO_1287 (O_1287,N_13796,N_14725);
and UO_1288 (O_1288,N_14335,N_14519);
or UO_1289 (O_1289,N_13910,N_14040);
or UO_1290 (O_1290,N_14987,N_14911);
and UO_1291 (O_1291,N_14239,N_14726);
nor UO_1292 (O_1292,N_14505,N_14243);
and UO_1293 (O_1293,N_14687,N_14846);
and UO_1294 (O_1294,N_13966,N_14553);
nand UO_1295 (O_1295,N_13997,N_13777);
and UO_1296 (O_1296,N_14822,N_14320);
and UO_1297 (O_1297,N_13566,N_14784);
or UO_1298 (O_1298,N_13805,N_13733);
or UO_1299 (O_1299,N_13502,N_13791);
nand UO_1300 (O_1300,N_14522,N_14258);
xor UO_1301 (O_1301,N_13757,N_14542);
and UO_1302 (O_1302,N_14027,N_14417);
xor UO_1303 (O_1303,N_13771,N_14013);
nor UO_1304 (O_1304,N_14925,N_14887);
nand UO_1305 (O_1305,N_14657,N_14309);
or UO_1306 (O_1306,N_14665,N_14657);
nor UO_1307 (O_1307,N_14869,N_14412);
nor UO_1308 (O_1308,N_14584,N_14976);
and UO_1309 (O_1309,N_14823,N_13778);
and UO_1310 (O_1310,N_14367,N_14602);
nand UO_1311 (O_1311,N_14149,N_14735);
and UO_1312 (O_1312,N_14963,N_13750);
or UO_1313 (O_1313,N_13885,N_14202);
and UO_1314 (O_1314,N_14483,N_14445);
nand UO_1315 (O_1315,N_14669,N_13501);
xnor UO_1316 (O_1316,N_14427,N_14426);
nor UO_1317 (O_1317,N_14098,N_13647);
nor UO_1318 (O_1318,N_14227,N_13570);
or UO_1319 (O_1319,N_13763,N_14289);
xnor UO_1320 (O_1320,N_14702,N_14946);
or UO_1321 (O_1321,N_14296,N_14872);
nor UO_1322 (O_1322,N_13998,N_14644);
or UO_1323 (O_1323,N_13606,N_14932);
and UO_1324 (O_1324,N_14412,N_14774);
nor UO_1325 (O_1325,N_14647,N_14576);
or UO_1326 (O_1326,N_13946,N_13885);
and UO_1327 (O_1327,N_13850,N_14544);
nor UO_1328 (O_1328,N_13540,N_13766);
and UO_1329 (O_1329,N_14215,N_14460);
nor UO_1330 (O_1330,N_14937,N_13877);
and UO_1331 (O_1331,N_13902,N_13731);
nand UO_1332 (O_1332,N_14966,N_13605);
nand UO_1333 (O_1333,N_14760,N_13546);
nor UO_1334 (O_1334,N_13872,N_14101);
and UO_1335 (O_1335,N_14338,N_13641);
or UO_1336 (O_1336,N_14475,N_14017);
nand UO_1337 (O_1337,N_13849,N_14334);
and UO_1338 (O_1338,N_13902,N_13881);
or UO_1339 (O_1339,N_13611,N_14892);
nand UO_1340 (O_1340,N_14671,N_14579);
xor UO_1341 (O_1341,N_13947,N_14648);
or UO_1342 (O_1342,N_14217,N_13582);
nand UO_1343 (O_1343,N_13951,N_14019);
xnor UO_1344 (O_1344,N_14011,N_13583);
nor UO_1345 (O_1345,N_14657,N_14266);
nand UO_1346 (O_1346,N_13988,N_14894);
or UO_1347 (O_1347,N_14436,N_14931);
nand UO_1348 (O_1348,N_13727,N_14378);
and UO_1349 (O_1349,N_14944,N_13978);
nand UO_1350 (O_1350,N_13813,N_14001);
and UO_1351 (O_1351,N_13636,N_14239);
nand UO_1352 (O_1352,N_14012,N_13763);
and UO_1353 (O_1353,N_14124,N_14627);
nand UO_1354 (O_1354,N_14364,N_14491);
and UO_1355 (O_1355,N_13706,N_14174);
and UO_1356 (O_1356,N_13997,N_14317);
and UO_1357 (O_1357,N_14217,N_13873);
nand UO_1358 (O_1358,N_13673,N_13808);
nand UO_1359 (O_1359,N_13731,N_14138);
or UO_1360 (O_1360,N_14943,N_14874);
and UO_1361 (O_1361,N_14990,N_13833);
and UO_1362 (O_1362,N_14759,N_14736);
nor UO_1363 (O_1363,N_13965,N_14753);
xnor UO_1364 (O_1364,N_14102,N_14974);
nand UO_1365 (O_1365,N_13646,N_14544);
and UO_1366 (O_1366,N_13917,N_14454);
or UO_1367 (O_1367,N_13729,N_14025);
nand UO_1368 (O_1368,N_13763,N_14117);
xor UO_1369 (O_1369,N_14795,N_14970);
nand UO_1370 (O_1370,N_13682,N_14044);
or UO_1371 (O_1371,N_14467,N_14230);
nand UO_1372 (O_1372,N_13731,N_13993);
nor UO_1373 (O_1373,N_13603,N_14180);
nand UO_1374 (O_1374,N_13947,N_13670);
nand UO_1375 (O_1375,N_14617,N_14648);
nand UO_1376 (O_1376,N_13576,N_13548);
or UO_1377 (O_1377,N_13856,N_14679);
nor UO_1378 (O_1378,N_13669,N_14790);
nand UO_1379 (O_1379,N_14047,N_14149);
nand UO_1380 (O_1380,N_13699,N_14424);
and UO_1381 (O_1381,N_14279,N_14110);
nor UO_1382 (O_1382,N_14421,N_13976);
nand UO_1383 (O_1383,N_14850,N_13969);
xor UO_1384 (O_1384,N_14517,N_14671);
xor UO_1385 (O_1385,N_13911,N_14438);
or UO_1386 (O_1386,N_14910,N_14987);
and UO_1387 (O_1387,N_14718,N_14735);
and UO_1388 (O_1388,N_13962,N_13589);
xnor UO_1389 (O_1389,N_13592,N_14683);
or UO_1390 (O_1390,N_14078,N_14825);
and UO_1391 (O_1391,N_14570,N_14393);
and UO_1392 (O_1392,N_14438,N_14204);
or UO_1393 (O_1393,N_13704,N_13803);
nor UO_1394 (O_1394,N_14792,N_14722);
nand UO_1395 (O_1395,N_14929,N_14759);
or UO_1396 (O_1396,N_14929,N_14605);
nand UO_1397 (O_1397,N_13905,N_14483);
nor UO_1398 (O_1398,N_14432,N_14146);
and UO_1399 (O_1399,N_14339,N_13766);
xnor UO_1400 (O_1400,N_14690,N_14598);
nand UO_1401 (O_1401,N_14535,N_14157);
nor UO_1402 (O_1402,N_14968,N_14682);
and UO_1403 (O_1403,N_13553,N_14796);
and UO_1404 (O_1404,N_13698,N_14973);
and UO_1405 (O_1405,N_14431,N_14458);
or UO_1406 (O_1406,N_13704,N_14919);
and UO_1407 (O_1407,N_13685,N_14021);
and UO_1408 (O_1408,N_14778,N_14901);
nor UO_1409 (O_1409,N_14700,N_14339);
xor UO_1410 (O_1410,N_13729,N_13560);
nand UO_1411 (O_1411,N_14565,N_13707);
and UO_1412 (O_1412,N_14652,N_13530);
and UO_1413 (O_1413,N_14729,N_13598);
nand UO_1414 (O_1414,N_14955,N_13906);
nor UO_1415 (O_1415,N_14800,N_14109);
or UO_1416 (O_1416,N_14911,N_14477);
xnor UO_1417 (O_1417,N_14804,N_14369);
nand UO_1418 (O_1418,N_14595,N_14637);
nor UO_1419 (O_1419,N_14755,N_14999);
nand UO_1420 (O_1420,N_14835,N_14654);
and UO_1421 (O_1421,N_14714,N_14246);
and UO_1422 (O_1422,N_14866,N_14326);
nor UO_1423 (O_1423,N_14386,N_14288);
or UO_1424 (O_1424,N_14877,N_14140);
nand UO_1425 (O_1425,N_13829,N_13711);
xor UO_1426 (O_1426,N_13764,N_14211);
nand UO_1427 (O_1427,N_14150,N_14247);
nor UO_1428 (O_1428,N_14678,N_14529);
or UO_1429 (O_1429,N_14634,N_14510);
and UO_1430 (O_1430,N_14794,N_14907);
xor UO_1431 (O_1431,N_13696,N_14852);
nand UO_1432 (O_1432,N_14172,N_13756);
xnor UO_1433 (O_1433,N_14927,N_14104);
and UO_1434 (O_1434,N_14146,N_14540);
and UO_1435 (O_1435,N_14854,N_14260);
and UO_1436 (O_1436,N_13840,N_13757);
nand UO_1437 (O_1437,N_13667,N_13661);
nand UO_1438 (O_1438,N_14692,N_13811);
or UO_1439 (O_1439,N_14993,N_13886);
and UO_1440 (O_1440,N_13835,N_14415);
nand UO_1441 (O_1441,N_13803,N_14116);
and UO_1442 (O_1442,N_13534,N_13803);
nand UO_1443 (O_1443,N_13644,N_14827);
or UO_1444 (O_1444,N_13653,N_14697);
or UO_1445 (O_1445,N_13947,N_14715);
or UO_1446 (O_1446,N_14843,N_14872);
nor UO_1447 (O_1447,N_14952,N_14646);
nand UO_1448 (O_1448,N_13537,N_13546);
xor UO_1449 (O_1449,N_13684,N_13599);
or UO_1450 (O_1450,N_14110,N_14115);
nand UO_1451 (O_1451,N_13534,N_13924);
nand UO_1452 (O_1452,N_14711,N_13973);
nor UO_1453 (O_1453,N_14741,N_13819);
xnor UO_1454 (O_1454,N_14038,N_14509);
and UO_1455 (O_1455,N_14876,N_14560);
and UO_1456 (O_1456,N_13556,N_14030);
nor UO_1457 (O_1457,N_13905,N_13638);
xnor UO_1458 (O_1458,N_14398,N_14631);
or UO_1459 (O_1459,N_13746,N_13564);
xor UO_1460 (O_1460,N_13865,N_14112);
nor UO_1461 (O_1461,N_14337,N_14473);
nor UO_1462 (O_1462,N_14696,N_14887);
nor UO_1463 (O_1463,N_14517,N_14851);
or UO_1464 (O_1464,N_14194,N_14968);
nand UO_1465 (O_1465,N_13573,N_13991);
or UO_1466 (O_1466,N_14619,N_13880);
and UO_1467 (O_1467,N_13955,N_14294);
or UO_1468 (O_1468,N_14849,N_14743);
nor UO_1469 (O_1469,N_14813,N_14416);
nor UO_1470 (O_1470,N_13710,N_14525);
and UO_1471 (O_1471,N_14262,N_13617);
nand UO_1472 (O_1472,N_13617,N_13792);
xnor UO_1473 (O_1473,N_13582,N_13694);
and UO_1474 (O_1474,N_13736,N_13913);
xnor UO_1475 (O_1475,N_13581,N_14102);
xor UO_1476 (O_1476,N_13992,N_14002);
nor UO_1477 (O_1477,N_14224,N_14930);
nand UO_1478 (O_1478,N_14805,N_13863);
and UO_1479 (O_1479,N_13996,N_13573);
nor UO_1480 (O_1480,N_14467,N_14416);
nor UO_1481 (O_1481,N_13762,N_14605);
and UO_1482 (O_1482,N_13845,N_13862);
nand UO_1483 (O_1483,N_14971,N_14357);
and UO_1484 (O_1484,N_13580,N_14968);
nor UO_1485 (O_1485,N_13930,N_13932);
and UO_1486 (O_1486,N_14523,N_13758);
and UO_1487 (O_1487,N_13735,N_13885);
nor UO_1488 (O_1488,N_13893,N_13896);
and UO_1489 (O_1489,N_14680,N_14878);
or UO_1490 (O_1490,N_14514,N_14340);
and UO_1491 (O_1491,N_13602,N_13866);
nand UO_1492 (O_1492,N_14034,N_14395);
and UO_1493 (O_1493,N_14033,N_14177);
and UO_1494 (O_1494,N_14489,N_14795);
and UO_1495 (O_1495,N_13688,N_14094);
and UO_1496 (O_1496,N_14216,N_14887);
or UO_1497 (O_1497,N_14199,N_13718);
and UO_1498 (O_1498,N_13974,N_14894);
xnor UO_1499 (O_1499,N_13736,N_14488);
nand UO_1500 (O_1500,N_14928,N_14528);
and UO_1501 (O_1501,N_14943,N_14395);
and UO_1502 (O_1502,N_13825,N_14563);
and UO_1503 (O_1503,N_13808,N_14528);
xor UO_1504 (O_1504,N_13744,N_14302);
and UO_1505 (O_1505,N_14929,N_13878);
xor UO_1506 (O_1506,N_13845,N_14760);
nor UO_1507 (O_1507,N_14965,N_13585);
nor UO_1508 (O_1508,N_14574,N_14152);
nand UO_1509 (O_1509,N_13705,N_14162);
nor UO_1510 (O_1510,N_14778,N_14260);
or UO_1511 (O_1511,N_14351,N_13644);
and UO_1512 (O_1512,N_14503,N_13639);
and UO_1513 (O_1513,N_13668,N_14775);
nand UO_1514 (O_1514,N_13725,N_13794);
nor UO_1515 (O_1515,N_13919,N_13679);
or UO_1516 (O_1516,N_14235,N_14596);
nor UO_1517 (O_1517,N_14651,N_13938);
or UO_1518 (O_1518,N_14004,N_13557);
and UO_1519 (O_1519,N_13652,N_14400);
or UO_1520 (O_1520,N_13797,N_14858);
or UO_1521 (O_1521,N_13728,N_13717);
or UO_1522 (O_1522,N_14716,N_13975);
nand UO_1523 (O_1523,N_14528,N_13860);
nor UO_1524 (O_1524,N_14037,N_14224);
nand UO_1525 (O_1525,N_14499,N_14719);
nand UO_1526 (O_1526,N_14971,N_14903);
nor UO_1527 (O_1527,N_14425,N_14291);
and UO_1528 (O_1528,N_14691,N_13729);
nor UO_1529 (O_1529,N_14837,N_14219);
nand UO_1530 (O_1530,N_14847,N_14823);
nand UO_1531 (O_1531,N_14175,N_13736);
or UO_1532 (O_1532,N_14439,N_14161);
and UO_1533 (O_1533,N_13703,N_13819);
and UO_1534 (O_1534,N_14958,N_13780);
or UO_1535 (O_1535,N_13945,N_14523);
nand UO_1536 (O_1536,N_14885,N_14572);
nand UO_1537 (O_1537,N_14502,N_14826);
nor UO_1538 (O_1538,N_13649,N_14499);
xnor UO_1539 (O_1539,N_14357,N_14849);
and UO_1540 (O_1540,N_14181,N_13890);
or UO_1541 (O_1541,N_14475,N_14574);
nor UO_1542 (O_1542,N_14242,N_14432);
xor UO_1543 (O_1543,N_13923,N_13799);
or UO_1544 (O_1544,N_14849,N_14909);
or UO_1545 (O_1545,N_13898,N_13895);
and UO_1546 (O_1546,N_14062,N_14907);
or UO_1547 (O_1547,N_13779,N_14842);
nor UO_1548 (O_1548,N_13554,N_13949);
and UO_1549 (O_1549,N_14608,N_13885);
or UO_1550 (O_1550,N_14251,N_14479);
and UO_1551 (O_1551,N_14569,N_13823);
nand UO_1552 (O_1552,N_14738,N_13893);
or UO_1553 (O_1553,N_14011,N_13508);
nor UO_1554 (O_1554,N_14317,N_14734);
nand UO_1555 (O_1555,N_14797,N_14538);
or UO_1556 (O_1556,N_14805,N_14243);
nor UO_1557 (O_1557,N_14423,N_13625);
nand UO_1558 (O_1558,N_14056,N_14900);
and UO_1559 (O_1559,N_14944,N_14433);
nor UO_1560 (O_1560,N_14883,N_13605);
or UO_1561 (O_1561,N_14222,N_14286);
or UO_1562 (O_1562,N_13653,N_14093);
nor UO_1563 (O_1563,N_13739,N_14096);
and UO_1564 (O_1564,N_14077,N_14625);
and UO_1565 (O_1565,N_14114,N_13636);
nor UO_1566 (O_1566,N_13981,N_13890);
nor UO_1567 (O_1567,N_13802,N_14323);
xor UO_1568 (O_1568,N_14924,N_14168);
and UO_1569 (O_1569,N_13538,N_13819);
xor UO_1570 (O_1570,N_14540,N_14350);
xnor UO_1571 (O_1571,N_13977,N_13773);
nor UO_1572 (O_1572,N_13504,N_13501);
nand UO_1573 (O_1573,N_13512,N_14711);
nor UO_1574 (O_1574,N_13746,N_14764);
nand UO_1575 (O_1575,N_14936,N_14267);
or UO_1576 (O_1576,N_14631,N_14551);
or UO_1577 (O_1577,N_14109,N_13928);
xnor UO_1578 (O_1578,N_13770,N_14218);
nor UO_1579 (O_1579,N_14836,N_14212);
nand UO_1580 (O_1580,N_13719,N_14213);
nand UO_1581 (O_1581,N_13547,N_13656);
xnor UO_1582 (O_1582,N_14007,N_13880);
nor UO_1583 (O_1583,N_14077,N_14744);
nand UO_1584 (O_1584,N_14008,N_13839);
and UO_1585 (O_1585,N_13640,N_14318);
and UO_1586 (O_1586,N_14733,N_14963);
nand UO_1587 (O_1587,N_14961,N_14721);
nand UO_1588 (O_1588,N_14819,N_14853);
or UO_1589 (O_1589,N_14599,N_14589);
and UO_1590 (O_1590,N_14995,N_14524);
xnor UO_1591 (O_1591,N_13596,N_14192);
or UO_1592 (O_1592,N_14806,N_14805);
nor UO_1593 (O_1593,N_13898,N_13693);
and UO_1594 (O_1594,N_14835,N_13913);
and UO_1595 (O_1595,N_14562,N_14507);
and UO_1596 (O_1596,N_14908,N_13589);
or UO_1597 (O_1597,N_14038,N_14684);
nor UO_1598 (O_1598,N_13599,N_14295);
or UO_1599 (O_1599,N_13560,N_14711);
or UO_1600 (O_1600,N_14954,N_14873);
or UO_1601 (O_1601,N_14567,N_14181);
nand UO_1602 (O_1602,N_14033,N_14845);
or UO_1603 (O_1603,N_14702,N_13653);
nor UO_1604 (O_1604,N_14311,N_14359);
or UO_1605 (O_1605,N_14494,N_14853);
xnor UO_1606 (O_1606,N_13722,N_14288);
and UO_1607 (O_1607,N_14601,N_14796);
xnor UO_1608 (O_1608,N_14208,N_13760);
or UO_1609 (O_1609,N_14827,N_14564);
nand UO_1610 (O_1610,N_14226,N_14675);
and UO_1611 (O_1611,N_13749,N_14264);
and UO_1612 (O_1612,N_14071,N_13618);
nor UO_1613 (O_1613,N_14231,N_14366);
xnor UO_1614 (O_1614,N_13610,N_13751);
nand UO_1615 (O_1615,N_13731,N_14487);
nand UO_1616 (O_1616,N_14822,N_14053);
and UO_1617 (O_1617,N_13999,N_13990);
nor UO_1618 (O_1618,N_14346,N_13982);
nor UO_1619 (O_1619,N_14843,N_13513);
xor UO_1620 (O_1620,N_14267,N_13541);
nand UO_1621 (O_1621,N_13748,N_14558);
nand UO_1622 (O_1622,N_14959,N_14078);
nand UO_1623 (O_1623,N_14414,N_14615);
nand UO_1624 (O_1624,N_13827,N_13734);
nor UO_1625 (O_1625,N_14576,N_14542);
nor UO_1626 (O_1626,N_14389,N_14023);
xnor UO_1627 (O_1627,N_13926,N_14963);
or UO_1628 (O_1628,N_14358,N_13791);
or UO_1629 (O_1629,N_13744,N_13932);
and UO_1630 (O_1630,N_13990,N_13931);
and UO_1631 (O_1631,N_14236,N_14566);
and UO_1632 (O_1632,N_14303,N_13926);
or UO_1633 (O_1633,N_13655,N_13788);
nor UO_1634 (O_1634,N_14441,N_14367);
nor UO_1635 (O_1635,N_14446,N_14495);
nor UO_1636 (O_1636,N_13982,N_14034);
or UO_1637 (O_1637,N_14513,N_14780);
xor UO_1638 (O_1638,N_13559,N_14011);
nor UO_1639 (O_1639,N_14085,N_13570);
xnor UO_1640 (O_1640,N_14285,N_13504);
nor UO_1641 (O_1641,N_13953,N_14476);
and UO_1642 (O_1642,N_13708,N_14303);
nand UO_1643 (O_1643,N_14209,N_13874);
or UO_1644 (O_1644,N_14704,N_13601);
and UO_1645 (O_1645,N_14117,N_13772);
xnor UO_1646 (O_1646,N_13674,N_13530);
nand UO_1647 (O_1647,N_14853,N_14972);
nor UO_1648 (O_1648,N_14521,N_13542);
and UO_1649 (O_1649,N_14217,N_14834);
and UO_1650 (O_1650,N_14401,N_13894);
or UO_1651 (O_1651,N_14717,N_14844);
and UO_1652 (O_1652,N_14619,N_13543);
or UO_1653 (O_1653,N_13705,N_14254);
nand UO_1654 (O_1654,N_14334,N_14549);
and UO_1655 (O_1655,N_14772,N_14738);
nand UO_1656 (O_1656,N_13894,N_14213);
or UO_1657 (O_1657,N_14383,N_13893);
and UO_1658 (O_1658,N_13825,N_13866);
and UO_1659 (O_1659,N_13819,N_14273);
or UO_1660 (O_1660,N_14708,N_14611);
nand UO_1661 (O_1661,N_14764,N_14625);
nand UO_1662 (O_1662,N_14195,N_14951);
and UO_1663 (O_1663,N_13747,N_14289);
and UO_1664 (O_1664,N_14624,N_14522);
nand UO_1665 (O_1665,N_13841,N_14594);
or UO_1666 (O_1666,N_14013,N_14711);
and UO_1667 (O_1667,N_14640,N_14688);
nor UO_1668 (O_1668,N_14409,N_13937);
or UO_1669 (O_1669,N_14026,N_13804);
xnor UO_1670 (O_1670,N_14235,N_14914);
xor UO_1671 (O_1671,N_14813,N_14303);
nor UO_1672 (O_1672,N_14224,N_14068);
and UO_1673 (O_1673,N_14038,N_13560);
nand UO_1674 (O_1674,N_14761,N_13779);
xor UO_1675 (O_1675,N_14800,N_13880);
and UO_1676 (O_1676,N_13937,N_14727);
nor UO_1677 (O_1677,N_13842,N_14360);
nand UO_1678 (O_1678,N_14090,N_14685);
xnor UO_1679 (O_1679,N_14402,N_13889);
and UO_1680 (O_1680,N_13878,N_14931);
nor UO_1681 (O_1681,N_14699,N_13967);
nor UO_1682 (O_1682,N_14494,N_14246);
xor UO_1683 (O_1683,N_13588,N_13595);
or UO_1684 (O_1684,N_14663,N_14931);
nor UO_1685 (O_1685,N_13941,N_14813);
and UO_1686 (O_1686,N_14668,N_13653);
nor UO_1687 (O_1687,N_13519,N_14155);
nand UO_1688 (O_1688,N_14971,N_13727);
xor UO_1689 (O_1689,N_14375,N_14069);
nand UO_1690 (O_1690,N_14223,N_14106);
nand UO_1691 (O_1691,N_14968,N_13659);
xnor UO_1692 (O_1692,N_14540,N_14536);
and UO_1693 (O_1693,N_14759,N_14909);
or UO_1694 (O_1694,N_14691,N_13589);
nor UO_1695 (O_1695,N_14868,N_14688);
nand UO_1696 (O_1696,N_13845,N_14944);
nand UO_1697 (O_1697,N_13883,N_14438);
or UO_1698 (O_1698,N_14252,N_13599);
xor UO_1699 (O_1699,N_14713,N_13794);
nand UO_1700 (O_1700,N_14152,N_13528);
xor UO_1701 (O_1701,N_14234,N_14601);
nor UO_1702 (O_1702,N_14221,N_14654);
nand UO_1703 (O_1703,N_14189,N_14208);
and UO_1704 (O_1704,N_14258,N_14808);
or UO_1705 (O_1705,N_14178,N_13591);
xnor UO_1706 (O_1706,N_13508,N_14726);
nor UO_1707 (O_1707,N_14131,N_14419);
or UO_1708 (O_1708,N_13885,N_13886);
xor UO_1709 (O_1709,N_14104,N_14299);
and UO_1710 (O_1710,N_14798,N_14942);
or UO_1711 (O_1711,N_14136,N_14075);
nor UO_1712 (O_1712,N_14632,N_14237);
xor UO_1713 (O_1713,N_13675,N_14632);
or UO_1714 (O_1714,N_14034,N_13917);
or UO_1715 (O_1715,N_14341,N_13893);
xor UO_1716 (O_1716,N_13856,N_13554);
nand UO_1717 (O_1717,N_14682,N_14565);
or UO_1718 (O_1718,N_14761,N_14840);
and UO_1719 (O_1719,N_14059,N_14565);
nor UO_1720 (O_1720,N_13518,N_14000);
and UO_1721 (O_1721,N_14737,N_13732);
nor UO_1722 (O_1722,N_14405,N_13642);
and UO_1723 (O_1723,N_14697,N_13754);
xor UO_1724 (O_1724,N_14052,N_13709);
or UO_1725 (O_1725,N_14006,N_14680);
nor UO_1726 (O_1726,N_13705,N_14902);
xnor UO_1727 (O_1727,N_14546,N_14025);
nor UO_1728 (O_1728,N_14106,N_14625);
nor UO_1729 (O_1729,N_14020,N_13926);
nor UO_1730 (O_1730,N_13995,N_14919);
nand UO_1731 (O_1731,N_13586,N_13851);
and UO_1732 (O_1732,N_14813,N_14251);
and UO_1733 (O_1733,N_14154,N_14861);
nand UO_1734 (O_1734,N_14304,N_14924);
nand UO_1735 (O_1735,N_14541,N_14730);
nor UO_1736 (O_1736,N_13509,N_14914);
or UO_1737 (O_1737,N_13941,N_13554);
and UO_1738 (O_1738,N_14655,N_14531);
nand UO_1739 (O_1739,N_13754,N_14710);
or UO_1740 (O_1740,N_13672,N_14213);
nor UO_1741 (O_1741,N_14671,N_14203);
or UO_1742 (O_1742,N_14658,N_14408);
nor UO_1743 (O_1743,N_14604,N_14917);
or UO_1744 (O_1744,N_13943,N_14462);
nor UO_1745 (O_1745,N_13758,N_14123);
nand UO_1746 (O_1746,N_13874,N_14322);
xor UO_1747 (O_1747,N_14261,N_14064);
nand UO_1748 (O_1748,N_14737,N_14816);
xnor UO_1749 (O_1749,N_14657,N_14158);
nor UO_1750 (O_1750,N_14066,N_14260);
nor UO_1751 (O_1751,N_14518,N_14288);
or UO_1752 (O_1752,N_14004,N_14266);
xnor UO_1753 (O_1753,N_13986,N_14058);
xor UO_1754 (O_1754,N_14818,N_14846);
nand UO_1755 (O_1755,N_13985,N_13762);
and UO_1756 (O_1756,N_13604,N_13681);
nand UO_1757 (O_1757,N_14646,N_13523);
nor UO_1758 (O_1758,N_14112,N_14313);
and UO_1759 (O_1759,N_14448,N_13753);
nor UO_1760 (O_1760,N_14695,N_14185);
or UO_1761 (O_1761,N_13597,N_14089);
or UO_1762 (O_1762,N_13935,N_14916);
nand UO_1763 (O_1763,N_14502,N_13614);
xnor UO_1764 (O_1764,N_13957,N_13948);
and UO_1765 (O_1765,N_13954,N_13615);
nand UO_1766 (O_1766,N_14689,N_14827);
and UO_1767 (O_1767,N_13870,N_14055);
and UO_1768 (O_1768,N_14908,N_14632);
or UO_1769 (O_1769,N_14794,N_13863);
and UO_1770 (O_1770,N_14751,N_13666);
or UO_1771 (O_1771,N_13821,N_14959);
xnor UO_1772 (O_1772,N_14853,N_14409);
nand UO_1773 (O_1773,N_14000,N_14076);
and UO_1774 (O_1774,N_14759,N_14602);
nor UO_1775 (O_1775,N_14170,N_14135);
nor UO_1776 (O_1776,N_14553,N_14959);
nand UO_1777 (O_1777,N_14685,N_14634);
and UO_1778 (O_1778,N_13870,N_14155);
nand UO_1779 (O_1779,N_14240,N_14716);
nand UO_1780 (O_1780,N_13609,N_13574);
and UO_1781 (O_1781,N_14587,N_13623);
nand UO_1782 (O_1782,N_14563,N_14205);
nand UO_1783 (O_1783,N_14585,N_14320);
nor UO_1784 (O_1784,N_14875,N_14269);
and UO_1785 (O_1785,N_14143,N_13847);
nor UO_1786 (O_1786,N_14888,N_13966);
nor UO_1787 (O_1787,N_14412,N_13964);
xor UO_1788 (O_1788,N_14633,N_14321);
or UO_1789 (O_1789,N_13795,N_13849);
or UO_1790 (O_1790,N_13634,N_14459);
and UO_1791 (O_1791,N_14464,N_14578);
nor UO_1792 (O_1792,N_14758,N_14083);
nand UO_1793 (O_1793,N_14793,N_14849);
and UO_1794 (O_1794,N_14156,N_14398);
xnor UO_1795 (O_1795,N_14238,N_14973);
nand UO_1796 (O_1796,N_14943,N_14668);
nor UO_1797 (O_1797,N_14154,N_14187);
and UO_1798 (O_1798,N_14841,N_13973);
nor UO_1799 (O_1799,N_13821,N_13602);
or UO_1800 (O_1800,N_14560,N_13683);
and UO_1801 (O_1801,N_14190,N_14171);
xnor UO_1802 (O_1802,N_13567,N_14187);
nand UO_1803 (O_1803,N_14660,N_13980);
nor UO_1804 (O_1804,N_14390,N_13527);
nor UO_1805 (O_1805,N_13856,N_13861);
and UO_1806 (O_1806,N_14760,N_14293);
nand UO_1807 (O_1807,N_14842,N_14674);
and UO_1808 (O_1808,N_14210,N_13516);
or UO_1809 (O_1809,N_13639,N_13531);
nor UO_1810 (O_1810,N_13503,N_14399);
nor UO_1811 (O_1811,N_13789,N_13879);
or UO_1812 (O_1812,N_14014,N_13975);
or UO_1813 (O_1813,N_14608,N_14707);
nand UO_1814 (O_1814,N_13773,N_14359);
and UO_1815 (O_1815,N_14009,N_14120);
nand UO_1816 (O_1816,N_14452,N_14830);
nand UO_1817 (O_1817,N_14246,N_14147);
nor UO_1818 (O_1818,N_14746,N_14854);
nand UO_1819 (O_1819,N_13827,N_13598);
nand UO_1820 (O_1820,N_14750,N_14388);
xor UO_1821 (O_1821,N_14133,N_14521);
nor UO_1822 (O_1822,N_13972,N_13997);
or UO_1823 (O_1823,N_13870,N_13893);
or UO_1824 (O_1824,N_13827,N_13796);
or UO_1825 (O_1825,N_14065,N_14771);
or UO_1826 (O_1826,N_13729,N_13578);
nand UO_1827 (O_1827,N_14595,N_14145);
or UO_1828 (O_1828,N_14269,N_13997);
or UO_1829 (O_1829,N_14787,N_13742);
nor UO_1830 (O_1830,N_14052,N_14970);
nor UO_1831 (O_1831,N_13861,N_14568);
xor UO_1832 (O_1832,N_13831,N_13730);
or UO_1833 (O_1833,N_13922,N_14096);
nand UO_1834 (O_1834,N_13629,N_13645);
xor UO_1835 (O_1835,N_14886,N_14003);
nor UO_1836 (O_1836,N_14426,N_13670);
nor UO_1837 (O_1837,N_14526,N_14096);
nand UO_1838 (O_1838,N_14498,N_13582);
xnor UO_1839 (O_1839,N_14240,N_14575);
nor UO_1840 (O_1840,N_14836,N_13522);
and UO_1841 (O_1841,N_14041,N_14066);
and UO_1842 (O_1842,N_14854,N_14618);
xnor UO_1843 (O_1843,N_13634,N_13732);
and UO_1844 (O_1844,N_13935,N_14203);
and UO_1845 (O_1845,N_14111,N_14676);
and UO_1846 (O_1846,N_13831,N_14899);
xnor UO_1847 (O_1847,N_14346,N_13791);
and UO_1848 (O_1848,N_13749,N_14434);
xnor UO_1849 (O_1849,N_14563,N_13704);
and UO_1850 (O_1850,N_14333,N_14162);
or UO_1851 (O_1851,N_14163,N_14007);
nor UO_1852 (O_1852,N_14572,N_13678);
and UO_1853 (O_1853,N_13916,N_13922);
nor UO_1854 (O_1854,N_14752,N_14776);
nand UO_1855 (O_1855,N_14238,N_13627);
or UO_1856 (O_1856,N_14220,N_14882);
and UO_1857 (O_1857,N_14031,N_14846);
nor UO_1858 (O_1858,N_14871,N_14044);
nor UO_1859 (O_1859,N_14184,N_14896);
and UO_1860 (O_1860,N_14392,N_14545);
and UO_1861 (O_1861,N_14536,N_13797);
nand UO_1862 (O_1862,N_14019,N_13526);
nand UO_1863 (O_1863,N_14947,N_14786);
or UO_1864 (O_1864,N_14571,N_14601);
or UO_1865 (O_1865,N_13521,N_13669);
nor UO_1866 (O_1866,N_14602,N_14084);
nand UO_1867 (O_1867,N_13723,N_14358);
or UO_1868 (O_1868,N_13853,N_13852);
nor UO_1869 (O_1869,N_14961,N_14230);
nand UO_1870 (O_1870,N_14483,N_13779);
nor UO_1871 (O_1871,N_14163,N_14282);
nor UO_1872 (O_1872,N_13627,N_14714);
nand UO_1873 (O_1873,N_14301,N_14219);
nor UO_1874 (O_1874,N_14519,N_13649);
and UO_1875 (O_1875,N_14893,N_14490);
nor UO_1876 (O_1876,N_14984,N_13720);
and UO_1877 (O_1877,N_14409,N_14570);
nand UO_1878 (O_1878,N_13899,N_13873);
nor UO_1879 (O_1879,N_14983,N_13738);
and UO_1880 (O_1880,N_14479,N_14093);
and UO_1881 (O_1881,N_14506,N_14110);
nand UO_1882 (O_1882,N_14465,N_13898);
and UO_1883 (O_1883,N_14543,N_13996);
or UO_1884 (O_1884,N_14727,N_13891);
or UO_1885 (O_1885,N_14237,N_14736);
nand UO_1886 (O_1886,N_14367,N_14292);
or UO_1887 (O_1887,N_14841,N_14872);
nor UO_1888 (O_1888,N_14733,N_13583);
xnor UO_1889 (O_1889,N_14495,N_13648);
nor UO_1890 (O_1890,N_14777,N_14588);
or UO_1891 (O_1891,N_14914,N_14734);
nor UO_1892 (O_1892,N_14901,N_13780);
nor UO_1893 (O_1893,N_14191,N_14879);
nand UO_1894 (O_1894,N_14722,N_13733);
or UO_1895 (O_1895,N_14973,N_13544);
nand UO_1896 (O_1896,N_14198,N_14638);
and UO_1897 (O_1897,N_14450,N_14726);
nor UO_1898 (O_1898,N_14227,N_14369);
or UO_1899 (O_1899,N_14243,N_14022);
nand UO_1900 (O_1900,N_13865,N_14848);
nor UO_1901 (O_1901,N_14794,N_13849);
nor UO_1902 (O_1902,N_13612,N_14382);
xor UO_1903 (O_1903,N_14329,N_13983);
or UO_1904 (O_1904,N_13655,N_14461);
nand UO_1905 (O_1905,N_14424,N_14623);
and UO_1906 (O_1906,N_14610,N_13745);
nor UO_1907 (O_1907,N_13510,N_14226);
or UO_1908 (O_1908,N_14240,N_14180);
nor UO_1909 (O_1909,N_14926,N_14582);
or UO_1910 (O_1910,N_14233,N_13799);
and UO_1911 (O_1911,N_14801,N_14798);
nand UO_1912 (O_1912,N_14912,N_14330);
nand UO_1913 (O_1913,N_14230,N_14577);
and UO_1914 (O_1914,N_14826,N_14561);
nor UO_1915 (O_1915,N_14877,N_14638);
nor UO_1916 (O_1916,N_13822,N_14334);
nand UO_1917 (O_1917,N_13710,N_14917);
nand UO_1918 (O_1918,N_14835,N_14849);
nand UO_1919 (O_1919,N_14359,N_14929);
xor UO_1920 (O_1920,N_14105,N_13687);
or UO_1921 (O_1921,N_13579,N_14265);
and UO_1922 (O_1922,N_13872,N_14923);
xnor UO_1923 (O_1923,N_14401,N_13740);
nor UO_1924 (O_1924,N_14134,N_14693);
nand UO_1925 (O_1925,N_13994,N_13837);
nand UO_1926 (O_1926,N_14148,N_14187);
xor UO_1927 (O_1927,N_13728,N_13744);
and UO_1928 (O_1928,N_13950,N_14669);
nor UO_1929 (O_1929,N_14312,N_13522);
nor UO_1930 (O_1930,N_13563,N_14517);
xnor UO_1931 (O_1931,N_13610,N_13518);
or UO_1932 (O_1932,N_13820,N_13714);
and UO_1933 (O_1933,N_14748,N_14314);
nor UO_1934 (O_1934,N_14800,N_14043);
or UO_1935 (O_1935,N_14622,N_14638);
xnor UO_1936 (O_1936,N_13572,N_14249);
and UO_1937 (O_1937,N_14423,N_13631);
or UO_1938 (O_1938,N_14198,N_13965);
nor UO_1939 (O_1939,N_13794,N_13859);
nand UO_1940 (O_1940,N_14760,N_14834);
and UO_1941 (O_1941,N_14089,N_14429);
and UO_1942 (O_1942,N_14047,N_14383);
or UO_1943 (O_1943,N_14335,N_14995);
and UO_1944 (O_1944,N_13672,N_13634);
xor UO_1945 (O_1945,N_14610,N_14304);
and UO_1946 (O_1946,N_13607,N_14838);
and UO_1947 (O_1947,N_13548,N_13724);
and UO_1948 (O_1948,N_13939,N_14093);
xor UO_1949 (O_1949,N_13990,N_13612);
and UO_1950 (O_1950,N_14794,N_13581);
nor UO_1951 (O_1951,N_14249,N_14686);
xor UO_1952 (O_1952,N_13780,N_14015);
nand UO_1953 (O_1953,N_13986,N_14184);
and UO_1954 (O_1954,N_13654,N_13853);
or UO_1955 (O_1955,N_13628,N_14743);
nor UO_1956 (O_1956,N_14778,N_14583);
and UO_1957 (O_1957,N_13807,N_13849);
nor UO_1958 (O_1958,N_13707,N_13866);
or UO_1959 (O_1959,N_14023,N_13535);
nor UO_1960 (O_1960,N_14785,N_13912);
xnor UO_1961 (O_1961,N_14477,N_14674);
and UO_1962 (O_1962,N_14347,N_14925);
nand UO_1963 (O_1963,N_14831,N_13782);
or UO_1964 (O_1964,N_13895,N_14166);
xor UO_1965 (O_1965,N_13550,N_14444);
nor UO_1966 (O_1966,N_13685,N_14652);
xor UO_1967 (O_1967,N_14401,N_14633);
and UO_1968 (O_1968,N_14790,N_13724);
or UO_1969 (O_1969,N_13645,N_14318);
xor UO_1970 (O_1970,N_14119,N_14088);
nand UO_1971 (O_1971,N_14082,N_14193);
nor UO_1972 (O_1972,N_14032,N_13882);
or UO_1973 (O_1973,N_14820,N_14613);
nor UO_1974 (O_1974,N_13624,N_13770);
nand UO_1975 (O_1975,N_14830,N_14998);
nand UO_1976 (O_1976,N_13726,N_13684);
nor UO_1977 (O_1977,N_14110,N_13659);
nor UO_1978 (O_1978,N_14228,N_13947);
xnor UO_1979 (O_1979,N_14419,N_14279);
or UO_1980 (O_1980,N_14287,N_14924);
nor UO_1981 (O_1981,N_14488,N_14158);
nand UO_1982 (O_1982,N_14071,N_13835);
nor UO_1983 (O_1983,N_13689,N_14523);
nand UO_1984 (O_1984,N_14559,N_14570);
or UO_1985 (O_1985,N_13687,N_14338);
nand UO_1986 (O_1986,N_14638,N_14864);
or UO_1987 (O_1987,N_14394,N_13531);
xor UO_1988 (O_1988,N_14340,N_14184);
and UO_1989 (O_1989,N_14422,N_14070);
nor UO_1990 (O_1990,N_13814,N_14104);
and UO_1991 (O_1991,N_13873,N_14631);
nor UO_1992 (O_1992,N_13758,N_14976);
nand UO_1993 (O_1993,N_13605,N_14863);
xnor UO_1994 (O_1994,N_14282,N_14353);
or UO_1995 (O_1995,N_14306,N_14524);
nor UO_1996 (O_1996,N_14829,N_14224);
and UO_1997 (O_1997,N_14515,N_14712);
nor UO_1998 (O_1998,N_14995,N_13567);
xnor UO_1999 (O_1999,N_13880,N_13995);
endmodule