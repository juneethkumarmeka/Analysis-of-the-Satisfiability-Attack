module basic_3000_30000_3500_100_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nor U0 (N_0,In_781,In_201);
nor U1 (N_1,In_1355,In_871);
nor U2 (N_2,In_890,In_2853);
and U3 (N_3,In_353,In_2123);
and U4 (N_4,In_2557,In_2074);
or U5 (N_5,In_468,In_753);
nand U6 (N_6,In_2717,In_2513);
nor U7 (N_7,In_959,In_2452);
xnor U8 (N_8,In_553,In_739);
and U9 (N_9,In_1906,In_2715);
and U10 (N_10,In_1196,In_84);
nand U11 (N_11,In_918,In_2460);
xnor U12 (N_12,In_2940,In_2810);
nand U13 (N_13,In_1835,In_2827);
nand U14 (N_14,In_760,In_2353);
nand U15 (N_15,In_1113,In_2366);
or U16 (N_16,In_926,In_1107);
nand U17 (N_17,In_2785,In_1216);
nand U18 (N_18,In_600,In_1825);
nand U19 (N_19,In_1000,In_2442);
and U20 (N_20,In_183,In_639);
or U21 (N_21,In_2328,In_378);
nand U22 (N_22,In_2743,In_1548);
or U23 (N_23,In_991,In_2739);
nor U24 (N_24,In_2484,In_822);
nand U25 (N_25,In_2969,In_1023);
and U26 (N_26,In_2536,In_908);
xnor U27 (N_27,In_2582,In_386);
or U28 (N_28,In_847,In_1086);
and U29 (N_29,In_2517,In_2677);
nand U30 (N_30,In_566,In_2134);
nand U31 (N_31,In_1637,In_1124);
xor U32 (N_32,In_2858,In_776);
xor U33 (N_33,In_2069,In_529);
or U34 (N_34,In_491,In_1406);
and U35 (N_35,In_1274,In_191);
xnor U36 (N_36,In_157,In_584);
xnor U37 (N_37,In_1927,In_2211);
nand U38 (N_38,In_669,In_1450);
nand U39 (N_39,In_2464,In_689);
nor U40 (N_40,In_2100,In_1270);
xnor U41 (N_41,In_2054,In_1775);
xnor U42 (N_42,In_924,In_2002);
nor U43 (N_43,In_696,In_2917);
nand U44 (N_44,In_608,In_2846);
and U45 (N_45,In_1440,In_1332);
nand U46 (N_46,In_1117,In_1601);
and U47 (N_47,In_87,In_1587);
and U48 (N_48,In_603,In_2222);
xor U49 (N_49,In_2908,In_454);
nor U50 (N_50,In_2400,In_121);
xnor U51 (N_51,In_2833,In_1719);
nand U52 (N_52,In_403,In_1593);
or U53 (N_53,In_1870,In_2560);
nand U54 (N_54,In_2662,In_1572);
nand U55 (N_55,In_2927,In_2550);
or U56 (N_56,In_86,In_658);
xnor U57 (N_57,In_2840,In_2558);
and U58 (N_58,In_619,In_1620);
xnor U59 (N_59,In_1946,In_376);
and U60 (N_60,In_686,In_740);
and U61 (N_61,In_1701,In_107);
nor U62 (N_62,In_176,In_2546);
or U63 (N_63,In_1389,In_2842);
xor U64 (N_64,In_1281,In_1191);
nand U65 (N_65,In_1673,In_1848);
nor U66 (N_66,In_2518,In_458);
nor U67 (N_67,In_2206,In_2479);
and U68 (N_68,In_1763,In_2773);
or U69 (N_69,In_1371,In_2961);
xor U70 (N_70,In_2880,In_2174);
nor U71 (N_71,In_2487,In_1517);
xor U72 (N_72,In_2352,In_2017);
nand U73 (N_73,In_902,In_1223);
and U74 (N_74,In_1001,In_2247);
and U75 (N_75,In_1081,In_1143);
and U76 (N_76,In_1592,In_481);
or U77 (N_77,In_1791,In_2294);
xor U78 (N_78,In_1758,In_1888);
xnor U79 (N_79,In_2433,In_2339);
xor U80 (N_80,In_2824,In_1509);
xor U81 (N_81,In_2989,In_2707);
nor U82 (N_82,In_1879,In_744);
and U83 (N_83,In_2208,In_1853);
xor U84 (N_84,In_2673,In_74);
xor U85 (N_85,In_2796,In_967);
or U86 (N_86,In_1268,In_2637);
nand U87 (N_87,In_2516,In_2543);
nor U88 (N_88,In_2616,In_1790);
nand U89 (N_89,In_718,In_361);
nand U90 (N_90,In_2886,In_2173);
or U91 (N_91,In_1602,In_104);
nor U92 (N_92,In_1305,In_35);
nand U93 (N_93,In_2732,In_1686);
or U94 (N_94,In_1662,In_2899);
or U95 (N_95,In_1063,In_866);
and U96 (N_96,In_1165,In_162);
nor U97 (N_97,In_2468,In_2344);
nand U98 (N_98,In_475,In_1512);
nand U99 (N_99,In_2018,In_1074);
or U100 (N_100,In_1530,In_2923);
nand U101 (N_101,In_1882,In_1590);
nand U102 (N_102,In_2085,In_1499);
and U103 (N_103,In_715,In_2008);
nor U104 (N_104,In_1626,In_1609);
nand U105 (N_105,In_793,In_25);
nor U106 (N_106,In_2434,In_1582);
nand U107 (N_107,In_670,In_1967);
xnor U108 (N_108,In_2248,In_2057);
and U109 (N_109,In_2843,In_1257);
or U110 (N_110,In_1142,In_1958);
nor U111 (N_111,In_2795,In_1994);
or U112 (N_112,In_466,In_2777);
and U113 (N_113,In_1072,In_752);
xnor U114 (N_114,In_1015,In_1319);
nor U115 (N_115,In_220,In_873);
nor U116 (N_116,In_592,In_938);
nor U117 (N_117,In_2430,In_936);
and U118 (N_118,In_1487,In_805);
nor U119 (N_119,In_2591,In_212);
nor U120 (N_120,In_2341,In_344);
nand U121 (N_121,In_1161,In_732);
xor U122 (N_122,In_268,In_775);
nor U123 (N_123,In_1738,In_1784);
nand U124 (N_124,In_802,In_1349);
nor U125 (N_125,In_1042,In_2976);
and U126 (N_126,In_1410,In_175);
nand U127 (N_127,In_2161,In_1523);
nor U128 (N_128,In_1412,In_2201);
nor U129 (N_129,In_562,In_645);
nand U130 (N_130,In_459,In_1394);
nor U131 (N_131,In_996,In_874);
or U132 (N_132,In_1811,In_1433);
xnor U133 (N_133,In_2348,In_569);
nor U134 (N_134,In_2738,In_1537);
and U135 (N_135,In_1698,In_390);
and U136 (N_136,In_1060,In_319);
xor U137 (N_137,In_1919,In_2242);
nor U138 (N_138,In_834,In_2067);
and U139 (N_139,In_618,In_13);
nand U140 (N_140,In_554,In_433);
nor U141 (N_141,In_1164,In_30);
nor U142 (N_142,In_1226,In_124);
and U143 (N_143,In_1114,In_714);
or U144 (N_144,In_722,In_1489);
nand U145 (N_145,In_197,In_666);
xnor U146 (N_146,In_248,In_1744);
nand U147 (N_147,In_2455,In_2727);
or U148 (N_148,In_214,In_2357);
xnor U149 (N_149,In_964,In_688);
nor U150 (N_150,In_1938,In_2236);
and U151 (N_151,In_2159,In_556);
or U152 (N_152,In_611,In_2481);
and U153 (N_153,In_245,In_1400);
nor U154 (N_154,In_602,In_1373);
nand U155 (N_155,In_1646,In_1043);
or U156 (N_156,In_1136,In_2572);
xor U157 (N_157,In_1195,In_2412);
or U158 (N_158,In_1631,In_1842);
or U159 (N_159,In_2102,In_1581);
xor U160 (N_160,In_637,In_1640);
nor U161 (N_161,In_1261,In_2011);
or U162 (N_162,In_1295,In_763);
nor U163 (N_163,In_1735,In_1426);
or U164 (N_164,In_422,In_2836);
xor U165 (N_165,In_2553,In_633);
and U166 (N_166,In_2866,In_2469);
and U167 (N_167,In_2802,In_416);
nor U168 (N_168,In_2830,In_494);
xnor U169 (N_169,In_2723,In_1491);
xor U170 (N_170,In_1108,In_2167);
nand U171 (N_171,In_2999,In_889);
or U172 (N_172,In_1183,In_995);
and U173 (N_173,In_517,In_1167);
or U174 (N_174,In_1265,In_1334);
nor U175 (N_175,In_2661,In_2408);
nor U176 (N_176,In_2522,In_2537);
xnor U177 (N_177,In_2774,In_1352);
nand U178 (N_178,In_1025,In_2407);
xor U179 (N_179,In_1773,In_1545);
or U180 (N_180,In_1013,In_2741);
or U181 (N_181,In_2091,In_2942);
xor U182 (N_182,In_396,In_1999);
nand U183 (N_183,In_661,In_853);
and U184 (N_184,In_406,In_1428);
and U185 (N_185,In_14,In_506);
xnor U186 (N_186,In_2768,In_258);
or U187 (N_187,In_755,In_2784);
xor U188 (N_188,In_1497,In_2718);
or U189 (N_189,In_356,In_1052);
nor U190 (N_190,In_146,In_143);
nor U191 (N_191,In_693,In_903);
nor U192 (N_192,In_557,In_2454);
or U193 (N_193,In_2992,In_1568);
xnor U194 (N_194,In_1316,In_1418);
nor U195 (N_195,In_1681,In_2960);
and U196 (N_196,In_572,In_1263);
nor U197 (N_197,In_892,In_698);
nor U198 (N_198,In_1665,In_2971);
xor U199 (N_199,In_2429,In_1365);
nor U200 (N_200,In_2640,In_765);
nand U201 (N_201,In_1241,In_2178);
xor U202 (N_202,In_424,In_180);
xnor U203 (N_203,In_1467,In_1213);
xnor U204 (N_204,In_2751,In_742);
nand U205 (N_205,In_646,In_2132);
and U206 (N_206,In_695,In_2444);
nand U207 (N_207,In_2139,In_904);
nor U208 (N_208,In_723,In_614);
nor U209 (N_209,In_72,In_2036);
or U210 (N_210,In_1127,In_23);
xor U211 (N_211,In_1617,In_2311);
nor U212 (N_212,In_2150,In_1901);
and U213 (N_213,In_2631,In_2221);
and U214 (N_214,In_128,In_333);
nand U215 (N_215,In_2828,In_2354);
or U216 (N_216,In_2890,In_2082);
or U217 (N_217,In_1722,In_2233);
nor U218 (N_218,In_2165,In_1580);
or U219 (N_219,In_109,In_2622);
xor U220 (N_220,In_4,In_257);
and U221 (N_221,In_1947,In_2577);
xnor U222 (N_222,In_660,In_2789);
and U223 (N_223,In_1903,In_563);
xor U224 (N_224,In_408,In_1873);
nor U225 (N_225,In_1745,In_982);
and U226 (N_226,In_502,In_624);
xor U227 (N_227,In_2531,In_304);
and U228 (N_228,In_2745,In_1885);
nand U229 (N_229,In_253,In_2656);
and U230 (N_230,In_2879,In_313);
nand U231 (N_231,In_2690,In_2682);
or U232 (N_232,In_894,In_2847);
xor U233 (N_233,In_1147,In_2919);
nand U234 (N_234,In_2657,In_1973);
xnor U235 (N_235,In_741,In_240);
or U236 (N_236,In_816,In_2169);
xor U237 (N_237,In_1469,In_1178);
or U238 (N_238,In_896,In_1514);
nand U239 (N_239,In_1621,In_218);
xnor U240 (N_240,In_1379,In_301);
xnor U241 (N_241,In_535,In_1623);
xnor U242 (N_242,In_1799,In_1900);
or U243 (N_243,In_298,In_2255);
or U244 (N_244,In_418,In_172);
or U245 (N_245,In_1669,In_2116);
and U246 (N_246,In_587,In_2146);
and U247 (N_247,In_1482,In_920);
nand U248 (N_248,In_2392,In_420);
nand U249 (N_249,In_1854,In_1571);
or U250 (N_250,In_1367,In_2826);
nand U251 (N_251,In_2972,In_708);
nand U252 (N_252,In_34,In_1920);
and U253 (N_253,In_2393,In_610);
or U254 (N_254,In_1207,In_2049);
or U255 (N_255,In_914,In_346);
xor U256 (N_256,In_125,In_2136);
nand U257 (N_257,In_1474,In_2514);
nor U258 (N_258,In_370,In_1106);
and U259 (N_259,In_225,In_2642);
and U260 (N_260,In_2483,In_311);
xor U261 (N_261,In_2540,In_574);
nand U262 (N_262,In_151,In_1085);
nor U263 (N_263,In_1310,In_2544);
or U264 (N_264,In_1990,In_374);
and U265 (N_265,In_2694,In_1886);
nand U266 (N_266,In_2816,In_2291);
xnor U267 (N_267,In_1579,In_2463);
nand U268 (N_268,In_2566,In_2959);
or U269 (N_269,In_260,In_546);
nor U270 (N_270,In_96,In_1012);
or U271 (N_271,In_1370,In_129);
xnor U272 (N_272,In_858,In_2901);
xnor U273 (N_273,In_2440,In_2417);
nand U274 (N_274,In_456,In_1109);
nand U275 (N_275,In_1359,In_1140);
nand U276 (N_276,In_1851,In_721);
nor U277 (N_277,In_812,In_2494);
or U278 (N_278,In_2027,In_2368);
nor U279 (N_279,In_397,In_483);
or U280 (N_280,In_2965,In_2046);
or U281 (N_281,In_919,In_1170);
and U282 (N_282,In_813,In_2697);
xor U283 (N_283,In_2274,In_2218);
and U284 (N_284,In_1283,In_208);
or U285 (N_285,In_532,In_206);
or U286 (N_286,In_1997,In_989);
nand U287 (N_287,In_2395,In_103);
and U288 (N_288,In_580,In_543);
xor U289 (N_289,In_2944,In_1566);
nor U290 (N_290,In_1133,In_2678);
and U291 (N_291,In_323,In_1856);
xor U292 (N_292,In_2099,In_1963);
and U293 (N_293,In_1859,In_1690);
xor U294 (N_294,In_1556,In_530);
or U295 (N_295,In_2439,In_1527);
xor U296 (N_296,In_426,In_2451);
nor U297 (N_297,In_2849,In_1761);
and U298 (N_298,In_943,In_1078);
or U299 (N_299,In_36,In_2115);
or U300 (N_300,In_2180,In_2421);
xnor U301 (N_301,In_2892,In_2336);
and U302 (N_302,In_2192,In_1276);
and U303 (N_303,In_2883,In_527);
and U304 (N_304,In_165,In_2384);
or U305 (N_305,N_46,In_2142);
and U306 (N_306,In_2051,In_1076);
or U307 (N_307,In_2109,In_193);
or U308 (N_308,In_1262,In_264);
nor U309 (N_309,In_949,In_2764);
and U310 (N_310,In_2474,In_1600);
or U311 (N_311,In_1457,In_2948);
and U312 (N_312,In_1102,In_1751);
nor U313 (N_313,In_878,In_2508);
nor U314 (N_314,N_260,In_250);
or U315 (N_315,In_1157,In_2427);
or U316 (N_316,In_879,In_1176);
or U317 (N_317,In_2725,In_237);
or U318 (N_318,In_2811,In_1361);
nor U319 (N_319,In_1717,In_1629);
and U320 (N_320,In_933,N_236);
and U321 (N_321,In_882,In_1059);
nand U322 (N_322,In_2576,In_2032);
xnor U323 (N_323,In_2962,In_1964);
and U324 (N_324,In_2356,N_259);
nor U325 (N_325,In_1695,In_2753);
nand U326 (N_326,In_152,In_2282);
nor U327 (N_327,In_1710,N_273);
xnor U328 (N_328,In_2106,In_1056);
nand U329 (N_329,In_2893,In_20);
nor U330 (N_330,In_2943,In_451);
nor U331 (N_331,In_792,In_728);
nor U332 (N_332,In_2997,In_2369);
nand U333 (N_333,In_1702,In_430);
xor U334 (N_334,In_2462,In_169);
nor U335 (N_335,In_1046,In_241);
xor U336 (N_336,In_280,In_2914);
nor U337 (N_337,In_687,In_368);
and U338 (N_338,In_1639,In_1050);
nand U339 (N_339,In_1041,In_203);
xor U340 (N_340,In_1477,In_2575);
and U341 (N_341,In_588,N_20);
nand U342 (N_342,In_1184,In_520);
nand U343 (N_343,In_667,In_1871);
xor U344 (N_344,In_2330,In_2335);
nor U345 (N_345,In_2580,In_1930);
or U346 (N_346,In_2070,In_1346);
and U347 (N_347,In_484,In_1655);
and U348 (N_348,In_2258,N_11);
or U349 (N_349,In_1335,In_1192);
xor U350 (N_350,N_6,In_1526);
and U351 (N_351,In_188,In_2787);
xnor U352 (N_352,In_1245,In_1360);
xor U353 (N_353,In_1622,In_2823);
xnor U354 (N_354,N_74,In_2612);
nor U355 (N_355,In_2014,In_1091);
nand U356 (N_356,In_992,In_1895);
or U357 (N_357,In_796,In_769);
and U358 (N_358,In_2670,In_1766);
and U359 (N_359,In_56,In_1887);
and U360 (N_360,In_1728,In_1700);
nor U361 (N_361,In_1510,In_2851);
nor U362 (N_362,In_1030,In_1553);
and U363 (N_363,In_2119,In_2559);
nor U364 (N_364,N_198,In_1080);
or U365 (N_365,In_762,In_2418);
or U366 (N_366,In_2175,In_1754);
or U367 (N_367,In_174,N_201);
and U368 (N_368,In_2910,N_166);
xnor U369 (N_369,In_2991,In_1126);
or U370 (N_370,In_2666,In_2658);
xnor U371 (N_371,In_1031,In_607);
and U372 (N_372,In_1857,In_1552);
xnor U373 (N_373,In_1541,In_2446);
nor U374 (N_374,In_2238,In_61);
nor U375 (N_375,In_2187,In_831);
and U376 (N_376,N_179,N_174);
xor U377 (N_377,In_1278,In_1405);
nor U378 (N_378,In_1670,In_1933);
and U379 (N_379,N_192,In_629);
and U380 (N_380,In_2592,In_2845);
nor U381 (N_381,In_1009,In_952);
xnor U382 (N_382,In_1716,In_1704);
nor U383 (N_383,In_6,In_1303);
and U384 (N_384,In_90,In_754);
xor U385 (N_385,N_266,In_998);
nand U386 (N_386,In_842,In_1275);
xor U387 (N_387,In_2272,In_2437);
or U388 (N_388,In_1808,In_962);
xor U389 (N_389,In_673,N_67);
nor U390 (N_390,In_1188,In_665);
nand U391 (N_391,In_821,In_1696);
nor U392 (N_392,In_419,In_635);
nand U393 (N_393,In_851,N_26);
xnor U394 (N_394,In_1255,In_10);
nand U395 (N_395,In_482,N_289);
and U396 (N_396,In_2689,In_1211);
and U397 (N_397,In_1792,In_163);
xnor U398 (N_398,In_1535,In_766);
nand U399 (N_399,In_2750,In_2915);
xnor U400 (N_400,In_1088,In_477);
and U401 (N_401,In_1819,In_707);
xnor U402 (N_402,In_1153,In_653);
nand U403 (N_403,In_1843,In_2549);
or U404 (N_404,In_2604,In_1366);
nor U405 (N_405,In_2327,In_318);
nand U406 (N_406,In_2438,In_1380);
nor U407 (N_407,In_473,In_2148);
and U408 (N_408,In_1219,In_683);
nand U409 (N_409,In_85,In_2138);
and U410 (N_410,In_380,In_100);
or U411 (N_411,In_2981,In_89);
or U412 (N_412,In_2402,In_1569);
nand U413 (N_413,In_1180,N_224);
and U414 (N_414,In_761,In_1232);
or U415 (N_415,N_3,N_292);
and U416 (N_416,N_293,In_1082);
xnor U417 (N_417,In_97,In_1777);
and U418 (N_418,In_78,In_1197);
nand U419 (N_419,In_2194,In_694);
nor U420 (N_420,In_1402,N_111);
and U421 (N_421,In_692,In_1902);
nor U422 (N_422,In_1508,In_1960);
nor U423 (N_423,In_1026,In_2435);
nand U424 (N_424,N_90,In_1331);
nor U425 (N_425,In_2918,In_2834);
nand U426 (N_426,In_1989,In_1287);
nor U427 (N_427,N_253,In_797);
or U428 (N_428,In_28,In_1048);
nand U429 (N_429,In_1976,In_2020);
nor U430 (N_430,In_2263,In_616);
or U431 (N_431,In_156,In_2312);
or U432 (N_432,In_888,In_2094);
and U433 (N_433,In_432,N_167);
nor U434 (N_434,In_2310,In_1653);
and U435 (N_435,In_2308,In_2377);
or U436 (N_436,In_647,In_1326);
nand U437 (N_437,In_917,In_411);
or U438 (N_438,In_631,In_1090);
xor U439 (N_439,In_0,In_2770);
nand U440 (N_440,N_221,In_1844);
or U441 (N_441,In_644,In_355);
nor U442 (N_442,In_2414,In_863);
xnor U443 (N_443,In_922,In_1028);
xor U444 (N_444,N_156,In_147);
nor U445 (N_445,In_2984,In_428);
nand U446 (N_446,In_2696,In_2583);
and U447 (N_447,In_93,In_1543);
nand U448 (N_448,In_2854,N_222);
nor U449 (N_449,In_1229,In_1576);
or U450 (N_450,In_305,In_1236);
nand U451 (N_451,In_1908,N_269);
and U452 (N_452,In_2620,In_861);
nor U453 (N_453,In_2567,In_2246);
nor U454 (N_454,In_1228,In_657);
or U455 (N_455,In_155,In_895);
xor U456 (N_456,In_1193,In_293);
xor U457 (N_457,In_2135,In_2144);
nor U458 (N_458,In_1064,In_2602);
nand U459 (N_459,In_2664,In_492);
and U460 (N_460,In_724,In_1551);
and U461 (N_461,In_860,In_210);
xnor U462 (N_462,In_2737,In_2736);
and U463 (N_463,In_1692,In_839);
xnor U464 (N_464,In_2952,In_1813);
or U465 (N_465,In_713,N_76);
nor U466 (N_466,In_815,In_231);
nand U467 (N_467,In_794,In_1540);
and U468 (N_468,In_1309,In_1838);
nor U469 (N_469,In_2005,N_91);
or U470 (N_470,In_1520,In_2683);
nand U471 (N_471,In_2062,In_1171);
and U472 (N_472,In_827,In_1847);
or U473 (N_473,In_897,In_1691);
and U474 (N_474,N_54,In_1417);
or U475 (N_475,N_53,In_2103);
nand U476 (N_476,In_2470,N_33);
xor U477 (N_477,In_2378,In_643);
xnor U478 (N_478,In_699,N_104);
nor U479 (N_479,N_83,In_440);
or U480 (N_480,In_613,In_538);
nand U481 (N_481,In_196,In_1019);
nand U482 (N_482,In_1430,In_2362);
xor U483 (N_483,In_1269,In_771);
xnor U484 (N_484,In_1354,In_2756);
or U485 (N_485,In_2023,In_1159);
nand U486 (N_486,In_940,In_443);
and U487 (N_487,In_2275,N_187);
xor U488 (N_488,In_2269,N_160);
nand U489 (N_489,In_1444,In_1242);
or U490 (N_490,In_488,In_476);
or U491 (N_491,In_2698,In_434);
xor U492 (N_492,In_737,In_944);
or U493 (N_493,In_1011,In_2818);
or U494 (N_494,In_568,In_2154);
and U495 (N_495,In_1397,N_249);
nor U496 (N_496,In_640,In_2276);
nor U497 (N_497,In_1125,N_113);
xor U498 (N_498,In_749,In_68);
xor U499 (N_499,In_2290,In_1614);
or U500 (N_500,In_111,In_465);
nor U501 (N_501,In_2829,In_654);
and U502 (N_502,In_2087,In_2542);
and U503 (N_503,In_656,N_161);
nand U504 (N_504,In_2261,In_1585);
xor U505 (N_505,In_736,N_213);
xor U506 (N_506,N_130,In_2848);
xor U507 (N_507,In_2510,In_1473);
nor U508 (N_508,In_1787,In_1243);
xor U509 (N_509,In_69,In_2945);
and U510 (N_510,In_2241,In_2045);
xnor U511 (N_511,In_2855,In_168);
xnor U512 (N_512,In_528,In_807);
xnor U513 (N_513,In_1720,In_676);
and U514 (N_514,In_400,In_1531);
or U515 (N_515,In_778,In_734);
nand U516 (N_516,In_2988,In_1588);
and U517 (N_517,In_2552,In_1876);
or U518 (N_518,In_2808,In_1279);
nand U519 (N_519,In_1066,In_678);
or U520 (N_520,In_758,In_2108);
nand U521 (N_521,In_1969,In_2405);
nand U522 (N_522,In_425,In_1478);
nor U523 (N_523,In_2935,In_638);
or U524 (N_524,In_636,N_212);
nor U525 (N_525,In_965,In_2713);
nor U526 (N_526,In_2098,In_2782);
nor U527 (N_527,In_1929,In_1432);
nor U528 (N_528,In_2679,In_1603);
nor U529 (N_529,In_1010,N_219);
nor U530 (N_530,N_239,In_1105);
nand U531 (N_531,In_2215,In_891);
or U532 (N_532,In_598,In_1141);
or U533 (N_533,In_1658,In_358);
and U534 (N_534,N_60,In_1247);
and U535 (N_535,N_136,In_2486);
nor U536 (N_536,In_2156,In_2963);
or U537 (N_537,In_1935,In_2447);
xnor U538 (N_538,In_2244,N_112);
xnor U539 (N_539,In_265,In_2381);
nand U540 (N_540,In_2556,In_2033);
nor U541 (N_541,In_2964,In_837);
and U542 (N_542,In_1534,In_1968);
or U543 (N_543,In_1996,In_91);
nor U544 (N_544,In_2922,In_544);
and U545 (N_545,N_153,In_1324);
and U546 (N_546,In_79,In_1706);
and U547 (N_547,In_1893,N_120);
xor U548 (N_548,In_178,In_1393);
nor U549 (N_549,In_1476,In_961);
and U550 (N_550,In_1409,In_1353);
or U551 (N_551,In_2224,In_2031);
nand U552 (N_552,In_1864,In_2325);
or U553 (N_553,In_259,In_179);
or U554 (N_554,In_2500,N_251);
nor U555 (N_555,In_738,In_1427);
nor U556 (N_556,In_585,In_2204);
and U557 (N_557,In_1437,In_1944);
xor U558 (N_558,N_135,In_1411);
xor U559 (N_559,In_1982,In_1767);
nand U560 (N_560,N_243,In_1699);
or U561 (N_561,In_2632,In_398);
and U562 (N_562,In_1413,In_1490);
or U563 (N_563,In_486,In_452);
nand U564 (N_564,In_3,In_2355);
and U565 (N_565,In_2515,In_2776);
nor U566 (N_566,In_659,In_876);
nor U567 (N_567,In_2004,In_2097);
xor U568 (N_568,In_1387,In_1089);
nor U569 (N_569,In_2279,In_1805);
nand U570 (N_570,In_2239,N_237);
xor U571 (N_571,In_2473,In_1659);
nand U572 (N_572,In_267,In_1231);
nor U573 (N_573,In_2509,In_209);
and U574 (N_574,In_446,In_76);
nand U575 (N_575,In_1244,In_2111);
nor U576 (N_576,In_1925,In_2596);
xnor U577 (N_577,In_1459,In_509);
nand U578 (N_578,In_1583,In_2183);
nor U579 (N_579,In_541,In_2681);
nor U580 (N_580,In_2699,In_2535);
nand U581 (N_581,In_2404,In_1746);
nand U582 (N_582,In_1796,N_284);
nand U583 (N_583,In_2000,In_1495);
or U584 (N_584,In_1458,In_1561);
xnor U585 (N_585,In_2920,In_2264);
and U586 (N_586,In_1014,In_1965);
nor U587 (N_587,In_263,In_1338);
nor U588 (N_588,In_980,In_1649);
nand U589 (N_589,In_1977,In_1118);
or U590 (N_590,In_120,N_286);
xnor U591 (N_591,N_124,In_278);
and U592 (N_592,In_364,In_1212);
xnor U593 (N_593,In_829,N_268);
nor U594 (N_594,In_521,In_561);
and U595 (N_595,In_1194,In_1119);
and U596 (N_596,In_1896,In_1252);
or U597 (N_597,In_559,In_153);
nand U598 (N_598,In_501,In_1521);
xor U599 (N_599,In_18,In_1970);
or U600 (N_600,In_1618,N_416);
nand U601 (N_601,In_2300,In_972);
xnor U602 (N_602,In_921,In_297);
xor U603 (N_603,In_2386,In_2155);
and U604 (N_604,In_573,In_2973);
or U605 (N_605,In_1376,In_930);
and U606 (N_606,In_2076,N_359);
nor U607 (N_607,N_207,In_2498);
nand U608 (N_608,N_315,In_2996);
and U609 (N_609,In_2374,N_461);
xnor U610 (N_610,N_1,In_194);
nor U611 (N_611,In_700,In_2902);
nor U612 (N_612,In_768,N_87);
and U613 (N_613,In_746,N_48);
and U614 (N_614,In_2547,In_1372);
or U615 (N_615,In_1884,In_384);
nor U616 (N_616,In_2379,N_186);
xor U617 (N_617,In_2013,In_1115);
xor U618 (N_618,N_12,N_155);
and U619 (N_619,N_142,In_2329);
nand U620 (N_620,N_431,In_2184);
nand U621 (N_621,In_974,In_2299);
nor U622 (N_622,N_152,In_5);
nand U623 (N_623,In_190,In_1455);
nor U624 (N_624,In_854,In_859);
and U625 (N_625,In_2872,In_388);
xnor U626 (N_626,In_63,In_429);
and U627 (N_627,In_2709,In_224);
xnor U628 (N_628,In_73,In_472);
and U629 (N_629,N_473,N_463);
nand U630 (N_630,N_449,In_1092);
nand U631 (N_631,N_519,In_1800);
nand U632 (N_632,N_573,In_1827);
nand U633 (N_633,In_2450,In_375);
xnor U634 (N_634,In_2804,In_885);
or U635 (N_635,In_1821,In_289);
or U636 (N_636,In_2614,In_2456);
nor U637 (N_637,In_1802,In_2083);
nand U638 (N_638,In_463,In_1454);
and U639 (N_639,In_2249,In_565);
xnor U640 (N_640,N_478,In_232);
nor U641 (N_641,In_2929,In_2747);
nand U642 (N_642,In_328,In_2316);
xor U643 (N_643,In_560,In_92);
xnor U644 (N_644,In_1038,N_533);
or U645 (N_645,In_322,In_671);
nor U646 (N_646,In_77,N_590);
and U647 (N_647,In_1209,N_240);
nand U648 (N_648,In_251,In_2692);
nor U649 (N_649,In_1726,In_1936);
or U650 (N_650,N_410,In_1916);
nor U651 (N_651,In_531,In_1542);
or U652 (N_652,In_801,N_23);
and U653 (N_653,N_528,In_1516);
and U654 (N_654,In_2871,In_236);
xnor U655 (N_655,N_429,In_2629);
nand U656 (N_656,In_2317,In_2792);
or U657 (N_657,In_2086,In_2528);
nand U658 (N_658,N_27,In_2101);
xnor U659 (N_659,In_335,In_2597);
and U660 (N_660,N_390,In_625);
nand U661 (N_661,In_2571,N_388);
and U662 (N_662,In_469,In_2593);
nand U663 (N_663,In_2058,In_1611);
nand U664 (N_664,N_394,In_2080);
nor U665 (N_665,In_756,In_1251);
and U666 (N_666,In_1364,In_16);
nand U667 (N_667,N_574,In_1032);
xor U668 (N_668,In_2198,In_757);
xnor U669 (N_669,In_2906,In_2037);
xor U670 (N_670,In_2432,In_1308);
or U671 (N_671,In_1718,In_2283);
nor U672 (N_672,N_481,N_149);
xnor U673 (N_673,In_1672,In_453);
or U674 (N_674,In_132,In_2225);
nand U675 (N_675,In_1154,In_1830);
or U676 (N_676,In_1320,In_2769);
and U677 (N_677,In_1714,In_2523);
xnor U678 (N_678,In_247,N_115);
nand U679 (N_679,In_2122,N_535);
or U680 (N_680,In_987,In_748);
or U681 (N_681,In_2060,N_176);
and U682 (N_682,In_880,In_2254);
xor U683 (N_683,In_1139,In_729);
or U684 (N_684,In_2193,In_275);
nand U685 (N_685,In_772,In_537);
nor U686 (N_686,N_329,In_1388);
xnor U687 (N_687,In_2061,In_825);
and U688 (N_688,In_1904,N_556);
xor U689 (N_689,In_391,In_2232);
nand U690 (N_690,N_35,In_2394);
xnor U691 (N_691,In_150,In_1912);
or U692 (N_692,In_909,In_2599);
nand U693 (N_693,N_474,In_2877);
nand U694 (N_694,N_370,In_2889);
xnor U695 (N_695,In_2941,In_1172);
xnor U696 (N_696,N_172,In_83);
nor U697 (N_697,In_2130,N_68);
nor U698 (N_698,N_417,In_261);
or U699 (N_699,In_1452,In_2501);
nor U700 (N_700,In_988,N_158);
xor U701 (N_701,In_571,N_72);
nor U702 (N_702,In_2653,N_325);
or U703 (N_703,In_1330,N_21);
nand U704 (N_704,In_2554,In_2655);
nor U705 (N_705,N_50,In_2321);
and U706 (N_706,In_2708,In_1222);
or U707 (N_707,N_13,In_254);
xor U708 (N_708,In_1407,In_1984);
and U709 (N_709,N_313,In_421);
or U710 (N_710,In_1987,N_570);
or U711 (N_711,In_2197,In_840);
nor U712 (N_712,In_609,In_1301);
and U713 (N_713,N_215,N_314);
nand U714 (N_714,In_1134,In_1748);
nand U715 (N_715,N_317,In_782);
or U716 (N_716,In_1221,N_312);
nand U717 (N_717,In_612,In_862);
nand U718 (N_718,In_731,In_1798);
xor U719 (N_719,In_1166,N_458);
xnor U720 (N_720,In_788,N_209);
nor U721 (N_721,In_957,In_1234);
nand U722 (N_722,In_2798,In_285);
xnor U723 (N_723,In_2788,In_1384);
nor U724 (N_724,In_593,In_2617);
nand U725 (N_725,In_1343,In_710);
nand U726 (N_726,In_1855,In_522);
nand U727 (N_727,In_2608,In_2372);
and U728 (N_728,In_229,In_994);
or U729 (N_729,In_819,In_2035);
or U730 (N_730,In_1158,In_1539);
nor U731 (N_731,In_401,N_568);
xor U732 (N_732,N_14,N_119);
nand U733 (N_733,In_586,In_2284);
or U734 (N_734,In_1959,In_2831);
and U735 (N_735,In_1280,In_2758);
nand U736 (N_736,In_342,In_2589);
and U737 (N_737,In_779,In_1045);
xnor U738 (N_738,In_33,N_361);
nor U739 (N_739,In_1980,In_1667);
or U740 (N_740,In_2805,In_2985);
xor U741 (N_741,In_664,In_963);
nor U742 (N_742,In_2921,N_483);
nor U743 (N_743,In_1550,In_705);
or U744 (N_744,N_294,N_513);
and U745 (N_745,N_285,N_382);
and U746 (N_746,N_92,In_2105);
nand U747 (N_747,In_1190,In_2323);
or U748 (N_748,In_490,In_2007);
nand U749 (N_749,In_551,In_620);
or U750 (N_750,In_2579,In_2493);
and U751 (N_751,In_906,In_2268);
nor U752 (N_752,N_238,In_1456);
nor U753 (N_753,In_1679,N_118);
nor U754 (N_754,In_227,In_2701);
and U755 (N_755,In_2297,In_2693);
nor U756 (N_756,In_1121,N_377);
and U757 (N_757,In_2635,N_436);
nor U758 (N_758,In_1267,N_495);
xnor U759 (N_759,In_2093,In_867);
and U760 (N_760,N_541,In_634);
and U761 (N_761,In_1797,In_798);
and U762 (N_762,In_1922,N_502);
or U763 (N_763,N_101,N_7);
xnor U764 (N_764,In_510,In_550);
or U765 (N_765,N_256,N_450);
nor U766 (N_766,In_2044,In_1058);
and U767 (N_767,In_362,N_177);
and U768 (N_768,N_395,In_1163);
nor U769 (N_769,N_122,In_1564);
or U770 (N_770,N_415,N_501);
nand U771 (N_771,In_941,In_1823);
nor U772 (N_772,In_711,In_2118);
and U773 (N_773,In_493,In_1494);
nand U774 (N_774,In_1524,In_836);
nor U775 (N_775,In_1554,In_703);
and U776 (N_776,N_392,In_244);
nand U777 (N_777,N_228,In_2641);
and U778 (N_778,In_1307,In_727);
or U779 (N_779,N_279,In_399);
or U780 (N_780,In_1345,In_848);
nor U781 (N_781,In_1322,In_2507);
xor U782 (N_782,N_323,In_627);
nand U783 (N_783,In_720,In_2491);
and U784 (N_784,In_2170,In_1177);
xnor U785 (N_785,In_2595,N_169);
or U786 (N_786,In_1486,N_109);
nand U787 (N_787,In_2755,N_216);
or U788 (N_788,In_1961,N_99);
xnor U789 (N_789,In_211,N_116);
or U790 (N_790,N_426,In_461);
or U791 (N_791,In_205,N_71);
and U792 (N_792,In_295,N_456);
and U793 (N_793,N_252,N_599);
nor U794 (N_794,In_2548,In_395);
nand U795 (N_795,In_1914,N_143);
and U796 (N_796,N_197,In_2133);
nor U797 (N_797,In_507,In_856);
nand U798 (N_798,In_29,In_1803);
xnor U799 (N_799,N_376,N_241);
and U800 (N_800,In_2199,In_817);
xnor U801 (N_801,In_1567,In_2562);
and U802 (N_802,In_1570,In_795);
nor U803 (N_803,In_44,In_946);
or U804 (N_804,In_485,In_101);
nor U805 (N_805,In_2112,In_1225);
and U806 (N_806,In_2129,In_784);
xnor U807 (N_807,In_1037,In_2286);
nand U808 (N_808,In_852,In_449);
nand U809 (N_809,In_2320,In_2767);
or U810 (N_810,In_605,N_522);
nand U811 (N_811,In_2485,In_2096);
nor U812 (N_812,In_1874,In_1503);
nand U813 (N_813,In_2809,In_2685);
and U814 (N_814,In_1463,In_595);
nand U815 (N_815,In_1753,N_345);
or U816 (N_816,In_2684,In_2025);
or U817 (N_817,In_1755,N_15);
nand U818 (N_818,In_1021,In_2399);
and U819 (N_819,In_1676,In_628);
and U820 (N_820,In_910,In_1129);
xor U821 (N_821,In_1863,In_2820);
and U822 (N_822,In_2630,In_339);
or U823 (N_823,N_397,N_138);
nor U824 (N_824,In_2410,N_425);
and U825 (N_825,N_248,In_2164);
xnor U826 (N_826,N_56,In_2065);
nor U827 (N_827,In_1390,In_148);
xnor U828 (N_828,N_98,N_499);
or U829 (N_829,N_185,In_2638);
or U830 (N_830,In_1525,In_1708);
nor U831 (N_831,In_662,In_372);
and U832 (N_832,In_315,In_747);
nor U833 (N_833,In_1067,In_2763);
or U834 (N_834,In_2628,In_2024);
nor U835 (N_835,In_1652,In_309);
or U836 (N_836,N_355,N_331);
nor U837 (N_837,In_1327,In_2465);
nand U838 (N_838,N_446,In_1546);
xnor U839 (N_839,N_438,N_512);
and U840 (N_840,In_1382,In_58);
and U841 (N_841,In_2887,N_396);
and U842 (N_842,In_1022,In_15);
or U843 (N_843,In_2760,In_1235);
xnor U844 (N_844,In_1498,In_651);
or U845 (N_845,In_1678,In_2039);
nand U846 (N_846,In_1101,N_421);
xor U847 (N_847,In_2607,In_2686);
or U848 (N_848,In_1734,In_726);
nor U849 (N_849,N_400,In_2147);
nand U850 (N_850,In_2613,In_1992);
xor U851 (N_851,In_1983,In_1804);
nand U852 (N_852,In_685,In_2322);
nor U853 (N_853,In_937,In_2530);
or U854 (N_854,In_2235,In_1029);
or U855 (N_855,In_135,In_913);
or U856 (N_856,In_2358,In_1318);
xnor U857 (N_857,In_596,N_347);
and U858 (N_858,In_1016,N_350);
or U859 (N_859,In_1302,In_877);
and U860 (N_860,In_1599,In_2600);
and U861 (N_861,In_272,N_36);
or U862 (N_862,In_1713,In_898);
and U863 (N_863,N_229,In_1425);
and U864 (N_864,In_1869,In_286);
nand U865 (N_865,In_680,In_450);
or U866 (N_866,In_2262,In_2151);
nand U867 (N_867,In_1664,In_1404);
and U868 (N_868,In_1339,In_1120);
xor U869 (N_869,In_2243,In_2957);
and U870 (N_870,In_2852,In_1991);
xor U871 (N_871,In_2946,In_2525);
or U872 (N_872,In_1416,N_183);
nor U873 (N_873,In_2229,In_288);
xnor U874 (N_874,In_2928,In_1277);
or U875 (N_875,In_2633,In_2042);
nor U876 (N_876,In_2574,In_2288);
and U877 (N_877,N_509,N_173);
nand U878 (N_878,In_1807,N_47);
nand U879 (N_879,In_2975,In_71);
nor U880 (N_880,In_2359,In_589);
nand U881 (N_881,N_582,In_479);
nand U882 (N_882,In_1071,In_2293);
or U883 (N_883,In_427,In_1506);
nand U884 (N_884,In_2048,In_1687);
and U885 (N_885,In_2223,In_1750);
and U886 (N_886,In_2207,In_2598);
nand U887 (N_887,In_1891,In_195);
and U888 (N_888,In_2415,In_2488);
nor U889 (N_889,In_2210,In_1377);
or U890 (N_890,In_2791,In_2752);
or U891 (N_891,In_1480,N_59);
nand U892 (N_892,In_242,In_2983);
nand U893 (N_893,N_383,N_262);
nand U894 (N_894,In_2380,In_887);
or U895 (N_895,In_945,In_750);
nand U896 (N_896,In_1606,In_2163);
nor U897 (N_897,In_57,N_559);
nor U898 (N_898,In_2066,In_1774);
and U899 (N_899,N_442,In_1921);
or U900 (N_900,N_850,In_1866);
and U901 (N_901,N_353,N_508);
and U902 (N_902,N_874,N_645);
nand U903 (N_903,In_1712,N_332);
nand U904 (N_904,In_1741,N_688);
or U905 (N_905,In_2680,N_681);
or U906 (N_906,In_1298,N_199);
nand U907 (N_907,N_290,N_510);
or U908 (N_908,N_680,N_470);
and U909 (N_909,N_32,N_235);
xnor U910 (N_910,In_2490,N_448);
or U911 (N_911,In_2623,In_299);
or U912 (N_912,In_387,In_1148);
or U913 (N_913,In_1949,N_627);
and U914 (N_914,N_648,N_326);
and U915 (N_915,In_392,N_433);
and U916 (N_916,N_847,In_405);
nand U917 (N_917,In_2333,In_1641);
nor U918 (N_918,In_958,In_1711);
and U919 (N_919,In_373,N_564);
nor U920 (N_920,In_1385,In_954);
nand U921 (N_921,In_516,In_1098);
nand U922 (N_922,In_1162,N_768);
nor U923 (N_923,N_511,In_1644);
xnor U924 (N_924,In_2780,In_2726);
nand U925 (N_925,In_1325,In_2937);
xnor U926 (N_926,In_394,In_828);
nor U927 (N_927,In_164,In_177);
nand U928 (N_928,In_173,In_606);
nor U929 (N_929,N_786,N_322);
nand U930 (N_930,In_845,N_351);
nor U931 (N_931,N_777,N_64);
or U932 (N_932,In_2588,N_861);
or U933 (N_933,N_428,N_836);
xor U934 (N_934,In_1150,In_835);
xor U935 (N_935,In_1979,In_2424);
and U936 (N_936,In_2990,In_366);
or U937 (N_937,In_2273,In_1926);
or U938 (N_938,In_2266,In_2555);
nor U939 (N_939,In_934,In_884);
and U940 (N_940,In_2314,N_267);
xnor U941 (N_941,In_2704,In_2064);
or U942 (N_942,In_2332,In_2606);
or U943 (N_943,In_2234,N_457);
xnor U944 (N_944,In_2896,In_2627);
or U945 (N_945,N_318,N_250);
or U946 (N_946,N_629,In_2059);
or U947 (N_947,In_199,In_970);
nand U948 (N_948,In_808,N_622);
or U949 (N_949,In_325,N_682);
nand U950 (N_950,N_838,N_299);
nand U951 (N_951,N_881,In_9);
xnor U952 (N_952,In_291,In_110);
nand U953 (N_953,In_256,In_1051);
nor U954 (N_954,In_1315,In_2383);
xor U955 (N_955,In_2939,In_2256);
and U956 (N_956,In_1429,In_1203);
or U957 (N_957,N_532,In_1654);
and U958 (N_958,In_118,N_487);
nand U959 (N_959,In_1233,N_148);
or U960 (N_960,In_39,N_697);
xor U961 (N_961,In_1998,In_2590);
xor U962 (N_962,In_1868,In_1068);
nor U963 (N_963,N_102,N_288);
and U964 (N_964,N_58,N_800);
or U965 (N_965,N_870,In_497);
and U966 (N_966,In_990,In_1271);
and U967 (N_967,N_650,In_2573);
nand U968 (N_968,In_615,In_414);
nand U969 (N_969,N_184,In_142);
xnor U970 (N_970,In_759,N_643);
nor U971 (N_971,In_2817,N_452);
and U972 (N_972,N_803,N_308);
xor U973 (N_973,In_2691,In_382);
xor U974 (N_974,N_22,In_2532);
and U975 (N_975,In_2113,In_2903);
and U976 (N_976,In_844,N_842);
nor U977 (N_977,In_2158,N_787);
xor U978 (N_978,In_2019,In_1529);
nor U979 (N_979,In_81,In_1594);
and U980 (N_980,In_2202,In_1675);
xnor U981 (N_981,In_663,N_711);
nor U982 (N_982,In_139,In_2426);
xor U983 (N_983,In_2980,In_1273);
nor U984 (N_984,N_134,In_691);
and U985 (N_985,N_233,N_200);
nand U986 (N_986,In_1689,In_2624);
nor U987 (N_987,In_122,In_350);
nand U988 (N_988,In_547,In_1917);
nand U989 (N_989,N_24,In_1836);
and U990 (N_990,N_17,In_1890);
or U991 (N_991,In_1227,In_770);
xnor U992 (N_992,In_2832,N_703);
or U993 (N_993,In_1660,In_1597);
xnor U994 (N_994,N_794,In_2982);
nor U995 (N_995,N_883,N_613);
nor U996 (N_996,In_2371,N_52);
nor U997 (N_997,N_379,In_2857);
nor U998 (N_998,In_1598,In_2343);
nor U999 (N_999,In_979,In_2260);
nand U1000 (N_1000,In_32,In_2219);
or U1001 (N_1001,In_1466,In_1485);
nor U1002 (N_1002,In_790,N_660);
nor U1003 (N_1003,In_843,In_1928);
nand U1004 (N_1004,In_2533,In_2865);
or U1005 (N_1005,N_867,In_1336);
xor U1006 (N_1006,In_2012,N_740);
nand U1007 (N_1007,In_438,N_123);
nand U1008 (N_1008,N_684,In_277);
nand U1009 (N_1009,N_261,N_10);
xnor U1010 (N_1010,In_1479,In_410);
xnor U1011 (N_1011,In_504,N_523);
nor U1012 (N_1012,In_993,In_1889);
and U1013 (N_1013,In_2797,In_228);
and U1014 (N_1014,In_45,In_1403);
and U1015 (N_1015,In_2191,In_1875);
nor U1016 (N_1016,In_2870,In_2861);
nand U1017 (N_1017,In_1168,In_2363);
nor U1018 (N_1018,In_2759,In_1084);
nor U1019 (N_1019,In_1381,N_733);
nand U1020 (N_1020,N_761,In_1112);
nor U1021 (N_1021,N_769,In_1104);
and U1022 (N_1022,N_588,In_717);
nor U1023 (N_1023,In_1100,In_925);
or U1024 (N_1024,N_69,In_1522);
and U1025 (N_1025,N_719,In_2873);
nor U1026 (N_1026,In_1461,In_1420);
or U1027 (N_1027,In_1130,In_341);
xnor U1028 (N_1028,In_2188,In_2397);
nand U1029 (N_1029,In_1464,In_1865);
or U1030 (N_1030,In_154,In_1574);
xnor U1031 (N_1031,In_1368,N_412);
nand U1032 (N_1032,In_2882,In_2209);
nor U1033 (N_1033,In_1008,In_2527);
or U1034 (N_1034,In_1073,N_159);
and U1035 (N_1035,In_2050,In_1781);
or U1036 (N_1036,N_387,N_306);
and U1037 (N_1037,In_2875,In_712);
nand U1038 (N_1038,In_648,In_1291);
nand U1039 (N_1039,N_716,In_1093);
or U1040 (N_1040,N_859,N_722);
xor U1041 (N_1041,In_2304,N_526);
nor U1042 (N_1042,In_1034,In_2461);
xnor U1043 (N_1043,In_2814,N_802);
nand U1044 (N_1044,In_1128,In_973);
nand U1045 (N_1045,In_192,In_548);
nor U1046 (N_1046,In_138,In_2885);
nand U1047 (N_1047,In_2619,In_2711);
and U1048 (N_1048,In_2916,In_1419);
or U1049 (N_1049,N_647,N_696);
and U1050 (N_1050,N_108,In_1351);
or U1051 (N_1051,In_1297,N_405);
nand U1052 (N_1052,In_2176,N_139);
xor U1053 (N_1053,N_813,In_2285);
and U1054 (N_1054,In_1877,N_467);
and U1055 (N_1055,In_650,N_73);
nor U1056 (N_1056,In_2307,In_2409);
xor U1057 (N_1057,In_2610,N_55);
or U1058 (N_1058,In_2909,N_283);
and U1059 (N_1059,In_1740,In_1173);
xnor U1060 (N_1060,N_793,In_2645);
xnor U1061 (N_1061,In_1386,In_1605);
nor U1062 (N_1062,In_1039,N_631);
nor U1063 (N_1063,N_517,In_2821);
or U1064 (N_1064,In_269,N_764);
nand U1065 (N_1065,In_348,In_1160);
and U1066 (N_1066,In_915,N_4);
nor U1067 (N_1067,In_2342,In_266);
nand U1068 (N_1068,In_239,N_178);
or U1069 (N_1069,In_2819,In_1972);
and U1070 (N_1070,In_601,In_2068);
xor U1071 (N_1071,In_1724,In_1246);
and U1072 (N_1072,N_789,N_304);
nor U1073 (N_1073,N_128,N_80);
or U1074 (N_1074,N_496,N_677);
nor U1075 (N_1075,N_62,In_1096);
nor U1076 (N_1076,In_2695,N_445);
xor U1077 (N_1077,In_2145,In_1344);
nor U1078 (N_1078,In_942,In_186);
xor U1079 (N_1079,In_1392,N_727);
or U1080 (N_1080,In_161,N_85);
or U1081 (N_1081,N_589,In_1348);
or U1082 (N_1082,In_1054,In_2190);
and U1083 (N_1083,In_1693,In_198);
or U1084 (N_1084,In_2949,In_1439);
xor U1085 (N_1085,In_80,In_2324);
or U1086 (N_1086,N_855,N_5);
xnor U1087 (N_1087,In_1723,In_881);
or U1088 (N_1088,In_330,In_649);
nor U1089 (N_1089,In_170,In_1595);
and U1090 (N_1090,N_686,In_1341);
or U1091 (N_1091,N_814,N_843);
and U1092 (N_1092,In_281,In_1475);
nand U1093 (N_1093,In_2006,N_298);
and U1094 (N_1094,In_60,In_672);
or U1095 (N_1095,In_271,In_1727);
nor U1096 (N_1096,N_860,In_2182);
nand U1097 (N_1097,N_817,N_825);
xor U1098 (N_1098,In_171,In_2979);
nand U1099 (N_1099,N_654,N_776);
nand U1100 (N_1100,In_2389,In_2453);
nand U1101 (N_1101,In_1765,In_2951);
and U1102 (N_1102,In_751,In_1442);
nor U1103 (N_1103,In_767,In_1975);
or U1104 (N_1104,In_2226,N_44);
or U1105 (N_1105,In_1408,N_661);
xor U1106 (N_1106,In_1978,In_534);
nand U1107 (N_1107,In_1259,N_81);
nor U1108 (N_1108,N_679,N_497);
nor U1109 (N_1109,In_1260,N_507);
and U1110 (N_1110,N_422,N_211);
nor U1111 (N_1111,In_2337,In_1528);
xnor U1112 (N_1112,In_677,In_948);
nor U1113 (N_1113,In_799,In_1097);
or U1114 (N_1114,N_628,In_94);
xnor U1115 (N_1115,In_1282,In_243);
xor U1116 (N_1116,In_2688,In_11);
nor U1117 (N_1117,In_55,N_675);
or U1118 (N_1118,In_1937,In_2716);
or U1119 (N_1119,In_478,In_404);
nand U1120 (N_1120,In_2472,N_620);
nand U1121 (N_1121,In_1648,N_100);
nand U1122 (N_1122,N_591,In_2868);
nand U1123 (N_1123,N_16,N_464);
nand U1124 (N_1124,In_1558,In_383);
xor U1125 (N_1125,N_171,In_1915);
xnor U1126 (N_1126,N_373,N_538);
and U1127 (N_1127,In_417,In_2793);
nand U1128 (N_1128,In_1532,In_1224);
nor U1129 (N_1129,N_466,In_810);
or U1130 (N_1130,In_2722,In_234);
nor U1131 (N_1131,In_2345,N_49);
nor U1132 (N_1132,In_379,N_451);
nand U1133 (N_1133,N_525,In_1421);
and U1134 (N_1134,N_888,In_1962);
xor U1135 (N_1135,In_37,In_1135);
nand U1136 (N_1136,N_544,In_542);
and U1137 (N_1137,In_1615,In_2950);
nor U1138 (N_1138,In_1656,N_839);
xor U1139 (N_1139,In_1286,In_1214);
and U1140 (N_1140,In_337,In_599);
nor U1141 (N_1141,N_303,In_1169);
and U1142 (N_1142,N_453,In_2425);
nor U1143 (N_1143,N_272,In_48);
or U1144 (N_1144,N_300,In_1860);
and U1145 (N_1145,In_2956,In_2280);
and U1146 (N_1146,N_57,In_1438);
nor U1147 (N_1147,N_110,In_1356);
nand U1148 (N_1148,In_2171,In_1187);
nand U1149 (N_1149,N_685,In_2179);
nor U1150 (N_1150,In_2041,In_1966);
nor U1151 (N_1151,In_1290,N_334);
nor U1152 (N_1152,N_882,In_2674);
and U1153 (N_1153,N_330,N_147);
or U1154 (N_1154,N_571,N_670);
xor U1155 (N_1155,N_743,N_107);
or U1156 (N_1156,In_1586,In_2911);
xor U1157 (N_1157,N_524,In_2603);
nor U1158 (N_1158,In_1472,In_2306);
nand U1159 (N_1159,In_1300,N_896);
and U1160 (N_1160,In_745,N_503);
nand U1161 (N_1161,In_1110,In_2626);
nand U1162 (N_1162,In_1736,In_1132);
nand U1163 (N_1163,N_706,N_691);
nand U1164 (N_1164,In_1215,In_719);
and U1165 (N_1165,In_984,N_884);
nand U1166 (N_1166,N_846,N_621);
and U1167 (N_1167,N_413,N_840);
nor U1168 (N_1168,In_2253,N_278);
nand U1169 (N_1169,In_789,N_666);
xnor U1170 (N_1170,In_2561,In_1513);
or U1171 (N_1171,N_29,In_1511);
nor U1172 (N_1172,N_898,In_1258);
and U1173 (N_1173,N_892,In_1518);
nand U1174 (N_1174,In_2257,In_1484);
xor U1175 (N_1175,In_1725,In_1831);
nor U1176 (N_1176,In_1995,In_2107);
or U1177 (N_1177,In_1069,In_496);
xnor U1178 (N_1178,In_978,In_2141);
nor U1179 (N_1179,In_2748,N_401);
nor U1180 (N_1180,N_206,In_2313);
or U1181 (N_1181,In_1832,In_1198);
xnor U1182 (N_1182,In_2489,In_803);
and U1183 (N_1183,N_594,In_1619);
and U1184 (N_1184,In_1694,In_252);
nor U1185 (N_1185,N_774,In_576);
nand U1186 (N_1186,N_287,In_2967);
or U1187 (N_1187,In_1663,In_832);
and U1188 (N_1188,In_849,In_235);
xor U1189 (N_1189,In_1913,N_545);
nand U1190 (N_1190,In_855,In_540);
nand U1191 (N_1191,In_2958,In_2413);
and U1192 (N_1192,In_2930,In_2749);
xor U1193 (N_1193,In_1256,In_2301);
xor U1194 (N_1194,In_2360,N_742);
xor U1195 (N_1195,In_1627,N_409);
nor U1196 (N_1196,In_1760,In_1547);
and U1197 (N_1197,N_791,In_1577);
and U1198 (N_1198,N_140,N_214);
nand U1199 (N_1199,In_1005,In_886);
nand U1200 (N_1200,N_601,In_2881);
nand U1201 (N_1201,In_1828,N_43);
nor U1202 (N_1202,In_2370,N_563);
and U1203 (N_1203,N_1194,In_233);
or U1204 (N_1204,In_316,N_748);
nor U1205 (N_1205,In_2594,N_665);
nor U1206 (N_1206,In_2075,In_2228);
and U1207 (N_1207,In_2584,In_2675);
xor U1208 (N_1208,N_577,N_583);
xor U1209 (N_1209,N_945,In_2746);
and U1210 (N_1210,N_1026,In_1786);
nor U1211 (N_1211,N_534,N_1130);
nor U1212 (N_1212,In_2079,In_1666);
and U1213 (N_1213,In_617,N_1095);
nand U1214 (N_1214,In_2466,N_1134);
nand U1215 (N_1215,N_819,N_1147);
xnor U1216 (N_1216,In_19,In_1024);
and U1217 (N_1217,In_2524,In_1205);
nand U1218 (N_1218,N_270,In_555);
nand U1219 (N_1219,N_792,In_471);
nor U1220 (N_1220,N_1150,In_1238);
or U1221 (N_1221,N_305,N_1156);
and U1222 (N_1222,In_1123,In_445);
and U1223 (N_1223,In_2894,In_2168);
and U1224 (N_1224,N_1041,N_598);
or U1225 (N_1225,In_2719,In_2277);
nand U1226 (N_1226,In_2931,N_230);
nor U1227 (N_1227,In_2900,In_2043);
and U1228 (N_1228,N_447,In_282);
nand U1229 (N_1229,N_34,In_123);
xor U1230 (N_1230,N_1098,N_617);
nand U1231 (N_1231,N_543,In_2667);
nand U1232 (N_1232,In_447,N_125);
xor U1233 (N_1233,In_302,In_2733);
and U1234 (N_1234,N_181,N_782);
xnor U1235 (N_1235,In_2212,In_320);
and U1236 (N_1236,N_145,In_2287);
xor U1237 (N_1237,In_1771,N_790);
and U1238 (N_1238,N_899,N_440);
xor U1239 (N_1239,In_47,In_1793);
nor U1240 (N_1240,In_273,N_721);
xor U1241 (N_1241,In_1878,In_2338);
or U1242 (N_1242,In_1850,N_806);
nand U1243 (N_1243,In_2898,In_2420);
or U1244 (N_1244,In_1810,N_921);
and U1245 (N_1245,In_2757,In_2431);
xor U1246 (N_1246,In_2449,N_1135);
or U1247 (N_1247,In_1628,In_1448);
and U1248 (N_1248,In_1715,In_2090);
xor U1249 (N_1249,In_1783,N_983);
nand U1250 (N_1250,In_1358,N_662);
nor U1251 (N_1251,In_1613,N_348);
nand U1252 (N_1252,In_219,In_911);
nor U1253 (N_1253,N_218,N_505);
nand U1254 (N_1254,In_1651,In_2092);
nor U1255 (N_1255,In_474,In_149);
nand U1256 (N_1256,In_1152,In_2504);
nand U1257 (N_1257,N_1015,N_984);
and U1258 (N_1258,N_455,N_63);
xor U1259 (N_1259,N_933,In_2936);
nor U1260 (N_1260,In_1643,N_117);
or U1261 (N_1261,N_831,In_552);
nand U1262 (N_1262,N_1022,In_960);
nor U1263 (N_1263,N_877,N_765);
xnor U1264 (N_1264,N_1078,In_1468);
and U1265 (N_1265,N_175,In_2888);
and U1266 (N_1266,In_1329,N_1033);
or U1267 (N_1267,In_697,N_1004);
nand U1268 (N_1268,In_216,In_2149);
nor U1269 (N_1269,N_307,N_203);
nand U1270 (N_1270,N_103,N_1090);
nor U1271 (N_1271,In_2503,N_1128);
or U1272 (N_1272,In_2117,N_25);
nor U1273 (N_1273,N_1084,In_2987);
xnor U1274 (N_1274,N_569,In_1839);
nor U1275 (N_1275,N_783,N_1120);
xnor U1276 (N_1276,In_2742,In_901);
and U1277 (N_1277,N_739,N_129);
and U1278 (N_1278,In_2807,In_470);
nor U1279 (N_1279,N_8,N_30);
nand U1280 (N_1280,In_1945,N_1159);
or U1281 (N_1281,In_1684,In_1006);
nand U1282 (N_1282,In_549,In_1299);
nand U1283 (N_1283,In_1721,In_513);
xnor U1284 (N_1284,In_1070,N_913);
xor U1285 (N_1285,In_2539,In_409);
nand U1286 (N_1286,In_1156,N_234);
and U1287 (N_1287,N_514,In_2072);
nand U1288 (N_1288,N_1046,In_2021);
or U1289 (N_1289,N_547,In_1289);
and U1290 (N_1290,In_630,In_1007);
xor U1291 (N_1291,In_1909,In_1940);
nand U1292 (N_1292,N_460,N_378);
nor U1293 (N_1293,N_639,In_389);
and U1294 (N_1294,N_937,N_1085);
and U1295 (N_1295,N_443,In_1707);
and U1296 (N_1296,In_2390,In_1816);
xnor U1297 (N_1297,In_2636,N_1176);
nand U1298 (N_1298,In_2364,In_2506);
or U1299 (N_1299,N_1066,In_2281);
nand U1300 (N_1300,N_1031,In_1794);
and U1301 (N_1301,N_923,N_897);
nor U1302 (N_1302,N_365,In_1941);
xnor U1303 (N_1303,In_327,N_700);
nor U1304 (N_1304,In_2459,In_51);
xor U1305 (N_1305,N_45,N_973);
nor U1306 (N_1306,N_835,In_582);
and U1307 (N_1307,In_158,In_412);
nand U1308 (N_1308,In_1099,N_1149);
and U1309 (N_1309,N_335,N_592);
nor U1310 (N_1310,In_2781,In_415);
or U1311 (N_1311,N_830,N_609);
xor U1312 (N_1312,N_1109,In_133);
or U1313 (N_1313,In_1002,In_655);
and U1314 (N_1314,In_98,In_2055);
or U1315 (N_1315,N_480,In_2644);
and U1316 (N_1316,N_1003,N_837);
or U1317 (N_1317,In_1304,In_2647);
and U1318 (N_1318,In_117,In_1762);
and U1319 (N_1319,N_911,In_2056);
or U1320 (N_1320,In_503,N_297);
or U1321 (N_1321,N_1162,In_217);
and U1322 (N_1322,N_1195,In_2482);
nand U1323 (N_1323,In_1616,In_2319);
nand U1324 (N_1324,In_809,In_1189);
and U1325 (N_1325,N_656,In_2974);
and U1326 (N_1326,N_1137,N_398);
nand U1327 (N_1327,N_539,In_864);
xor U1328 (N_1328,In_1682,N_309);
nand U1329 (N_1329,N_655,N_189);
nand U1330 (N_1330,N_1167,In_682);
xor U1331 (N_1331,In_393,N_1028);
nand U1332 (N_1332,In_1812,In_1953);
nor U1333 (N_1333,N_1192,N_762);
and U1334 (N_1334,N_51,In_1040);
and U1335 (N_1335,In_290,N_291);
xnor U1336 (N_1336,In_2585,N_1076);
nand U1337 (N_1337,In_2578,N_615);
or U1338 (N_1338,In_2052,In_2367);
nor U1339 (N_1339,In_1742,In_1911);
nand U1340 (N_1340,N_1179,N_255);
nor U1341 (N_1341,In_423,In_575);
or U1342 (N_1342,N_943,In_1500);
xnor U1343 (N_1343,N_1187,In_1144);
nand U1344 (N_1344,N_638,N_324);
xnor U1345 (N_1345,In_2615,In_2200);
nand U1346 (N_1346,In_1044,N_369);
nand U1347 (N_1347,In_75,N_974);
and U1348 (N_1348,N_865,In_1317);
nor U1349 (N_1349,In_2671,N_93);
and U1350 (N_1350,In_2471,In_1369);
nor U1351 (N_1351,N_490,In_2152);
and U1352 (N_1352,In_2,N_210);
xor U1353 (N_1353,In_2028,N_1125);
xor U1354 (N_1354,In_1208,In_2884);
xnor U1355 (N_1355,N_956,In_2040);
nor U1356 (N_1356,In_112,In_1415);
and U1357 (N_1357,In_1818,N_88);
nand U1358 (N_1358,In_681,In_1020);
nand U1359 (N_1359,In_2634,N_165);
nor U1360 (N_1360,In_2034,In_2534);
and U1361 (N_1361,In_519,N_454);
nor U1362 (N_1362,In_1083,N_150);
and U1363 (N_1363,N_1153,N_575);
or U1364 (N_1364,N_779,In_674);
nor U1365 (N_1365,In_1782,In_2411);
xnor U1366 (N_1366,In_2245,In_40);
or U1367 (N_1367,N_1042,In_525);
nor U1368 (N_1368,N_678,N_1062);
and U1369 (N_1369,In_2761,N_853);
xor U1370 (N_1370,N_848,N_824);
nor U1371 (N_1371,In_1942,N_493);
and U1372 (N_1372,In_431,In_2744);
nor U1373 (N_1373,N_1132,N_607);
and U1374 (N_1374,N_1057,In_2388);
nand U1375 (N_1375,N_372,N_862);
xor U1376 (N_1376,N_358,In_2305);
nor U1377 (N_1377,In_1817,In_2137);
or U1378 (N_1378,N_641,N_1013);
xor U1379 (N_1379,In_1465,N_341);
nor U1380 (N_1380,N_1010,N_737);
nand U1381 (N_1381,N_1054,N_402);
or U1382 (N_1382,In_500,In_1685);
nor U1383 (N_1383,N_775,N_530);
and U1384 (N_1384,In_2790,In_1881);
and U1385 (N_1385,In_999,In_2298);
or U1386 (N_1386,N_625,N_864);
or U1387 (N_1387,In_1789,N_935);
or U1388 (N_1388,N_618,In_2995);
and U1389 (N_1389,N_1044,In_167);
nand U1390 (N_1390,In_1957,N_1101);
nor U1391 (N_1391,N_1191,In_1635);
nor U1392 (N_1392,In_1555,In_1826);
xor U1393 (N_1393,In_1445,In_1202);
xnor U1394 (N_1394,N_492,N_133);
xor U1395 (N_1395,N_1172,In_2416);
nand U1396 (N_1396,In_642,In_321);
xnor U1397 (N_1397,N_924,In_1155);
and U1398 (N_1398,In_1743,N_844);
and U1399 (N_1399,N_195,In_1017);
and U1400 (N_1400,N_439,N_887);
or U1401 (N_1401,In_2867,N_658);
and U1402 (N_1402,In_489,In_2195);
nor U1403 (N_1403,N_459,N_295);
xnor U1404 (N_1404,N_997,In_332);
xnor U1405 (N_1405,N_942,N_391);
and U1406 (N_1406,In_907,In_1837);
xor U1407 (N_1407,N_816,N_606);
xnor U1408 (N_1408,In_1217,N_713);
nor U1409 (N_1409,In_467,In_413);
nor U1410 (N_1410,In_2186,In_1087);
xor U1411 (N_1411,N_975,In_1116);
nor U1412 (N_1412,In_2110,In_981);
xnor U1413 (N_1413,In_2665,N_484);
xnor U1414 (N_1414,In_997,N_1138);
and U1415 (N_1415,In_1732,N_1051);
and U1416 (N_1416,In_246,In_2181);
or U1417 (N_1417,In_2815,In_1661);
and U1418 (N_1418,In_2445,N_1106);
nand U1419 (N_1419,In_59,In_1248);
or U1420 (N_1420,N_828,In_2216);
or U1421 (N_1421,In_1849,In_536);
and U1422 (N_1422,In_1596,N_86);
xor U1423 (N_1423,N_465,N_893);
nor U1424 (N_1424,In_2863,In_2643);
or U1425 (N_1425,N_967,N_407);
nand U1426 (N_1426,N_106,N_217);
nand U1427 (N_1427,In_102,N_821);
and U1428 (N_1428,N_520,N_276);
xnor U1429 (N_1429,N_1032,In_70);
and U1430 (N_1430,N_476,N_798);
xnor U1431 (N_1431,In_872,In_2505);
xor U1432 (N_1432,In_106,N_1055);
xor U1433 (N_1433,In_371,N_925);
nand U1434 (N_1434,N_698,In_1321);
or U1435 (N_1435,In_1955,N_672);
xnor U1436 (N_1436,N_1122,In_369);
and U1437 (N_1437,N_747,In_1340);
nand U1438 (N_1438,In_2334,In_514);
nor U1439 (N_1439,N_610,N_1000);
nand U1440 (N_1440,N_362,In_12);
xnor U1441 (N_1441,In_457,In_2721);
and U1442 (N_1442,In_594,In_2172);
nor U1443 (N_1443,In_1328,N_188);
xor U1444 (N_1444,In_2121,In_42);
nand U1445 (N_1445,In_50,In_343);
nor U1446 (N_1446,In_2496,N_1035);
or U1447 (N_1447,N_1045,N_812);
nor U1448 (N_1448,In_2458,In_334);
nor U1449 (N_1449,N_316,N_1136);
and U1450 (N_1450,N_972,In_88);
nor U1451 (N_1451,N_759,N_845);
and U1452 (N_1452,N_65,N_938);
xor U1453 (N_1453,In_2289,N_1100);
and U1454 (N_1454,In_331,N_833);
nor U1455 (N_1455,N_724,N_926);
and U1456 (N_1456,N_1058,In_730);
or U1457 (N_1457,N_1114,In_690);
and U1458 (N_1458,In_564,In_1414);
xnor U1459 (N_1459,N_1048,In_1492);
or U1460 (N_1460,In_1470,N_529);
or U1461 (N_1461,N_906,N_580);
xor U1462 (N_1462,In_1515,In_1079);
nand U1463 (N_1463,In_2270,N_271);
and U1464 (N_1464,In_2497,In_2361);
xnor U1465 (N_1465,N_562,N_337);
nor U1466 (N_1466,In_2905,N_220);
xor U1467 (N_1467,N_1089,In_1785);
or U1468 (N_1468,In_1313,N_674);
xnor U1469 (N_1469,In_533,In_1633);
xor U1470 (N_1470,In_2331,In_1383);
nor U1471 (N_1471,In_2724,N_95);
xor U1472 (N_1472,N_1008,N_435);
or U1473 (N_1473,In_1905,N_1144);
and U1474 (N_1474,N_632,In_2650);
xor U1475 (N_1475,N_750,In_116);
xnor U1476 (N_1476,In_2001,In_1446);
nand U1477 (N_1477,In_706,In_578);
and U1478 (N_1478,In_1642,In_1883);
and U1479 (N_1479,N_668,In_1004);
xnor U1480 (N_1480,In_511,N_346);
xnor U1481 (N_1481,In_1462,N_1025);
and U1482 (N_1482,N_738,In_2126);
or U1483 (N_1483,N_399,In_95);
and U1484 (N_1484,N_1024,In_2214);
xnor U1485 (N_1485,In_1272,In_2350);
nor U1486 (N_1486,N_663,In_2250);
nand U1487 (N_1487,In_1650,N_876);
and U1488 (N_1488,In_137,N_1148);
nor U1489 (N_1489,In_652,In_2668);
and U1490 (N_1490,N_121,In_2340);
nor U1491 (N_1491,In_360,N_479);
nand U1492 (N_1492,In_791,N_873);
and U1493 (N_1493,N_822,N_1189);
nand U1494 (N_1494,In_2703,N_1067);
nand U1495 (N_1495,In_969,In_1952);
nand U1496 (N_1496,In_17,N_521);
or U1497 (N_1497,N_1163,In_2443);
nand U1498 (N_1498,In_1266,In_1292);
xnor U1499 (N_1499,N_560,N_1091);
or U1500 (N_1500,N_1407,In_2401);
or U1501 (N_1501,In_249,In_701);
or U1502 (N_1502,In_1801,N_1246);
nand U1503 (N_1503,In_317,N_1123);
or U1504 (N_1504,In_1731,N_1310);
nor U1505 (N_1505,N_1080,In_185);
nand U1506 (N_1506,N_223,In_2162);
and U1507 (N_1507,N_1426,N_1296);
or U1508 (N_1508,N_1392,In_7);
and U1509 (N_1509,In_1337,N_669);
xor U1510 (N_1510,N_941,In_716);
nor U1511 (N_1511,N_352,In_1824);
xor U1512 (N_1512,N_1227,N_1182);
xnor U1513 (N_1513,N_1419,N_1364);
or U1514 (N_1514,N_1294,In_912);
and U1515 (N_1515,N_1353,N_708);
nor U1516 (N_1516,N_1249,N_1216);
nor U1517 (N_1517,In_2786,In_1264);
nor U1518 (N_1518,N_551,N_1330);
nand U1519 (N_1519,N_1184,N_437);
nand U1520 (N_1520,N_1317,In_928);
xor U1521 (N_1521,N_832,In_307);
nor U1522 (N_1522,N_1324,N_1140);
xor U1523 (N_1523,In_1610,N_190);
and U1524 (N_1524,N_985,In_2955);
and U1525 (N_1525,N_797,N_734);
and U1526 (N_1526,N_1225,N_557);
xor U1527 (N_1527,In_1677,N_1235);
nand U1528 (N_1528,N_2,In_2841);
or U1529 (N_1529,N_380,N_1139);
nor U1530 (N_1530,In_2071,In_1507);
and U1531 (N_1531,N_718,In_1923);
nor U1532 (N_1532,N_1454,In_65);
nand U1533 (N_1533,N_1462,N_1369);
and U1534 (N_1534,In_2978,In_773);
nor U1535 (N_1535,N_695,N_1020);
xor U1536 (N_1536,In_1375,N_1372);
nor U1537 (N_1537,In_381,N_1115);
xor U1538 (N_1538,N_1455,N_603);
or U1539 (N_1539,N_531,In_1181);
nor U1540 (N_1540,N_970,N_500);
and U1541 (N_1541,In_735,N_728);
and U1542 (N_1542,N_1142,In_38);
and U1543 (N_1543,N_550,In_2078);
nor U1544 (N_1544,In_2705,In_2970);
nand U1545 (N_1545,In_351,In_2621);
and U1546 (N_1546,N_97,In_2403);
nand U1547 (N_1547,In_1779,In_2947);
and U1548 (N_1548,N_805,In_2398);
nor U1549 (N_1549,In_2478,In_2660);
or U1550 (N_1550,N_360,In_1053);
nor U1551 (N_1551,N_1269,In_2772);
nand U1552 (N_1552,In_223,In_2564);
and U1553 (N_1553,N_744,N_1061);
xor U1554 (N_1554,N_506,In_1943);
and U1555 (N_1555,N_953,N_406);
nor U1556 (N_1556,In_1709,In_1907);
xor U1557 (N_1557,N_980,N_1422);
xnor U1558 (N_1558,N_338,N_916);
xnor U1559 (N_1559,N_1319,N_948);
or U1560 (N_1560,In_144,In_1288);
nand U1561 (N_1561,N_1117,In_2526);
nor U1562 (N_1562,In_1422,N_1288);
or U1563 (N_1563,N_715,In_955);
or U1564 (N_1564,In_2932,In_1988);
or U1565 (N_1565,In_1591,N_910);
or U1566 (N_1566,N_1014,In_2659);
nand U1567 (N_1567,In_2081,In_2441);
nand U1568 (N_1568,N_1224,N_1488);
nor U1569 (N_1569,N_596,N_694);
xnor U1570 (N_1570,N_1447,N_1009);
and U1571 (N_1571,N_1424,N_579);
xor U1572 (N_1572,In_1504,N_1442);
nor U1573 (N_1573,In_1538,N_1457);
nor U1574 (N_1574,N_1209,N_732);
xor U1575 (N_1575,In_26,N_553);
xor U1576 (N_1576,N_1466,In_1820);
nor U1577 (N_1577,In_2376,N_418);
nor U1578 (N_1578,In_480,N_527);
and U1579 (N_1579,N_1380,N_915);
nand U1580 (N_1580,In_2835,In_985);
nand U1581 (N_1581,In_1932,N_94);
nand U1582 (N_1582,In_181,In_2271);
and U1583 (N_1583,N_1043,N_1190);
xor U1584 (N_1584,In_204,In_2512);
nor U1585 (N_1585,N_890,In_2924);
xor U1586 (N_1586,N_920,N_1291);
and U1587 (N_1587,N_649,In_1210);
and U1588 (N_1588,In_1769,In_2639);
xor U1589 (N_1589,N_1094,N_1469);
or U1590 (N_1590,N_1282,N_552);
or U1591 (N_1591,In_641,In_1483);
and U1592 (N_1592,In_1434,N_1157);
nor U1593 (N_1593,N_979,In_495);
and U1594 (N_1594,N_468,In_2153);
nor U1595 (N_1595,In_1872,N_114);
nand U1596 (N_1596,N_1409,N_1377);
nor U1597 (N_1597,N_781,In_951);
nor U1598 (N_1598,In_134,In_976);
xnor U1599 (N_1599,In_2010,In_570);
xor U1600 (N_1600,N_1493,N_1047);
nor U1601 (N_1601,N_1056,N_863);
nand U1602 (N_1602,N_1428,In_1806);
or U1603 (N_1603,In_2476,In_2499);
xnor U1604 (N_1604,In_1065,N_275);
nand U1605 (N_1605,In_2735,In_2131);
and U1606 (N_1606,In_1306,In_1199);
nor U1607 (N_1607,In_2986,N_1232);
and U1608 (N_1608,N_70,N_434);
or U1609 (N_1609,In_1396,In_2127);
or U1610 (N_1610,N_652,N_1475);
nor U1611 (N_1611,N_1073,In_2605);
and U1612 (N_1612,N_282,In_591);
nand U1613 (N_1613,N_644,N_1385);
nand U1614 (N_1614,In_2968,N_1443);
xnor U1615 (N_1615,N_624,In_439);
nor U1616 (N_1616,N_683,In_1350);
and U1617 (N_1617,N_301,In_1003);
xnor U1618 (N_1618,N_690,N_1335);
nor U1619 (N_1619,In_1201,N_872);
nor U1620 (N_1620,N_131,In_1075);
or U1621 (N_1621,N_955,N_852);
nand U1622 (N_1622,N_41,In_1357);
nand U1623 (N_1623,In_1284,In_329);
or U1624 (N_1624,In_524,In_1898);
and U1625 (N_1625,N_1145,In_140);
xor U1626 (N_1626,N_427,In_336);
nand U1627 (N_1627,In_1608,In_841);
or U1628 (N_1628,N_1266,In_846);
and U1629 (N_1629,In_1294,N_151);
and U1630 (N_1630,In_800,In_1632);
nor U1631 (N_1631,In_1146,N_586);
nor U1632 (N_1632,In_202,In_54);
and U1633 (N_1633,N_1487,N_1360);
and U1634 (N_1634,In_115,N_77);
nand U1635 (N_1635,N_441,In_53);
and U1636 (N_1636,In_2084,N_141);
and U1637 (N_1637,In_1149,N_403);
nand U1638 (N_1638,N_1370,In_824);
and U1639 (N_1639,N_889,N_1183);
or U1640 (N_1640,N_1119,In_2213);
nor U1641 (N_1641,N_226,N_595);
xnor U1642 (N_1642,In_2038,In_804);
and U1643 (N_1643,N_1060,In_367);
and U1644 (N_1644,In_1861,In_2813);
xnor U1645 (N_1645,In_508,N_749);
nand U1646 (N_1646,In_407,N_1284);
and U1647 (N_1647,N_1347,N_1069);
or U1648 (N_1648,N_1229,In_626);
or U1649 (N_1649,In_46,N_1270);
or U1650 (N_1650,In_2878,N_756);
nand U1651 (N_1651,N_1431,In_1253);
or U1652 (N_1652,In_820,In_213);
xnor U1653 (N_1653,N_1006,N_89);
xnor U1654 (N_1654,N_950,N_28);
or U1655 (N_1655,In_1956,N_785);
and U1656 (N_1656,In_893,N_1039);
nor U1657 (N_1657,N_84,N_1241);
xnor U1658 (N_1658,N_834,In_2387);
or U1659 (N_1659,N_667,N_1478);
xnor U1660 (N_1660,In_2230,In_1323);
nor U1661 (N_1661,In_2913,N_1260);
xnor U1662 (N_1662,N_549,N_1331);
or U1663 (N_1663,In_365,In_2754);
xor U1664 (N_1664,In_968,In_2825);
or U1665 (N_1665,In_2740,N_826);
xor U1666 (N_1666,N_1301,N_1433);
xnor U1667 (N_1667,In_811,N_635);
nand U1668 (N_1668,In_2912,N_1238);
xor U1669 (N_1669,N_1268,In_2016);
nand U1670 (N_1670,N_79,N_1316);
and U1671 (N_1671,N_205,N_1173);
xor U1672 (N_1672,N_1304,In_2838);
xor U1673 (N_1673,N_1420,N_815);
nand U1674 (N_1674,N_469,N_1197);
xnor U1675 (N_1675,N_1289,In_1401);
nor U1676 (N_1676,In_402,In_255);
nand U1677 (N_1677,N_1387,N_1274);
and U1678 (N_1678,N_1483,N_1155);
xnor U1679 (N_1679,N_1121,N_385);
nand U1680 (N_1680,N_1093,N_961);
and U1681 (N_1681,N_1350,N_366);
xnor U1682 (N_1682,N_664,In_184);
xnor U1683 (N_1683,N_246,N_788);
and U1684 (N_1684,N_1244,N_96);
nand U1685 (N_1685,In_2651,N_971);
or U1686 (N_1686,N_992,N_328);
or U1687 (N_1687,N_1338,In_2806);
nand U1688 (N_1688,In_2217,In_2160);
or U1689 (N_1689,N_1359,N_1313);
and U1690 (N_1690,In_136,N_1391);
nor U1691 (N_1691,N_265,N_1437);
xnor U1692 (N_1692,In_1894,In_2029);
nor U1693 (N_1693,N_707,In_1841);
nor U1694 (N_1694,In_1993,In_900);
nand U1695 (N_1695,N_1171,N_78);
nand U1696 (N_1696,N_1300,N_9);
xor U1697 (N_1697,In_515,N_1245);
or U1698 (N_1698,N_1005,N_567);
or U1699 (N_1699,In_1705,N_1256);
and U1700 (N_1700,N_919,N_1393);
nand U1701 (N_1701,N_996,In_1951);
nor U1702 (N_1702,N_758,N_689);
nor U1703 (N_1703,N_633,N_194);
nand U1704 (N_1704,In_512,In_352);
nand U1705 (N_1705,N_1297,N_1474);
nand U1706 (N_1706,N_264,In_1668);
nand U1707 (N_1707,In_1505,In_113);
nor U1708 (N_1708,N_857,N_1065);
and U1709 (N_1709,In_292,N_193);
and U1710 (N_1710,In_187,N_1450);
and U1711 (N_1711,In_2382,In_875);
or U1712 (N_1712,N_951,In_2347);
and U1713 (N_1713,In_1174,N_676);
nand U1714 (N_1714,In_579,In_1502);
xnor U1715 (N_1715,N_126,N_702);
or U1716 (N_1716,N_561,In_1451);
and U1717 (N_1717,In_159,N_994);
xor U1718 (N_1718,N_1050,N_1206);
and U1719 (N_1719,In_437,N_917);
nor U1720 (N_1720,N_1204,In_632);
or U1721 (N_1721,N_1485,N_957);
and U1722 (N_1722,In_1563,In_1049);
or U1723 (N_1723,In_215,In_1840);
xor U1724 (N_1724,In_2166,N_912);
xor U1725 (N_1725,N_1479,In_338);
nand U1726 (N_1726,In_1250,N_1152);
nor U1727 (N_1727,In_780,N_471);
and U1728 (N_1728,N_504,In_1145);
nor U1729 (N_1729,N_1314,In_230);
or U1730 (N_1730,In_1931,N_1063);
and U1731 (N_1731,N_1435,N_1396);
nand U1732 (N_1732,In_276,In_1095);
nand U1733 (N_1733,N_1165,N_880);
xnor U1734 (N_1734,In_2720,In_1612);
or U1735 (N_1735,N_486,In_1636);
and U1736 (N_1736,N_602,In_2422);
nor U1737 (N_1737,N_1401,N_518);
nand U1738 (N_1738,In_1391,In_2876);
nand U1739 (N_1739,N_820,N_196);
nor U1740 (N_1740,In_1,In_2315);
or U1741 (N_1741,In_975,In_1645);
and U1742 (N_1742,In_1077,N_1390);
nand U1743 (N_1743,In_1186,N_162);
nor U1744 (N_1744,In_1363,N_263);
xnor U1745 (N_1745,In_1756,N_634);
xnor U1746 (N_1746,In_927,In_1657);
nor U1747 (N_1747,N_1328,N_1034);
xor U1748 (N_1748,In_1607,In_448);
and U1749 (N_1749,In_1453,In_2822);
and U1750 (N_1750,In_2897,N_1262);
xnor U1751 (N_1751,In_114,N_1308);
or U1752 (N_1752,N_593,In_2326);
xnor U1753 (N_1753,N_371,In_2669);
nand U1754 (N_1754,In_1897,In_2850);
nor U1755 (N_1755,N_1305,In_182);
nand U1756 (N_1756,In_1934,In_1449);
and U1757 (N_1757,N_939,In_279);
nor U1758 (N_1758,N_208,In_455);
or U1759 (N_1759,N_342,N_1242);
or U1760 (N_1760,N_735,In_2267);
nand U1761 (N_1761,N_432,N_154);
or U1762 (N_1762,N_204,N_375);
nand U1763 (N_1763,N_630,N_491);
nor U1764 (N_1764,In_870,N_1410);
or U1765 (N_1765,In_787,In_2009);
nand U1766 (N_1766,In_2799,N_1030);
nor U1767 (N_1767,N_1215,In_2492);
nand U1768 (N_1768,In_1237,In_1342);
and U1769 (N_1769,N_1416,In_2053);
or U1770 (N_1770,N_730,In_2022);
or U1771 (N_1771,In_1314,N_225);
and U1772 (N_1772,N_964,In_2296);
nand U1773 (N_1773,N_946,In_99);
or U1774 (N_1774,In_2648,In_764);
nor U1775 (N_1775,N_717,N_928);
nand U1776 (N_1776,N_1210,In_2095);
nor U1777 (N_1777,N_374,In_1398);
and U1778 (N_1778,N_693,In_1950);
xor U1779 (N_1779,N_753,In_1285);
and U1780 (N_1780,N_849,N_105);
xor U1781 (N_1781,N_132,N_771);
and U1782 (N_1782,N_1082,N_1275);
or U1783 (N_1783,N_949,In_2375);
xor U1784 (N_1784,In_1954,In_523);
nand U1785 (N_1785,N_993,N_31);
or U1786 (N_1786,In_1057,N_1087);
nand U1787 (N_1787,In_2125,N_1208);
and U1788 (N_1788,In_1035,In_2237);
or U1789 (N_1789,N_1345,In_2519);
nand U1790 (N_1790,In_1822,In_1910);
nor U1791 (N_1791,N_1252,In_702);
or U1792 (N_1792,N_1448,N_1470);
xnor U1793 (N_1793,In_1362,N_657);
or U1794 (N_1794,N_1077,N_357);
nor U1795 (N_1795,N_934,N_554);
or U1796 (N_1796,N_1318,In_823);
or U1797 (N_1797,In_2385,N_807);
and U1798 (N_1798,In_2837,N_1311);
xor U1799 (N_1799,In_349,N_605);
and U1800 (N_1800,N_1570,In_2480);
and U1801 (N_1801,In_2545,In_2436);
and U1802 (N_1802,In_130,N_1665);
nand U1803 (N_1803,N_1012,N_710);
nor U1804 (N_1804,In_108,N_1516);
nor U1805 (N_1805,In_621,In_1220);
nand U1806 (N_1806,In_460,N_1271);
or U1807 (N_1807,N_1783,N_1445);
xnor U1808 (N_1808,N_1560,In_1055);
or U1809 (N_1809,In_1688,N_885);
nand U1810 (N_1810,N_1750,In_1565);
xor U1811 (N_1811,In_82,In_1703);
and U1812 (N_1812,N_1366,In_2346);
nor U1813 (N_1813,In_590,N_932);
and U1814 (N_1814,N_640,In_1206);
xnor U1815 (N_1815,In_733,N_485);
nand U1816 (N_1816,N_386,N_1543);
nor U1817 (N_1817,N_494,N_1257);
nand U1818 (N_1818,N_990,N_66);
xnor U1819 (N_1819,N_1415,In_1441);
nand U1820 (N_1820,N_900,N_930);
or U1821 (N_1821,In_2448,N_1592);
or U1822 (N_1822,N_1730,N_1444);
nor U1823 (N_1823,N_1436,N_959);
xor U1824 (N_1824,In_2654,N_1512);
or U1825 (N_1825,N_1361,In_1488);
xnor U1826 (N_1826,In_2762,In_956);
nand U1827 (N_1827,In_363,In_119);
xor U1828 (N_1828,N_1645,N_986);
nor U1829 (N_1829,N_1663,In_462);
or U1830 (N_1830,N_1749,N_38);
and U1831 (N_1831,N_1200,In_2731);
and U1832 (N_1832,In_2088,N_1752);
nand U1833 (N_1833,In_2869,N_801);
nand U1834 (N_1834,N_1354,In_62);
nand U1835 (N_1835,N_1577,N_1344);
nor U1836 (N_1836,N_327,N_424);
xnor U1837 (N_1837,N_1620,N_1341);
xor U1838 (N_1838,In_1752,N_1086);
xor U1839 (N_1839,In_2812,In_857);
nand U1840 (N_1840,N_1686,N_637);
nor U1841 (N_1841,N_1799,N_1207);
nand U1842 (N_1842,N_1343,N_1666);
nand U1843 (N_1843,In_1218,N_1452);
nand U1844 (N_1844,N_1482,In_1604);
or U1845 (N_1845,N_1217,In_2874);
nor U1846 (N_1846,N_1541,In_2177);
xor U1847 (N_1847,N_1507,N_704);
nor U1848 (N_1848,N_182,N_1309);
nor U1849 (N_1849,N_1563,In_2862);
nor U1850 (N_1850,N_878,N_1471);
xnor U1851 (N_1851,N_1212,N_1695);
xor U1852 (N_1852,N_1386,In_2120);
nand U1853 (N_1853,N_1672,N_1351);
nor U1854 (N_1854,N_725,In_2143);
nand U1855 (N_1855,N_1124,N_1565);
nand U1856 (N_1856,N_1792,N_1237);
and U1857 (N_1857,N_1320,N_1637);
nand U1858 (N_1858,In_577,N_1669);
nor U1859 (N_1859,N_1389,N_851);
xor U1860 (N_1860,N_1786,In_2601);
or U1861 (N_1861,In_1103,In_2672);
xnor U1862 (N_1862,In_2714,In_1768);
xnor U1863 (N_1863,In_1481,N_1612);
nor U1864 (N_1864,In_539,N_42);
and U1865 (N_1865,N_868,N_1617);
and U1866 (N_1866,N_1605,N_1705);
and U1867 (N_1867,N_180,In_2551);
or U1868 (N_1868,In_1562,N_321);
xnor U1869 (N_1869,In_287,In_1435);
nand U1870 (N_1870,N_1213,N_1203);
or U1871 (N_1871,N_1589,In_826);
nor U1872 (N_1872,In_518,N_1710);
nand U1873 (N_1873,N_1264,N_858);
xor U1874 (N_1874,N_1747,N_1405);
or U1875 (N_1875,N_1733,In_1584);
nor U1876 (N_1876,N_1576,N_1129);
or U1877 (N_1877,N_537,In_436);
and U1878 (N_1878,In_2586,In_66);
or U1879 (N_1879,N_1530,N_1583);
nand U1880 (N_1880,N_841,N_1181);
nand U1881 (N_1881,N_1631,In_303);
nor U1882 (N_1882,N_799,N_244);
nor U1883 (N_1883,In_2259,N_1439);
and U1884 (N_1884,In_1249,N_1691);
or U1885 (N_1885,In_1347,In_1697);
nor U1886 (N_1886,In_2318,N_1248);
xor U1887 (N_1887,N_1337,N_1598);
and U1888 (N_1888,N_1107,N_1394);
nor U1889 (N_1889,N_1169,N_1768);
xor U1890 (N_1890,In_704,In_583);
or U1891 (N_1891,N_741,In_2710);
and U1892 (N_1892,N_1704,N_1722);
nor U1893 (N_1893,N_1524,N_1538);
nor U1894 (N_1894,N_1406,N_257);
or U1895 (N_1895,In_200,N_1326);
nor U1896 (N_1896,In_238,N_1703);
and U1897 (N_1897,In_2934,N_918);
nand U1898 (N_1898,In_935,In_1624);
and U1899 (N_1899,In_818,In_2391);
or U1900 (N_1900,N_1606,N_1644);
and U1901 (N_1901,N_597,In_1795);
nor U1902 (N_1902,N_1739,In_1460);
and U1903 (N_1903,N_1534,N_277);
and U1904 (N_1904,N_1585,N_168);
nand U1905 (N_1905,N_1408,In_2734);
nor U1906 (N_1906,N_578,N_1717);
nor U1907 (N_1907,N_1234,N_280);
or U1908 (N_1908,N_1336,N_1529);
or U1909 (N_1909,In_2303,N_1547);
or U1910 (N_1910,N_1647,N_1535);
or U1911 (N_1911,N_1740,In_49);
nand U1912 (N_1912,N_1616,N_1019);
and U1913 (N_1913,N_1412,In_1254);
xor U1914 (N_1914,N_1052,In_2251);
or U1915 (N_1915,N_1795,N_1484);
xor U1916 (N_1916,N_1654,In_2292);
xor U1917 (N_1917,In_1519,N_770);
nand U1918 (N_1918,N_1160,N_1295);
nor U1919 (N_1919,N_823,N_1681);
and U1920 (N_1920,In_1647,N_1021);
xor U1921 (N_1921,In_1986,N_311);
or U1922 (N_1922,N_1720,N_636);
nor U1923 (N_1923,N_576,N_1685);
nand U1924 (N_1924,In_2801,N_1675);
xnor U1925 (N_1925,N_1254,N_1402);
xnor U1926 (N_1926,In_2895,N_1568);
or U1927 (N_1927,N_1280,N_1682);
nand U1928 (N_1928,N_1127,N_1782);
nand U1929 (N_1929,N_1554,N_1712);
and U1930 (N_1930,N_163,In_377);
or U1931 (N_1931,In_1780,N_1239);
or U1932 (N_1932,N_1092,In_2124);
nand U1933 (N_1933,N_963,N_1688);
nand U1934 (N_1934,In_679,N_1158);
and U1935 (N_1935,N_1357,In_939);
and U1936 (N_1936,N_1143,In_2779);
and U1937 (N_1937,N_1223,N_976);
and U1938 (N_1938,In_505,N_1597);
or U1939 (N_1939,N_1536,N_1713);
and U1940 (N_1940,N_1755,N_1643);
nand U1941 (N_1941,In_2495,N_1677);
or U1942 (N_1942,N_1011,In_1436);
and U1943 (N_1943,In_2568,N_1465);
and U1944 (N_1944,N_1762,N_626);
or U1945 (N_1945,N_931,N_1615);
xor U1946 (N_1946,N_1413,N_1567);
or U1947 (N_1947,N_1709,N_720);
or U1948 (N_1948,N_1578,N_1706);
nand U1949 (N_1949,N_1517,In_274);
nand U1950 (N_1950,In_1573,N_555);
or U1951 (N_1951,In_1378,N_444);
or U1952 (N_1952,N_1629,N_1040);
nand U1953 (N_1953,N_1684,In_262);
and U1954 (N_1954,N_245,In_2140);
or U1955 (N_1955,In_1739,In_675);
xnor U1956 (N_1956,N_1103,N_1151);
nor U1957 (N_1957,N_1676,N_1352);
or U1958 (N_1958,N_1588,In_435);
nor U1959 (N_1959,In_971,N_1774);
nor U1960 (N_1960,N_339,N_1521);
xor U1961 (N_1961,N_1542,N_767);
and U1962 (N_1962,N_1477,In_1399);
and U1963 (N_1963,In_306,N_1594);
or U1964 (N_1964,In_2203,N_1557);
or U1965 (N_1965,N_1425,N_709);
nor U1966 (N_1966,N_1580,In_2015);
and U1967 (N_1967,In_2205,N_1404);
nor U1968 (N_1968,N_1368,N_1562);
and U1969 (N_1969,N_1027,In_1185);
and U1970 (N_1970,N_616,In_1985);
xor U1971 (N_1971,In_2766,N_1007);
nand U1972 (N_1972,In_1924,N_1398);
or U1973 (N_1973,In_354,N_922);
nor U1974 (N_1974,In_314,N_1417);
nand U1975 (N_1975,N_1481,N_1689);
nand U1976 (N_1976,N_760,In_1036);
nor U1977 (N_1977,N_1604,In_1674);
xnor U1978 (N_1978,In_207,In_145);
and U1979 (N_1979,N_1221,N_809);
or U1980 (N_1980,N_1253,N_1214);
or U1981 (N_1981,In_2104,In_2730);
xnor U1982 (N_1982,In_1974,In_160);
xor U1983 (N_1983,N_585,N_1596);
nand U1984 (N_1984,N_40,N_146);
xor U1985 (N_1985,N_489,N_1719);
and U1986 (N_1986,N_1619,In_2521);
nand U1987 (N_1987,N_1399,N_1607);
nand U1988 (N_1988,N_1708,N_1388);
or U1989 (N_1989,N_1178,N_1584);
or U1990 (N_1990,N_1718,N_1243);
or U1991 (N_1991,N_1778,In_2775);
or U1992 (N_1992,N_1504,N_296);
and U1993 (N_1993,N_419,In_2663);
and U1994 (N_1994,N_1177,N_903);
and U1995 (N_1995,In_2047,N_1141);
nor U1996 (N_1996,N_565,In_296);
or U1997 (N_1997,N_1287,In_2196);
or U1998 (N_1998,In_1737,N_701);
nand U1999 (N_1999,N_1108,N_1356);
and U2000 (N_2000,In_1814,N_1104);
nand U2001 (N_2001,N_1429,N_1323);
or U2002 (N_2002,N_1322,In_131);
xor U2003 (N_2003,N_1552,N_1549);
or U2004 (N_2004,N_389,N_1508);
nand U2005 (N_2005,In_2227,In_905);
nand U2006 (N_2006,In_2925,N_905);
xnor U2007 (N_2007,N_1099,N_772);
and U2008 (N_2008,In_2706,N_1226);
and U2009 (N_2009,In_1200,N_894);
nand U2010 (N_2010,In_2933,In_2477);
nor U2011 (N_2011,In_1557,In_899);
xor U2012 (N_2012,N_1075,N_1290);
nor U2013 (N_2013,N_745,In_2676);
xnor U2014 (N_2014,N_1037,N_1327);
nand U2015 (N_2015,N_1081,In_464);
and U2016 (N_2016,In_326,N_1414);
or U2017 (N_2017,N_1511,N_1298);
or U2018 (N_2018,N_1168,In_1151);
or U2019 (N_2019,N_1472,N_581);
nor U2020 (N_2020,N_1403,N_795);
xor U2021 (N_2021,In_1536,N_1339);
or U2022 (N_2022,N_1609,In_442);
nand U2023 (N_2023,N_1759,N_1312);
nor U2024 (N_2024,N_1559,N_1649);
or U2025 (N_2025,In_777,In_1131);
and U2026 (N_2026,N_1468,N_909);
nand U2027 (N_2027,In_357,In_2502);
or U2028 (N_2028,In_983,In_2728);
xnor U2029 (N_2029,In_929,In_1575);
nand U2030 (N_2030,N_1434,N_1784);
nor U2031 (N_2031,N_901,In_1094);
or U2032 (N_2032,N_1240,N_1579);
or U2033 (N_2033,N_723,In_774);
and U2034 (N_2034,In_441,In_2998);
nand U2035 (N_2035,N_1180,In_2220);
or U2036 (N_2036,N_1701,In_1496);
xnor U2037 (N_2037,N_1088,In_359);
nor U2038 (N_2038,N_1741,N_1608);
xnor U2039 (N_2039,N_1146,N_61);
nand U2040 (N_2040,N_1251,In_1829);
nor U2041 (N_2041,In_2520,N_854);
nor U2042 (N_2042,N_202,N_977);
or U2043 (N_2043,In_743,N_736);
nand U2044 (N_2044,In_2351,N_751);
nor U2045 (N_2045,N_1628,In_545);
and U2046 (N_2046,N_947,N_1769);
xnor U2047 (N_2047,In_622,N_1038);
and U2048 (N_2048,N_1707,N_1651);
nor U2049 (N_2049,In_868,In_2026);
nor U2050 (N_2050,In_2565,N_1766);
and U2051 (N_2051,In_1533,N_875);
nand U2052 (N_2052,N_1315,N_1285);
nor U2053 (N_2053,N_1735,N_1738);
or U2054 (N_2054,In_347,N_1626);
nand U2055 (N_2055,N_1116,In_1443);
nor U2056 (N_2056,N_1446,In_668);
nor U2057 (N_2057,N_1110,N_673);
or U2058 (N_2058,N_1794,N_886);
or U2059 (N_2059,In_294,N_1497);
nor U2060 (N_2060,N_1776,In_2295);
xor U2061 (N_2061,In_2157,In_597);
or U2062 (N_2062,N_936,N_1788);
and U2063 (N_2063,In_684,In_1680);
nor U2064 (N_2064,N_1764,N_1639);
nand U2065 (N_2065,N_1188,N_1737);
xnor U2066 (N_2066,N_1233,In_2609);
nand U2067 (N_2067,N_367,In_1757);
xnor U2068 (N_2068,N_1537,In_883);
xor U2069 (N_2069,N_891,In_1333);
or U2070 (N_2070,N_811,N_1586);
xnor U2071 (N_2071,N_1453,In_2467);
and U2072 (N_2072,In_8,N_1381);
and U2073 (N_2073,N_1111,N_254);
nor U2074 (N_2074,In_1374,In_1230);
nand U2075 (N_2075,In_222,N_1166);
nor U2076 (N_2076,N_1029,N_1734);
xnor U2077 (N_2077,N_1627,In_2926);
nand U2078 (N_2078,N_829,N_1791);
or U2079 (N_2079,N_1687,N_1395);
nor U2080 (N_2080,N_1724,In_1918);
and U2081 (N_2081,In_869,N_1690);
nor U2082 (N_2082,N_1798,N_1533);
xor U2083 (N_2083,N_1514,In_105);
xnor U2084 (N_2084,N_1490,N_1590);
xor U2085 (N_2085,N_157,N_1219);
and U2086 (N_2086,N_1519,N_968);
and U2087 (N_2087,In_623,N_75);
nand U2088 (N_2088,N_1787,In_2687);
nand U2089 (N_2089,N_1083,In_141);
nor U2090 (N_2090,In_838,N_1748);
xor U2091 (N_2091,In_1501,In_2538);
and U2092 (N_2092,N_1793,In_2783);
and U2093 (N_2093,In_22,N_1379);
nor U2094 (N_2094,In_300,N_1211);
and U2095 (N_2095,In_1671,N_671);
nand U2096 (N_2096,N_1726,N_1625);
or U2097 (N_2097,N_1397,N_1463);
xor U2098 (N_2098,In_1549,In_953);
nor U2099 (N_2099,N_546,In_2625);
nor U2100 (N_2100,N_2073,In_2611);
nand U2101 (N_2101,N_1979,N_927);
xor U2102 (N_2102,N_1126,N_1725);
and U2103 (N_2103,N_1551,N_1558);
or U2104 (N_2104,N_2068,N_1118);
xor U2105 (N_2105,N_39,In_2938);
or U2106 (N_2106,N_1656,N_1384);
nor U2107 (N_2107,In_1867,N_808);
xnor U2108 (N_2108,N_1857,N_2039);
xnor U2109 (N_2109,N_1494,In_1899);
or U2110 (N_2110,In_2089,N_1325);
and U2111 (N_2111,N_978,N_1767);
and U2112 (N_2112,In_1447,N_2071);
nor U2113 (N_2113,N_82,N_1496);
nand U2114 (N_2114,In_950,N_1648);
nor U2115 (N_2115,N_1810,N_731);
and U2116 (N_2116,N_2007,N_1600);
and U2117 (N_2117,N_988,N_2095);
or U2118 (N_2118,N_1796,N_2040);
nand U2119 (N_2119,In_2800,N_1375);
or U2120 (N_2120,N_1860,In_1175);
nor U2121 (N_2121,N_1836,N_908);
or U2122 (N_2122,N_2046,N_1674);
nor U2123 (N_2123,In_1018,In_1892);
nor U2124 (N_2124,In_830,N_1694);
and U2125 (N_2125,N_1640,In_966);
and U2126 (N_2126,In_2529,N_1660);
or U2127 (N_2127,In_604,N_1273);
nor U2128 (N_2128,N_2052,In_1471);
xnor U2129 (N_2129,In_21,N_804);
xnor U2130 (N_2130,N_2028,N_1017);
and U2131 (N_2131,N_2015,In_67);
nand U2132 (N_2132,In_1638,N_540);
or U2133 (N_2133,N_1460,N_1963);
xnor U2134 (N_2134,N_827,N_1459);
or U2135 (N_2135,N_566,N_1829);
or U2136 (N_2136,N_515,N_1659);
and U2137 (N_2137,N_281,N_381);
nand U2138 (N_2138,N_1988,N_1785);
xnor U2139 (N_2139,N_1635,N_1913);
nor U2140 (N_2140,N_2054,N_2080);
and U2141 (N_2141,N_1614,N_1222);
nor U2142 (N_2142,N_1849,N_1321);
or U2143 (N_2143,In_1179,In_487);
nand U2144 (N_2144,In_1733,N_2085);
xor U2145 (N_2145,N_344,N_726);
nand U2146 (N_2146,N_1198,In_1138);
and U2147 (N_2147,N_1936,N_2076);
or U2148 (N_2148,N_1967,N_1458);
nor U2149 (N_2149,N_2032,N_998);
or U2150 (N_2150,N_1872,In_1311);
or U2151 (N_2151,N_995,N_1427);
or U2152 (N_2152,N_895,In_226);
nor U2153 (N_2153,N_1880,N_1279);
nand U2154 (N_2154,In_2396,N_1850);
nor U2155 (N_2155,N_1852,N_1884);
and U2156 (N_2156,N_310,N_1881);
or U2157 (N_2157,N_1991,N_1342);
xnor U2158 (N_2158,In_2302,N_1303);
or U2159 (N_2159,N_2082,N_1771);
xor U2160 (N_2160,N_981,N_1957);
xor U2161 (N_2161,N_1673,In_2765);
and U2162 (N_2162,In_2618,N_752);
nand U2163 (N_2163,N_1770,N_1499);
nand U2164 (N_2164,N_1461,N_1779);
xor U2165 (N_2165,N_2066,N_302);
and U2166 (N_2166,N_2025,N_2014);
xnor U2167 (N_2167,N_1550,In_166);
xnor U2168 (N_2168,N_411,In_814);
or U2169 (N_2169,N_18,N_902);
and U2170 (N_2170,N_1801,N_1680);
xnor U2171 (N_2171,N_1951,N_1874);
nand U2172 (N_2172,N_879,N_191);
and U2173 (N_2173,N_1848,In_783);
or U2174 (N_2174,N_1068,N_1819);
and U2175 (N_2175,N_1652,N_1814);
xor U2176 (N_2176,N_1876,N_1636);
nor U2177 (N_2177,N_1154,N_1696);
nand U2178 (N_2178,N_1924,In_1293);
nand U2179 (N_2179,N_2030,In_1858);
xor U2180 (N_2180,N_600,In_2349);
nand U2181 (N_2181,N_1775,In_221);
nand U2182 (N_2182,In_2702,N_1281);
nor U2183 (N_2183,N_1112,N_1623);
or U2184 (N_2184,N_659,N_1802);
nor U2185 (N_2185,N_1981,N_1263);
or U2186 (N_2186,N_2079,In_1111);
xnor U2187 (N_2187,N_1231,N_1329);
or U2188 (N_2188,In_31,In_1296);
or U2189 (N_2189,N_914,N_1809);
nor U2190 (N_2190,N_1866,N_2061);
nand U2191 (N_2191,In_923,N_1272);
nand U2192 (N_2192,N_1820,N_1896);
nor U2193 (N_2193,N_343,N_1825);
and U2194 (N_2194,N_1823,N_1374);
nand U2195 (N_2195,N_1982,N_907);
xnor U2196 (N_2196,N_1833,N_1846);
nand U2197 (N_2197,N_349,N_954);
nand U2198 (N_2198,In_977,N_1276);
nor U2199 (N_2199,N_2059,N_1670);
or U2200 (N_2200,In_2652,N_1544);
or U2201 (N_2201,N_1869,N_1683);
and U2202 (N_2202,In_1630,N_488);
xnor U2203 (N_2203,N_1618,N_1736);
and U2204 (N_2204,N_1937,N_1727);
and U2205 (N_2205,In_2581,N_2055);
nor U2206 (N_2206,N_1464,N_1827);
and U2207 (N_2207,N_1418,In_2844);
and U2208 (N_2208,N_958,N_1818);
nand U2209 (N_2209,N_1261,N_1492);
and U2210 (N_2210,In_1204,N_1839);
nor U2211 (N_2211,N_1202,In_2649);
or U2212 (N_2212,N_482,N_1944);
nor U2213 (N_2213,N_1667,In_385);
or U2214 (N_2214,N_1096,N_1757);
and U2215 (N_2215,N_1079,N_2008);
xor U2216 (N_2216,In_64,In_2977);
and U2217 (N_2217,In_932,N_404);
or U2218 (N_2218,In_1137,N_1977);
or U2219 (N_2219,N_1830,In_1578);
nand U2220 (N_2220,N_780,N_962);
nand U2221 (N_2221,N_784,N_2044);
or U2222 (N_2222,N_2057,N_1700);
or U2223 (N_2223,N_1250,N_231);
nand U2224 (N_2224,N_1939,N_944);
or U2225 (N_2225,N_1699,In_1395);
nand U2226 (N_2226,N_2093,N_1506);
xnor U2227 (N_2227,N_2096,N_1307);
or U2228 (N_2228,N_1863,N_2091);
nor U2229 (N_2229,In_2003,N_766);
nor U2230 (N_2230,N_37,N_612);
xor U2231 (N_2231,N_1897,N_1449);
or U2232 (N_2232,N_1862,In_1852);
nand U2233 (N_2233,N_1915,In_567);
or U2234 (N_2234,N_1973,N_2023);
or U2235 (N_2235,In_2419,N_1016);
xnor U2236 (N_2236,N_796,N_1638);
and U2237 (N_2237,N_1515,N_687);
and U2238 (N_2238,N_2094,N_1362);
and U2239 (N_2239,N_2097,N_368);
or U2240 (N_2240,N_1985,N_1509);
nor U2241 (N_2241,In_1033,N_1070);
or U2242 (N_2242,N_137,In_284);
or U2243 (N_2243,N_1894,N_1886);
nand U2244 (N_2244,N_548,N_1838);
xor U2245 (N_2245,In_1815,N_2019);
or U2246 (N_2246,N_2062,N_2029);
and U2247 (N_2247,N_1732,N_1072);
and U2248 (N_2248,N_1573,In_2457);
or U2249 (N_2249,N_1927,In_2063);
nor U2250 (N_2250,N_1572,N_258);
or U2251 (N_2251,N_773,N_1882);
and U2252 (N_2252,N_1965,N_1918);
or U2253 (N_2253,In_806,N_1995);
nor U2254 (N_2254,N_692,N_2004);
and U2255 (N_2255,N_2074,N_1502);
nor U2256 (N_2256,N_1865,In_308);
nor U2257 (N_2257,N_1807,N_1624);
nand U2258 (N_2258,N_1925,N_1817);
and U2259 (N_2259,N_1969,In_126);
nand U2260 (N_2260,N_2001,In_1634);
nand U2261 (N_2261,In_1729,N_1763);
or U2262 (N_2262,N_1503,N_1834);
nand U2263 (N_2263,In_785,N_1980);
xnor U2264 (N_2264,In_2185,N_1292);
and U2265 (N_2265,In_2570,N_1761);
nor U2266 (N_2266,N_1945,In_2278);
or U2267 (N_2267,N_2060,N_1885);
or U2268 (N_2268,N_2009,N_1943);
xor U2269 (N_2269,N_1956,N_1723);
or U2270 (N_2270,In_2252,N_2099);
nand U2271 (N_2271,In_709,In_1845);
nand U2272 (N_2272,N_1679,N_1976);
nor U2273 (N_2273,In_581,N_2049);
nand U2274 (N_2274,N_1113,In_1424);
xnor U2275 (N_2275,N_1873,N_462);
xor U2276 (N_2276,In_526,N_1302);
xnor U2277 (N_2277,N_1642,N_2067);
nand U2278 (N_2278,N_1946,N_1744);
nor U2279 (N_2279,N_1489,N_2065);
and U2280 (N_2280,N_1824,N_1917);
nor U2281 (N_2281,N_1196,N_1641);
or U2282 (N_2282,In_1948,In_2856);
or U2283 (N_2283,N_2048,N_1716);
nor U2284 (N_2284,N_699,N_1358);
nand U2285 (N_2285,N_1938,In_1493);
nand U2286 (N_2286,N_1611,N_1230);
nor U2287 (N_2287,N_1828,N_1803);
or U2288 (N_2288,N_2006,N_1539);
xnor U2289 (N_2289,In_2966,N_2064);
xnor U2290 (N_2290,N_1001,N_477);
nor U2291 (N_2291,N_1653,N_1546);
and U2292 (N_2292,In_499,N_1161);
and U2293 (N_2293,N_1904,N_1854);
and U2294 (N_2294,N_1756,N_1815);
and U2295 (N_2295,N_651,N_1059);
nand U2296 (N_2296,N_810,N_2013);
and U2297 (N_2297,N_1002,N_1940);
and U2298 (N_2298,N_2083,N_2018);
nor U2299 (N_2299,N_1545,N_1835);
nand U2300 (N_2300,N_319,In_312);
nand U2301 (N_2301,N_1286,N_1970);
xor U2302 (N_2302,N_1650,N_1864);
nand U2303 (N_2303,N_1657,N_2024);
nand U2304 (N_2304,N_604,In_2309);
nor U2305 (N_2305,In_340,N_1950);
or U2306 (N_2306,N_340,N_2063);
nor U2307 (N_2307,N_1432,N_333);
or U2308 (N_2308,N_1971,N_1587);
nor U2309 (N_2309,In_1747,N_516);
or U2310 (N_2310,N_1500,N_1984);
or U2311 (N_2311,N_1954,In_2541);
or U2312 (N_2312,N_1348,N_1603);
xnor U2313 (N_2313,N_929,N_587);
nor U2314 (N_2314,N_1837,In_1776);
nand U2315 (N_2315,N_2078,N_969);
xor U2316 (N_2316,N_714,N_1480);
and U2317 (N_2317,N_1102,N_1958);
nor U2318 (N_2318,N_1968,N_1693);
nand U2319 (N_2319,N_1930,N_1664);
nor U2320 (N_2320,N_940,N_1498);
nand U2321 (N_2321,N_1868,N_1540);
nand U2322 (N_2322,N_1821,N_904);
nor U2323 (N_2323,N_1373,In_2428);
xnor U2324 (N_2324,N_2033,N_1994);
nor U2325 (N_2325,N_1258,N_1754);
or U2326 (N_2326,N_1871,In_43);
and U2327 (N_2327,N_1928,N_2000);
xor U2328 (N_2328,N_1174,N_1346);
and U2329 (N_2329,N_1332,N_1826);
and U2330 (N_2330,N_584,In_1788);
or U2331 (N_2331,N_1349,N_1856);
nand U2332 (N_2332,N_2003,In_2907);
or U2333 (N_2333,N_1935,N_1901);
and U2334 (N_2334,N_729,In_2475);
xnor U2335 (N_2335,N_227,In_2839);
nor U2336 (N_2336,N_642,In_1764);
nor U2337 (N_2337,N_1228,N_1646);
xnor U2338 (N_2338,N_1905,N_1853);
or U2339 (N_2339,N_1909,N_1920);
nor U2340 (N_2340,N_1186,N_1989);
xor U2341 (N_2341,N_1780,In_1312);
or U2342 (N_2342,N_247,N_1267);
or U2343 (N_2343,N_1575,N_1520);
or U2344 (N_2344,In_1971,In_1981);
nand U2345 (N_2345,N_1998,N_1340);
nand U2346 (N_2346,In_1560,N_1621);
nand U2347 (N_2347,In_24,In_850);
or U2348 (N_2348,In_2373,N_1952);
or U2349 (N_2349,N_1071,N_1278);
nand U2350 (N_2350,N_1753,N_475);
nand U2351 (N_2351,N_1858,N_778);
and U2352 (N_2352,N_1630,N_1531);
nor U2353 (N_2353,N_999,N_1382);
xnor U2354 (N_2354,In_1683,N_1879);
and U2355 (N_2355,In_2864,N_1602);
nor U2356 (N_2356,In_1240,N_960);
and U2357 (N_2357,N_558,N_242);
nand U2358 (N_2358,N_1678,N_1383);
nor U2359 (N_2359,N_2086,N_1996);
xnor U2360 (N_2360,N_2045,In_1759);
and U2361 (N_2361,N_2092,N_1986);
nand U2362 (N_2362,N_869,N_1595);
and U2363 (N_2363,In_1625,N_1746);
and U2364 (N_2364,N_1773,N_1036);
xor U2365 (N_2365,N_1934,In_1423);
and U2366 (N_2366,In_2953,N_966);
nand U2367 (N_2367,In_2904,N_1566);
nor U2368 (N_2368,N_1283,N_1842);
nand U2369 (N_2369,N_2012,N_1591);
nand U2370 (N_2370,N_1523,N_646);
and U2371 (N_2371,N_0,N_1633);
nand U2372 (N_2372,N_1175,N_866);
nor U2373 (N_2373,N_757,In_2712);
xnor U2374 (N_2374,N_1599,In_1778);
nor U2375 (N_2375,In_2587,N_1911);
or U2376 (N_2376,N_1922,N_1789);
and U2377 (N_2377,In_1182,N_1218);
nor U2378 (N_2378,N_1561,N_1800);
and U2379 (N_2379,In_725,N_623);
nor U2380 (N_2380,N_1870,N_420);
xnor U2381 (N_2381,N_2081,N_1655);
nand U2382 (N_2382,N_1526,N_818);
nand U2383 (N_2383,N_1265,N_1220);
nor U2384 (N_2384,N_408,N_1548);
nor U2385 (N_2385,N_1990,In_2077);
nor U2386 (N_2386,N_1105,In_1833);
nor U2387 (N_2387,N_1831,N_1743);
or U2388 (N_2388,N_965,In_2778);
nand U2389 (N_2389,N_1961,N_987);
xnor U2390 (N_2390,N_1236,N_423);
and U2391 (N_2391,In_986,N_1855);
or U2392 (N_2392,N_1875,In_2128);
xnor U2393 (N_2393,N_498,In_444);
and U2394 (N_2394,N_1505,In_1544);
nand U2395 (N_2395,N_1953,N_1522);
or U2396 (N_2396,N_2084,N_1889);
and U2397 (N_2397,N_1919,In_2771);
and U2398 (N_2398,In_1061,N_1247);
or U2399 (N_2399,N_1847,N_384);
xor U2400 (N_2400,N_1491,N_2206);
or U2401 (N_2401,N_2121,N_2192);
and U2402 (N_2402,N_1728,N_1742);
nor U2403 (N_2403,N_2297,N_2141);
or U2404 (N_2404,N_1813,N_2285);
or U2405 (N_2405,N_2201,N_2243);
or U2406 (N_2406,N_1299,N_2198);
or U2407 (N_2407,N_2363,N_2356);
nor U2408 (N_2408,N_2299,N_2209);
or U2409 (N_2409,N_705,N_1916);
or U2410 (N_2410,N_2252,N_2050);
and U2411 (N_2411,N_2186,N_1430);
xnor U2412 (N_2412,N_2290,N_2005);
and U2413 (N_2413,In_2189,N_2163);
nor U2414 (N_2414,N_2332,N_2233);
or U2415 (N_2415,N_430,N_2341);
xor U2416 (N_2416,N_2237,N_1974);
or U2417 (N_2417,N_1661,In_1559);
nand U2418 (N_2418,N_2282,N_2118);
nand U2419 (N_2419,N_2165,N_2178);
and U2420 (N_2420,N_2017,N_2392);
or U2421 (N_2421,N_1975,N_2292);
nor U2422 (N_2422,N_1074,N_1333);
nor U2423 (N_2423,N_1903,N_1812);
or U2424 (N_2424,N_2034,N_2120);
nor U2425 (N_2425,N_1164,N_1400);
and U2426 (N_2426,In_2803,In_1809);
nor U2427 (N_2427,N_2182,N_2344);
or U2428 (N_2428,N_2245,N_856);
or U2429 (N_2429,N_2300,N_2254);
xor U2430 (N_2430,N_2230,N_2368);
and U2431 (N_2431,N_2360,N_1805);
xor U2432 (N_2432,N_1808,N_2139);
or U2433 (N_2433,N_2333,N_2247);
nor U2434 (N_2434,N_2231,N_611);
or U2435 (N_2435,N_1893,N_1581);
nand U2436 (N_2436,N_1900,N_2106);
nor U2437 (N_2437,N_2278,N_2047);
or U2438 (N_2438,N_1843,N_1513);
xor U2439 (N_2439,N_1811,N_1999);
and U2440 (N_2440,N_2365,N_2132);
nand U2441 (N_2441,N_2124,N_1610);
nand U2442 (N_2442,N_2397,N_1185);
nor U2443 (N_2443,N_2327,N_2378);
xnor U2444 (N_2444,N_1467,N_2335);
or U2445 (N_2445,N_1698,N_1049);
xnor U2446 (N_2446,N_393,In_2994);
nor U2447 (N_2447,N_2339,N_1790);
xnor U2448 (N_2448,N_2102,N_2375);
or U2449 (N_2449,N_1334,In_27);
nor U2450 (N_2450,N_356,N_1293);
or U2451 (N_2451,N_2051,N_1822);
and U2452 (N_2452,N_1365,N_2340);
nand U2453 (N_2453,N_2196,N_1923);
nor U2454 (N_2454,N_1906,N_1841);
or U2455 (N_2455,In_2231,N_2373);
nor U2456 (N_2456,In_2240,N_2119);
nor U2457 (N_2457,N_2353,N_754);
or U2458 (N_2458,In_1062,N_2343);
and U2459 (N_2459,N_1992,N_1421);
or U2460 (N_2460,N_1571,In_2114);
or U2461 (N_2461,N_2330,In_865);
nor U2462 (N_2462,N_608,N_1851);
or U2463 (N_2463,N_2275,N_2153);
nor U2464 (N_2464,N_1926,N_1306);
nand U2465 (N_2465,N_2383,N_1721);
nand U2466 (N_2466,N_1959,N_2324);
xnor U2467 (N_2467,N_1574,N_1931);
or U2468 (N_2468,N_1942,N_2323);
xnor U2469 (N_2469,N_320,N_2200);
nand U2470 (N_2470,N_1510,N_2157);
nor U2471 (N_2471,N_2281,N_2114);
xnor U2472 (N_2472,N_2122,N_2152);
nor U2473 (N_2473,In_1880,N_2100);
xor U2474 (N_2474,N_2312,N_2123);
nand U2475 (N_2475,N_2160,N_2239);
and U2476 (N_2476,N_2117,N_2225);
and U2477 (N_2477,N_2125,In_833);
and U2478 (N_2478,N_2257,In_1862);
nand U2479 (N_2479,N_2269,N_2177);
nand U2480 (N_2480,N_2264,N_2204);
or U2481 (N_2481,N_1844,N_2002);
nor U2482 (N_2482,N_2352,N_2270);
nor U2483 (N_2483,In_189,In_1589);
or U2484 (N_2484,N_1473,N_2384);
nor U2485 (N_2485,N_2294,N_2035);
or U2486 (N_2486,N_2176,N_2208);
xnor U2487 (N_2487,N_2321,N_2334);
or U2488 (N_2488,N_2205,N_2190);
nor U2489 (N_2489,N_1532,N_1711);
or U2490 (N_2490,N_2164,N_2109);
nand U2491 (N_2491,N_2135,N_472);
or U2492 (N_2492,N_2161,N_2380);
and U2493 (N_2493,N_871,N_1715);
and U2494 (N_2494,N_1731,N_1964);
nand U2495 (N_2495,N_2315,N_1883);
xnor U2496 (N_2496,N_2170,N_2213);
nor U2497 (N_2497,N_1898,N_164);
xor U2498 (N_2498,N_1997,N_2336);
xor U2499 (N_2499,N_2219,N_2215);
xnor U2500 (N_2500,N_2179,In_1122);
or U2501 (N_2501,N_1702,In_2423);
and U2502 (N_2502,N_2207,N_2156);
xnor U2503 (N_2503,N_1949,N_1528);
xnor U2504 (N_2504,N_1816,N_2295);
and U2505 (N_2505,N_2151,N_653);
xnor U2506 (N_2506,In_52,N_2279);
and U2507 (N_2507,N_1962,N_2288);
xnor U2508 (N_2508,N_2370,In_1027);
and U2509 (N_2509,N_2016,N_2056);
nand U2510 (N_2510,In_1770,N_2173);
nand U2511 (N_2511,N_2347,N_2385);
xnor U2512 (N_2512,In_2646,N_619);
nor U2513 (N_2513,N_2202,In_2954);
and U2514 (N_2514,N_2262,N_1933);
or U2515 (N_2515,N_2296,N_1582);
or U2516 (N_2516,In_947,N_1758);
xnor U2517 (N_2517,N_1912,N_1966);
xnor U2518 (N_2518,N_2326,N_2342);
and U2519 (N_2519,N_2221,N_2116);
nor U2520 (N_2520,N_2162,In_127);
or U2521 (N_2521,N_2372,N_2246);
nor U2522 (N_2522,In_2030,N_1891);
nand U2523 (N_2523,N_1376,N_2218);
nand U2524 (N_2524,N_2187,N_1170);
nor U2525 (N_2525,N_1914,N_2355);
nor U2526 (N_2526,In_1772,N_2238);
or U2527 (N_2527,N_2301,N_1832);
and U2528 (N_2528,N_614,N_755);
and U2529 (N_2529,N_2235,N_2236);
xor U2530 (N_2530,N_2174,N_1255);
nand U2531 (N_2531,N_2346,In_41);
xor U2532 (N_2532,N_2189,N_2133);
nor U2533 (N_2533,N_2037,N_2226);
xnor U2534 (N_2534,N_2129,In_931);
or U2535 (N_2535,N_2302,N_2199);
nor U2536 (N_2536,N_2223,N_1668);
xnor U2537 (N_2537,N_1972,N_2331);
xnor U2538 (N_2538,N_2389,In_270);
and U2539 (N_2539,N_2140,N_1840);
or U2540 (N_2540,N_2195,In_2859);
and U2541 (N_2541,N_2090,N_1556);
nand U2542 (N_2542,N_991,N_1932);
nand U2543 (N_2543,N_2126,N_1662);
and U2544 (N_2544,N_2234,N_2088);
nand U2545 (N_2545,N_2276,N_1518);
nor U2546 (N_2546,N_2318,N_2131);
nor U2547 (N_2547,N_1555,N_2166);
or U2548 (N_2548,N_1908,N_1983);
nor U2549 (N_2549,N_2366,N_2266);
nand U2550 (N_2550,N_1729,N_1671);
and U2551 (N_2551,N_2185,N_363);
nand U2552 (N_2552,N_1525,N_1772);
nand U2553 (N_2553,N_2304,N_1692);
and U2554 (N_2554,N_2255,N_2111);
or U2555 (N_2555,N_2210,N_1423);
nand U2556 (N_2556,N_2329,N_2113);
xnor U2557 (N_2557,N_1613,N_2142);
nor U2558 (N_2558,N_2357,N_2379);
xnor U2559 (N_2559,N_1907,N_2042);
xnor U2560 (N_2560,N_2112,N_2354);
nor U2561 (N_2561,N_1569,N_1601);
and U2562 (N_2562,In_498,N_1053);
or U2563 (N_2563,N_336,N_1697);
xor U2564 (N_2564,N_2211,N_2313);
and U2565 (N_2565,In_2511,N_2229);
nand U2566 (N_2566,N_1978,N_2289);
and U2567 (N_2567,N_2038,In_1239);
nor U2568 (N_2568,N_1797,N_2228);
and U2569 (N_2569,N_763,N_1205);
xor U2570 (N_2570,N_1355,N_2350);
nor U2571 (N_2571,N_2359,N_1201);
nor U2572 (N_2572,In_2073,N_1745);
xor U2573 (N_2573,N_2271,N_2031);
xnor U2574 (N_2574,N_989,N_2053);
or U2575 (N_2575,N_2159,N_2169);
or U2576 (N_2576,N_2272,In_2365);
or U2577 (N_2577,N_2317,N_2303);
nor U2578 (N_2578,N_2058,N_364);
nand U2579 (N_2579,N_2130,N_2259);
nand U2580 (N_2580,N_1760,N_2098);
nand U2581 (N_2581,N_982,N_2386);
or U2582 (N_2582,N_2175,N_1411);
xor U2583 (N_2583,In_1730,N_2267);
nand U2584 (N_2584,N_1895,N_2087);
and U2585 (N_2585,N_2381,N_746);
or U2586 (N_2586,N_1888,N_2308);
and U2587 (N_2587,In_283,N_2149);
xnor U2588 (N_2588,N_2021,N_1948);
and U2589 (N_2589,N_354,N_2137);
xor U2590 (N_2590,N_1921,N_1367);
or U2591 (N_2591,N_1714,N_2367);
nand U2592 (N_2592,N_2168,N_2222);
nor U2593 (N_2593,N_2250,N_2136);
nand U2594 (N_2594,N_712,N_2184);
nor U2595 (N_2595,N_2319,N_2358);
or U2596 (N_2596,N_2286,N_1941);
or U2597 (N_2597,N_1199,N_2128);
and U2598 (N_2598,N_2345,N_1634);
nand U2599 (N_2599,N_1131,N_144);
xor U2600 (N_2600,N_274,N_2284);
xor U2601 (N_2601,N_2027,N_2077);
nor U2602 (N_2602,N_1622,N_1993);
xor U2603 (N_2603,N_1899,In_1431);
or U2604 (N_2604,N_1501,N_2311);
nor U2605 (N_2605,N_1593,N_2306);
and U2606 (N_2606,N_2146,N_2348);
xnor U2607 (N_2607,N_2349,N_2396);
nand U2608 (N_2608,N_2216,N_2010);
xnor U2609 (N_2609,N_2020,In_2729);
and U2610 (N_2610,N_1023,N_2307);
and U2611 (N_2611,N_1765,In_1047);
xnor U2612 (N_2612,N_2232,N_2265);
xnor U2613 (N_2613,N_2110,N_1867);
nand U2614 (N_2614,N_2217,N_2104);
nor U2615 (N_2615,N_2180,N_2171);
or U2616 (N_2616,N_1476,In_345);
nand U2617 (N_2617,N_2183,In_2993);
or U2618 (N_2618,N_2154,N_2398);
nand U2619 (N_2619,In_2563,N_1553);
or U2620 (N_2620,In_2700,N_2158);
and U2621 (N_2621,N_2188,N_1193);
xor U2622 (N_2622,N_1890,N_127);
and U2623 (N_2623,N_2022,N_2393);
nand U2624 (N_2624,N_2144,N_2399);
and U2625 (N_2625,N_2382,N_2328);
nand U2626 (N_2626,In_1939,N_2320);
nor U2627 (N_2627,N_1887,N_2291);
or U2628 (N_2628,N_1378,N_1097);
nor U2629 (N_2629,In_1846,N_2274);
nor U2630 (N_2630,N_1878,N_2394);
or U2631 (N_2631,N_2337,N_2101);
or U2632 (N_2632,N_2145,In_2569);
nand U2633 (N_2633,N_2212,N_1495);
xnor U2634 (N_2634,N_2361,N_2376);
nand U2635 (N_2635,N_2241,N_2224);
xor U2636 (N_2636,N_2167,N_1363);
or U2637 (N_2637,In_2406,N_2369);
nand U2638 (N_2638,N_2075,N_2127);
or U2639 (N_2639,N_2310,N_1877);
or U2640 (N_2640,N_2220,N_414);
xnor U2641 (N_2641,N_2043,N_2107);
nand U2642 (N_2642,N_2293,N_2362);
or U2643 (N_2643,N_1564,N_2374);
xnor U2644 (N_2644,N_2143,N_2388);
and U2645 (N_2645,N_2214,N_2248);
nand U2646 (N_2646,In_786,In_2794);
and U2647 (N_2647,N_2273,N_2138);
xor U2648 (N_2648,N_2072,N_1259);
nor U2649 (N_2649,N_1456,In_1749);
nand U2650 (N_2650,N_2240,N_2011);
and U2651 (N_2651,N_1133,N_1861);
xor U2652 (N_2652,In_558,N_2105);
nand U2653 (N_2653,N_1892,N_2242);
nor U2654 (N_2654,N_1781,In_916);
and U2655 (N_2655,N_1018,N_2193);
xor U2656 (N_2656,N_2115,N_2377);
xnor U2657 (N_2657,In_2265,N_2041);
nand U2658 (N_2658,N_2181,N_2325);
nand U2659 (N_2659,N_170,N_2134);
and U2660 (N_2660,N_2026,N_2287);
nor U2661 (N_2661,N_2227,N_1658);
nand U2662 (N_2662,N_2263,N_2197);
and U2663 (N_2663,N_1777,N_1845);
and U2664 (N_2664,N_2089,N_2261);
nor U2665 (N_2665,N_2249,N_1451);
and U2666 (N_2666,N_2316,N_1910);
nand U2667 (N_2667,N_2322,N_2305);
or U2668 (N_2668,N_2298,N_2148);
or U2669 (N_2669,N_2391,N_2351);
or U2670 (N_2670,In_2860,N_1751);
and U2671 (N_2671,N_2108,N_2147);
and U2672 (N_2672,N_2260,In_2891);
nand U2673 (N_2673,N_2251,N_19);
or U2674 (N_2674,N_2172,N_1806);
nor U2675 (N_2675,N_1371,N_232);
xnor U2676 (N_2676,N_2280,N_2194);
and U2677 (N_2677,N_1987,N_2395);
and U2678 (N_2678,N_2036,N_2364);
and U2679 (N_2679,In_310,N_1441);
and U2680 (N_2680,N_2371,N_2268);
or U2681 (N_2681,N_572,N_1955);
and U2682 (N_2682,N_2203,N_2258);
xnor U2683 (N_2683,N_2387,N_1902);
nor U2684 (N_2684,N_2283,N_1929);
nand U2685 (N_2685,N_2390,N_1804);
nand U2686 (N_2686,N_2191,In_324);
nand U2687 (N_2687,N_1486,N_952);
and U2688 (N_2688,N_1947,N_1438);
xor U2689 (N_2689,In_1834,N_2277);
xnor U2690 (N_2690,N_2155,N_1064);
xor U2691 (N_2691,N_536,N_1960);
nor U2692 (N_2692,N_2103,N_1440);
nor U2693 (N_2693,N_2256,N_1277);
and U2694 (N_2694,N_2314,N_542);
nand U2695 (N_2695,N_1632,N_2253);
or U2696 (N_2696,N_2070,N_2069);
and U2697 (N_2697,N_2338,N_2244);
xnor U2698 (N_2698,N_2309,N_1859);
xnor U2699 (N_2699,N_2150,N_1527);
nand U2700 (N_2700,N_2497,N_2499);
xor U2701 (N_2701,N_2430,N_2574);
xnor U2702 (N_2702,N_2498,N_2519);
nor U2703 (N_2703,N_2596,N_2484);
nand U2704 (N_2704,N_2661,N_2545);
or U2705 (N_2705,N_2567,N_2544);
and U2706 (N_2706,N_2621,N_2694);
and U2707 (N_2707,N_2415,N_2464);
nor U2708 (N_2708,N_2500,N_2440);
and U2709 (N_2709,N_2659,N_2495);
and U2710 (N_2710,N_2413,N_2429);
nand U2711 (N_2711,N_2691,N_2663);
xnor U2712 (N_2712,N_2487,N_2425);
and U2713 (N_2713,N_2409,N_2630);
xor U2714 (N_2714,N_2629,N_2411);
xor U2715 (N_2715,N_2428,N_2623);
and U2716 (N_2716,N_2472,N_2591);
or U2717 (N_2717,N_2664,N_2465);
nor U2718 (N_2718,N_2676,N_2521);
or U2719 (N_2719,N_2426,N_2656);
or U2720 (N_2720,N_2699,N_2561);
nand U2721 (N_2721,N_2575,N_2577);
and U2722 (N_2722,N_2622,N_2618);
nand U2723 (N_2723,N_2654,N_2400);
xnor U2724 (N_2724,N_2626,N_2452);
nor U2725 (N_2725,N_2640,N_2616);
and U2726 (N_2726,N_2491,N_2447);
xor U2727 (N_2727,N_2653,N_2463);
and U2728 (N_2728,N_2459,N_2693);
and U2729 (N_2729,N_2683,N_2688);
xnor U2730 (N_2730,N_2668,N_2414);
or U2731 (N_2731,N_2603,N_2520);
xor U2732 (N_2732,N_2407,N_2535);
or U2733 (N_2733,N_2681,N_2692);
nor U2734 (N_2734,N_2438,N_2560);
and U2735 (N_2735,N_2635,N_2558);
nor U2736 (N_2736,N_2476,N_2601);
and U2737 (N_2737,N_2402,N_2532);
nor U2738 (N_2738,N_2550,N_2581);
and U2739 (N_2739,N_2446,N_2537);
or U2740 (N_2740,N_2605,N_2647);
nand U2741 (N_2741,N_2408,N_2412);
or U2742 (N_2742,N_2637,N_2493);
xnor U2743 (N_2743,N_2424,N_2516);
xor U2744 (N_2744,N_2580,N_2613);
and U2745 (N_2745,N_2417,N_2434);
nor U2746 (N_2746,N_2582,N_2564);
nand U2747 (N_2747,N_2517,N_2671);
nor U2748 (N_2748,N_2492,N_2526);
or U2749 (N_2749,N_2557,N_2529);
and U2750 (N_2750,N_2538,N_2536);
or U2751 (N_2751,N_2505,N_2488);
xnor U2752 (N_2752,N_2543,N_2509);
nand U2753 (N_2753,N_2482,N_2477);
xor U2754 (N_2754,N_2607,N_2416);
nand U2755 (N_2755,N_2590,N_2669);
nand U2756 (N_2756,N_2523,N_2658);
and U2757 (N_2757,N_2540,N_2609);
xor U2758 (N_2758,N_2643,N_2566);
nand U2759 (N_2759,N_2649,N_2507);
nand U2760 (N_2760,N_2627,N_2436);
and U2761 (N_2761,N_2510,N_2645);
nand U2762 (N_2762,N_2443,N_2650);
and U2763 (N_2763,N_2644,N_2453);
and U2764 (N_2764,N_2524,N_2620);
nor U2765 (N_2765,N_2527,N_2485);
or U2766 (N_2766,N_2614,N_2502);
or U2767 (N_2767,N_2468,N_2432);
nand U2768 (N_2768,N_2617,N_2471);
or U2769 (N_2769,N_2625,N_2602);
xnor U2770 (N_2770,N_2454,N_2652);
nor U2771 (N_2771,N_2592,N_2587);
or U2772 (N_2772,N_2585,N_2483);
xnor U2773 (N_2773,N_2682,N_2486);
nor U2774 (N_2774,N_2554,N_2615);
and U2775 (N_2775,N_2501,N_2563);
nor U2776 (N_2776,N_2503,N_2455);
and U2777 (N_2777,N_2667,N_2462);
nand U2778 (N_2778,N_2642,N_2405);
xnor U2779 (N_2779,N_2695,N_2619);
or U2780 (N_2780,N_2628,N_2677);
or U2781 (N_2781,N_2457,N_2588);
xor U2782 (N_2782,N_2406,N_2624);
or U2783 (N_2783,N_2441,N_2696);
or U2784 (N_2784,N_2646,N_2690);
xnor U2785 (N_2785,N_2697,N_2480);
nand U2786 (N_2786,N_2546,N_2641);
or U2787 (N_2787,N_2684,N_2420);
nor U2788 (N_2788,N_2513,N_2444);
nor U2789 (N_2789,N_2565,N_2660);
or U2790 (N_2790,N_2490,N_2439);
nand U2791 (N_2791,N_2583,N_2633);
or U2792 (N_2792,N_2638,N_2665);
xor U2793 (N_2793,N_2572,N_2552);
and U2794 (N_2794,N_2674,N_2456);
nand U2795 (N_2795,N_2608,N_2458);
nor U2796 (N_2796,N_2651,N_2598);
or U2797 (N_2797,N_2422,N_2541);
nor U2798 (N_2798,N_2481,N_2573);
xor U2799 (N_2799,N_2556,N_2686);
nor U2800 (N_2800,N_2419,N_2512);
nand U2801 (N_2801,N_2451,N_2600);
nand U2802 (N_2802,N_2449,N_2533);
nor U2803 (N_2803,N_2442,N_2494);
nand U2804 (N_2804,N_2473,N_2469);
nand U2805 (N_2805,N_2648,N_2612);
or U2806 (N_2806,N_2662,N_2539);
nor U2807 (N_2807,N_2534,N_2479);
and U2808 (N_2808,N_2531,N_2655);
nand U2809 (N_2809,N_2673,N_2639);
xnor U2810 (N_2810,N_2470,N_2670);
nor U2811 (N_2811,N_2403,N_2549);
nand U2812 (N_2812,N_2597,N_2489);
or U2813 (N_2813,N_2461,N_2698);
nand U2814 (N_2814,N_2672,N_2421);
or U2815 (N_2815,N_2599,N_2448);
or U2816 (N_2816,N_2460,N_2576);
and U2817 (N_2817,N_2548,N_2594);
nor U2818 (N_2818,N_2475,N_2450);
xnor U2819 (N_2819,N_2562,N_2547);
and U2820 (N_2820,N_2437,N_2467);
nor U2821 (N_2821,N_2433,N_2496);
xnor U2822 (N_2822,N_2404,N_2525);
or U2823 (N_2823,N_2570,N_2571);
or U2824 (N_2824,N_2553,N_2687);
nor U2825 (N_2825,N_2542,N_2410);
and U2826 (N_2826,N_2401,N_2689);
or U2827 (N_2827,N_2518,N_2528);
nor U2828 (N_2828,N_2685,N_2504);
and U2829 (N_2829,N_2586,N_2474);
and U2830 (N_2830,N_2431,N_2606);
nand U2831 (N_2831,N_2632,N_2506);
xor U2832 (N_2832,N_2579,N_2522);
or U2833 (N_2833,N_2589,N_2423);
and U2834 (N_2834,N_2551,N_2478);
or U2835 (N_2835,N_2466,N_2555);
nand U2836 (N_2836,N_2530,N_2445);
and U2837 (N_2837,N_2418,N_2435);
and U2838 (N_2838,N_2427,N_2511);
nand U2839 (N_2839,N_2578,N_2666);
or U2840 (N_2840,N_2657,N_2611);
and U2841 (N_2841,N_2569,N_2634);
and U2842 (N_2842,N_2584,N_2675);
and U2843 (N_2843,N_2680,N_2568);
nor U2844 (N_2844,N_2631,N_2514);
or U2845 (N_2845,N_2559,N_2595);
and U2846 (N_2846,N_2679,N_2508);
nor U2847 (N_2847,N_2515,N_2610);
nor U2848 (N_2848,N_2678,N_2604);
nand U2849 (N_2849,N_2636,N_2593);
nor U2850 (N_2850,N_2510,N_2696);
or U2851 (N_2851,N_2510,N_2557);
or U2852 (N_2852,N_2514,N_2583);
xnor U2853 (N_2853,N_2489,N_2408);
and U2854 (N_2854,N_2457,N_2614);
nor U2855 (N_2855,N_2556,N_2521);
and U2856 (N_2856,N_2413,N_2549);
nand U2857 (N_2857,N_2457,N_2540);
nor U2858 (N_2858,N_2548,N_2651);
nor U2859 (N_2859,N_2669,N_2432);
and U2860 (N_2860,N_2664,N_2523);
and U2861 (N_2861,N_2481,N_2695);
nor U2862 (N_2862,N_2512,N_2552);
xnor U2863 (N_2863,N_2512,N_2413);
nor U2864 (N_2864,N_2559,N_2546);
xor U2865 (N_2865,N_2680,N_2433);
xnor U2866 (N_2866,N_2690,N_2572);
xor U2867 (N_2867,N_2560,N_2429);
nand U2868 (N_2868,N_2481,N_2433);
nand U2869 (N_2869,N_2572,N_2510);
or U2870 (N_2870,N_2468,N_2482);
xor U2871 (N_2871,N_2444,N_2626);
xnor U2872 (N_2872,N_2586,N_2656);
or U2873 (N_2873,N_2592,N_2672);
xnor U2874 (N_2874,N_2503,N_2459);
and U2875 (N_2875,N_2453,N_2501);
xnor U2876 (N_2876,N_2448,N_2600);
xor U2877 (N_2877,N_2455,N_2466);
and U2878 (N_2878,N_2518,N_2616);
nor U2879 (N_2879,N_2563,N_2553);
nand U2880 (N_2880,N_2486,N_2563);
xor U2881 (N_2881,N_2649,N_2623);
nor U2882 (N_2882,N_2667,N_2529);
and U2883 (N_2883,N_2409,N_2468);
nor U2884 (N_2884,N_2400,N_2463);
xnor U2885 (N_2885,N_2624,N_2483);
and U2886 (N_2886,N_2450,N_2402);
and U2887 (N_2887,N_2452,N_2597);
nand U2888 (N_2888,N_2554,N_2484);
or U2889 (N_2889,N_2505,N_2462);
xnor U2890 (N_2890,N_2514,N_2480);
xnor U2891 (N_2891,N_2469,N_2551);
nand U2892 (N_2892,N_2484,N_2619);
nor U2893 (N_2893,N_2658,N_2473);
nor U2894 (N_2894,N_2578,N_2512);
or U2895 (N_2895,N_2438,N_2643);
xor U2896 (N_2896,N_2601,N_2661);
xnor U2897 (N_2897,N_2443,N_2428);
or U2898 (N_2898,N_2571,N_2614);
nand U2899 (N_2899,N_2502,N_2675);
and U2900 (N_2900,N_2674,N_2687);
xnor U2901 (N_2901,N_2699,N_2483);
or U2902 (N_2902,N_2466,N_2589);
and U2903 (N_2903,N_2642,N_2434);
nor U2904 (N_2904,N_2476,N_2417);
and U2905 (N_2905,N_2692,N_2651);
nand U2906 (N_2906,N_2593,N_2488);
and U2907 (N_2907,N_2474,N_2431);
xor U2908 (N_2908,N_2432,N_2402);
xnor U2909 (N_2909,N_2571,N_2603);
nor U2910 (N_2910,N_2424,N_2421);
nor U2911 (N_2911,N_2578,N_2553);
nand U2912 (N_2912,N_2649,N_2484);
or U2913 (N_2913,N_2698,N_2462);
xnor U2914 (N_2914,N_2620,N_2455);
and U2915 (N_2915,N_2587,N_2664);
and U2916 (N_2916,N_2587,N_2527);
or U2917 (N_2917,N_2551,N_2613);
or U2918 (N_2918,N_2523,N_2650);
xor U2919 (N_2919,N_2460,N_2540);
xnor U2920 (N_2920,N_2677,N_2660);
or U2921 (N_2921,N_2554,N_2681);
or U2922 (N_2922,N_2515,N_2636);
and U2923 (N_2923,N_2522,N_2469);
nand U2924 (N_2924,N_2449,N_2575);
or U2925 (N_2925,N_2638,N_2410);
nor U2926 (N_2926,N_2626,N_2507);
xnor U2927 (N_2927,N_2424,N_2665);
nor U2928 (N_2928,N_2476,N_2490);
nand U2929 (N_2929,N_2698,N_2546);
nand U2930 (N_2930,N_2457,N_2482);
or U2931 (N_2931,N_2408,N_2589);
and U2932 (N_2932,N_2568,N_2429);
nand U2933 (N_2933,N_2446,N_2545);
xnor U2934 (N_2934,N_2486,N_2672);
nand U2935 (N_2935,N_2533,N_2475);
nand U2936 (N_2936,N_2425,N_2635);
and U2937 (N_2937,N_2421,N_2462);
and U2938 (N_2938,N_2599,N_2555);
and U2939 (N_2939,N_2493,N_2508);
xnor U2940 (N_2940,N_2683,N_2536);
nor U2941 (N_2941,N_2629,N_2678);
nor U2942 (N_2942,N_2433,N_2598);
or U2943 (N_2943,N_2607,N_2676);
nor U2944 (N_2944,N_2438,N_2635);
and U2945 (N_2945,N_2609,N_2453);
nor U2946 (N_2946,N_2553,N_2474);
nor U2947 (N_2947,N_2504,N_2577);
nand U2948 (N_2948,N_2591,N_2540);
xor U2949 (N_2949,N_2508,N_2585);
xor U2950 (N_2950,N_2487,N_2620);
and U2951 (N_2951,N_2680,N_2642);
and U2952 (N_2952,N_2666,N_2585);
nor U2953 (N_2953,N_2573,N_2556);
nand U2954 (N_2954,N_2508,N_2527);
nand U2955 (N_2955,N_2440,N_2658);
nor U2956 (N_2956,N_2603,N_2518);
nand U2957 (N_2957,N_2569,N_2633);
nor U2958 (N_2958,N_2517,N_2460);
nand U2959 (N_2959,N_2623,N_2484);
or U2960 (N_2960,N_2699,N_2600);
or U2961 (N_2961,N_2644,N_2510);
or U2962 (N_2962,N_2433,N_2609);
nand U2963 (N_2963,N_2603,N_2537);
xor U2964 (N_2964,N_2639,N_2691);
nand U2965 (N_2965,N_2499,N_2410);
and U2966 (N_2966,N_2648,N_2652);
or U2967 (N_2967,N_2645,N_2652);
xor U2968 (N_2968,N_2410,N_2446);
and U2969 (N_2969,N_2643,N_2693);
nor U2970 (N_2970,N_2642,N_2406);
xnor U2971 (N_2971,N_2491,N_2549);
nor U2972 (N_2972,N_2456,N_2585);
xnor U2973 (N_2973,N_2525,N_2423);
or U2974 (N_2974,N_2465,N_2665);
or U2975 (N_2975,N_2438,N_2585);
and U2976 (N_2976,N_2478,N_2580);
nand U2977 (N_2977,N_2527,N_2433);
or U2978 (N_2978,N_2678,N_2525);
and U2979 (N_2979,N_2452,N_2619);
nand U2980 (N_2980,N_2441,N_2547);
and U2981 (N_2981,N_2498,N_2417);
xnor U2982 (N_2982,N_2598,N_2697);
and U2983 (N_2983,N_2422,N_2674);
xnor U2984 (N_2984,N_2537,N_2498);
xnor U2985 (N_2985,N_2546,N_2570);
nand U2986 (N_2986,N_2661,N_2647);
xor U2987 (N_2987,N_2643,N_2617);
nor U2988 (N_2988,N_2696,N_2570);
or U2989 (N_2989,N_2648,N_2466);
or U2990 (N_2990,N_2662,N_2604);
and U2991 (N_2991,N_2483,N_2416);
and U2992 (N_2992,N_2428,N_2657);
or U2993 (N_2993,N_2455,N_2533);
nand U2994 (N_2994,N_2573,N_2471);
xnor U2995 (N_2995,N_2405,N_2679);
nand U2996 (N_2996,N_2517,N_2611);
and U2997 (N_2997,N_2647,N_2513);
and U2998 (N_2998,N_2686,N_2580);
nand U2999 (N_2999,N_2516,N_2581);
xnor U3000 (N_3000,N_2730,N_2725);
xnor U3001 (N_3001,N_2728,N_2822);
nor U3002 (N_3002,N_2931,N_2857);
or U3003 (N_3003,N_2946,N_2908);
and U3004 (N_3004,N_2731,N_2935);
or U3005 (N_3005,N_2726,N_2939);
nor U3006 (N_3006,N_2945,N_2794);
nand U3007 (N_3007,N_2910,N_2918);
nor U3008 (N_3008,N_2739,N_2973);
xnor U3009 (N_3009,N_2912,N_2807);
nor U3010 (N_3010,N_2865,N_2984);
xor U3011 (N_3011,N_2759,N_2907);
and U3012 (N_3012,N_2706,N_2987);
or U3013 (N_3013,N_2813,N_2764);
nand U3014 (N_3014,N_2815,N_2774);
nand U3015 (N_3015,N_2966,N_2883);
or U3016 (N_3016,N_2734,N_2817);
xnor U3017 (N_3017,N_2742,N_2927);
nand U3018 (N_3018,N_2701,N_2916);
xor U3019 (N_3019,N_2920,N_2801);
or U3020 (N_3020,N_2751,N_2995);
nor U3021 (N_3021,N_2834,N_2863);
nand U3022 (N_3022,N_2988,N_2762);
or U3023 (N_3023,N_2881,N_2993);
nand U3024 (N_3024,N_2944,N_2765);
or U3025 (N_3025,N_2778,N_2905);
nor U3026 (N_3026,N_2738,N_2796);
or U3027 (N_3027,N_2975,N_2775);
xnor U3028 (N_3028,N_2960,N_2870);
and U3029 (N_3029,N_2757,N_2906);
xor U3030 (N_3030,N_2962,N_2798);
xnor U3031 (N_3031,N_2885,N_2858);
and U3032 (N_3032,N_2886,N_2924);
xor U3033 (N_3033,N_2797,N_2882);
or U3034 (N_3034,N_2898,N_2768);
nand U3035 (N_3035,N_2824,N_2873);
nor U3036 (N_3036,N_2721,N_2951);
nand U3037 (N_3037,N_2785,N_2821);
and U3038 (N_3038,N_2800,N_2715);
and U3039 (N_3039,N_2736,N_2752);
or U3040 (N_3040,N_2753,N_2979);
and U3041 (N_3041,N_2702,N_2746);
nor U3042 (N_3042,N_2866,N_2896);
and U3043 (N_3043,N_2936,N_2878);
and U3044 (N_3044,N_2719,N_2783);
nand U3045 (N_3045,N_2799,N_2848);
nor U3046 (N_3046,N_2851,N_2754);
nand U3047 (N_3047,N_2816,N_2860);
xnor U3048 (N_3048,N_2720,N_2855);
xor U3049 (N_3049,N_2758,N_2940);
nand U3050 (N_3050,N_2814,N_2879);
and U3051 (N_3051,N_2989,N_2808);
nor U3052 (N_3052,N_2921,N_2709);
nand U3053 (N_3053,N_2887,N_2953);
xnor U3054 (N_3054,N_2845,N_2733);
nand U3055 (N_3055,N_2892,N_2868);
and U3056 (N_3056,N_2784,N_2938);
and U3057 (N_3057,N_2859,N_2847);
nand U3058 (N_3058,N_2704,N_2849);
or U3059 (N_3059,N_2780,N_2820);
nor U3060 (N_3060,N_2723,N_2915);
and U3061 (N_3061,N_2901,N_2974);
nor U3062 (N_3062,N_2963,N_2895);
nand U3063 (N_3063,N_2978,N_2894);
nand U3064 (N_3064,N_2729,N_2846);
nand U3065 (N_3065,N_2823,N_2934);
or U3066 (N_3066,N_2876,N_2790);
nand U3067 (N_3067,N_2923,N_2795);
xor U3068 (N_3068,N_2958,N_2707);
or U3069 (N_3069,N_2850,N_2972);
nor U3070 (N_3070,N_2714,N_2841);
nand U3071 (N_3071,N_2840,N_2932);
nand U3072 (N_3072,N_2812,N_2893);
and U3073 (N_3073,N_2871,N_2703);
and U3074 (N_3074,N_2925,N_2727);
xor U3075 (N_3075,N_2772,N_2833);
and U3076 (N_3076,N_2747,N_2804);
nand U3077 (N_3077,N_2740,N_2745);
nand U3078 (N_3078,N_2853,N_2880);
and U3079 (N_3079,N_2929,N_2968);
and U3080 (N_3080,N_2748,N_2999);
nor U3081 (N_3081,N_2969,N_2716);
nor U3082 (N_3082,N_2954,N_2710);
nor U3083 (N_3083,N_2787,N_2922);
nand U3084 (N_3084,N_2825,N_2782);
nor U3085 (N_3085,N_2718,N_2769);
or U3086 (N_3086,N_2844,N_2843);
nand U3087 (N_3087,N_2829,N_2826);
and U3088 (N_3088,N_2914,N_2750);
nand U3089 (N_3089,N_2835,N_2862);
nand U3090 (N_3090,N_2830,N_2947);
xor U3091 (N_3091,N_2836,N_2867);
or U3092 (N_3092,N_2991,N_2964);
xor U3093 (N_3093,N_2943,N_2897);
and U3094 (N_3094,N_2950,N_2819);
xnor U3095 (N_3095,N_2937,N_2856);
or U3096 (N_3096,N_2861,N_2766);
nor U3097 (N_3097,N_2971,N_2955);
or U3098 (N_3098,N_2977,N_2842);
or U3099 (N_3099,N_2970,N_2919);
and U3100 (N_3100,N_2902,N_2941);
nand U3101 (N_3101,N_2827,N_2994);
and U3102 (N_3102,N_2949,N_2722);
and U3103 (N_3103,N_2743,N_2985);
nor U3104 (N_3104,N_2724,N_2874);
xor U3105 (N_3105,N_2942,N_2763);
nor U3106 (N_3106,N_2712,N_2777);
and U3107 (N_3107,N_2805,N_2982);
and U3108 (N_3108,N_2705,N_2904);
nand U3109 (N_3109,N_2749,N_2875);
nand U3110 (N_3110,N_2864,N_2735);
and U3111 (N_3111,N_2990,N_2838);
nand U3112 (N_3112,N_2967,N_2983);
nand U3113 (N_3113,N_2852,N_2708);
nand U3114 (N_3114,N_2900,N_2806);
and U3115 (N_3115,N_2792,N_2773);
xnor U3116 (N_3116,N_2802,N_2890);
nand U3117 (N_3117,N_2803,N_2903);
or U3118 (N_3118,N_2788,N_2789);
xor U3119 (N_3119,N_2909,N_2831);
nand U3120 (N_3120,N_2961,N_2828);
nor U3121 (N_3121,N_2711,N_2761);
nor U3122 (N_3122,N_2776,N_2965);
xnor U3123 (N_3123,N_2986,N_2930);
nor U3124 (N_3124,N_2811,N_2957);
nor U3125 (N_3125,N_2891,N_2884);
xnor U3126 (N_3126,N_2700,N_2837);
nand U3127 (N_3127,N_2781,N_2832);
and U3128 (N_3128,N_2786,N_2717);
nor U3129 (N_3129,N_2872,N_2959);
or U3130 (N_3130,N_2767,N_2756);
or U3131 (N_3131,N_2899,N_2913);
xor U3132 (N_3132,N_2869,N_2809);
nor U3133 (N_3133,N_2732,N_2933);
xor U3134 (N_3134,N_2952,N_2760);
nand U3135 (N_3135,N_2737,N_2956);
or U3136 (N_3136,N_2779,N_2996);
and U3137 (N_3137,N_2713,N_2911);
and U3138 (N_3138,N_2771,N_2928);
xnor U3139 (N_3139,N_2839,N_2998);
nand U3140 (N_3140,N_2791,N_2810);
or U3141 (N_3141,N_2981,N_2976);
nand U3142 (N_3142,N_2877,N_2926);
nor U3143 (N_3143,N_2854,N_2755);
nand U3144 (N_3144,N_2997,N_2818);
and U3145 (N_3145,N_2980,N_2888);
nor U3146 (N_3146,N_2992,N_2948);
xor U3147 (N_3147,N_2741,N_2744);
and U3148 (N_3148,N_2917,N_2770);
nor U3149 (N_3149,N_2793,N_2889);
nor U3150 (N_3150,N_2996,N_2803);
and U3151 (N_3151,N_2846,N_2785);
and U3152 (N_3152,N_2875,N_2812);
xnor U3153 (N_3153,N_2723,N_2913);
xor U3154 (N_3154,N_2912,N_2789);
or U3155 (N_3155,N_2867,N_2918);
nand U3156 (N_3156,N_2815,N_2718);
or U3157 (N_3157,N_2712,N_2980);
xnor U3158 (N_3158,N_2849,N_2904);
nand U3159 (N_3159,N_2897,N_2809);
nand U3160 (N_3160,N_2893,N_2747);
or U3161 (N_3161,N_2700,N_2803);
nand U3162 (N_3162,N_2955,N_2784);
and U3163 (N_3163,N_2711,N_2942);
nand U3164 (N_3164,N_2828,N_2858);
xnor U3165 (N_3165,N_2993,N_2754);
xor U3166 (N_3166,N_2802,N_2746);
and U3167 (N_3167,N_2976,N_2796);
and U3168 (N_3168,N_2769,N_2852);
nand U3169 (N_3169,N_2794,N_2837);
and U3170 (N_3170,N_2791,N_2955);
and U3171 (N_3171,N_2989,N_2713);
and U3172 (N_3172,N_2992,N_2791);
or U3173 (N_3173,N_2736,N_2838);
nor U3174 (N_3174,N_2704,N_2770);
and U3175 (N_3175,N_2782,N_2901);
xnor U3176 (N_3176,N_2920,N_2766);
and U3177 (N_3177,N_2721,N_2849);
nor U3178 (N_3178,N_2753,N_2950);
or U3179 (N_3179,N_2856,N_2891);
xnor U3180 (N_3180,N_2901,N_2983);
and U3181 (N_3181,N_2806,N_2787);
or U3182 (N_3182,N_2852,N_2710);
nor U3183 (N_3183,N_2783,N_2945);
nor U3184 (N_3184,N_2989,N_2937);
nand U3185 (N_3185,N_2811,N_2854);
nor U3186 (N_3186,N_2717,N_2909);
or U3187 (N_3187,N_2997,N_2728);
nand U3188 (N_3188,N_2769,N_2727);
nor U3189 (N_3189,N_2898,N_2849);
xnor U3190 (N_3190,N_2871,N_2755);
nand U3191 (N_3191,N_2812,N_2852);
and U3192 (N_3192,N_2849,N_2949);
or U3193 (N_3193,N_2793,N_2925);
or U3194 (N_3194,N_2855,N_2986);
xor U3195 (N_3195,N_2723,N_2921);
or U3196 (N_3196,N_2890,N_2859);
or U3197 (N_3197,N_2900,N_2973);
xnor U3198 (N_3198,N_2886,N_2844);
xnor U3199 (N_3199,N_2752,N_2961);
nand U3200 (N_3200,N_2952,N_2818);
nor U3201 (N_3201,N_2973,N_2956);
and U3202 (N_3202,N_2857,N_2896);
or U3203 (N_3203,N_2953,N_2994);
nor U3204 (N_3204,N_2885,N_2788);
xor U3205 (N_3205,N_2904,N_2906);
xnor U3206 (N_3206,N_2990,N_2761);
or U3207 (N_3207,N_2808,N_2864);
and U3208 (N_3208,N_2862,N_2828);
xnor U3209 (N_3209,N_2802,N_2866);
or U3210 (N_3210,N_2864,N_2746);
or U3211 (N_3211,N_2793,N_2756);
and U3212 (N_3212,N_2976,N_2986);
or U3213 (N_3213,N_2995,N_2902);
xnor U3214 (N_3214,N_2738,N_2726);
xnor U3215 (N_3215,N_2943,N_2728);
xnor U3216 (N_3216,N_2828,N_2802);
xor U3217 (N_3217,N_2836,N_2986);
nand U3218 (N_3218,N_2753,N_2945);
xnor U3219 (N_3219,N_2730,N_2965);
nand U3220 (N_3220,N_2944,N_2797);
and U3221 (N_3221,N_2747,N_2751);
nand U3222 (N_3222,N_2716,N_2792);
and U3223 (N_3223,N_2843,N_2998);
xor U3224 (N_3224,N_2802,N_2818);
and U3225 (N_3225,N_2733,N_2705);
and U3226 (N_3226,N_2829,N_2747);
and U3227 (N_3227,N_2751,N_2789);
nand U3228 (N_3228,N_2882,N_2955);
nand U3229 (N_3229,N_2922,N_2896);
or U3230 (N_3230,N_2747,N_2901);
and U3231 (N_3231,N_2733,N_2707);
and U3232 (N_3232,N_2796,N_2897);
xnor U3233 (N_3233,N_2733,N_2910);
and U3234 (N_3234,N_2906,N_2977);
and U3235 (N_3235,N_2706,N_2939);
nor U3236 (N_3236,N_2853,N_2727);
nand U3237 (N_3237,N_2847,N_2737);
and U3238 (N_3238,N_2849,N_2836);
nor U3239 (N_3239,N_2935,N_2988);
or U3240 (N_3240,N_2914,N_2969);
nand U3241 (N_3241,N_2965,N_2783);
xor U3242 (N_3242,N_2909,N_2998);
or U3243 (N_3243,N_2765,N_2707);
nand U3244 (N_3244,N_2783,N_2910);
nor U3245 (N_3245,N_2929,N_2949);
nand U3246 (N_3246,N_2880,N_2723);
nor U3247 (N_3247,N_2929,N_2955);
nor U3248 (N_3248,N_2704,N_2881);
and U3249 (N_3249,N_2929,N_2744);
nand U3250 (N_3250,N_2941,N_2936);
and U3251 (N_3251,N_2765,N_2961);
nand U3252 (N_3252,N_2747,N_2874);
or U3253 (N_3253,N_2771,N_2992);
or U3254 (N_3254,N_2947,N_2760);
nor U3255 (N_3255,N_2931,N_2974);
nor U3256 (N_3256,N_2967,N_2883);
xnor U3257 (N_3257,N_2936,N_2965);
nand U3258 (N_3258,N_2740,N_2903);
or U3259 (N_3259,N_2923,N_2866);
nor U3260 (N_3260,N_2818,N_2981);
or U3261 (N_3261,N_2752,N_2895);
nand U3262 (N_3262,N_2843,N_2848);
xnor U3263 (N_3263,N_2843,N_2737);
xor U3264 (N_3264,N_2884,N_2773);
or U3265 (N_3265,N_2707,N_2750);
and U3266 (N_3266,N_2868,N_2829);
or U3267 (N_3267,N_2875,N_2804);
nand U3268 (N_3268,N_2904,N_2728);
or U3269 (N_3269,N_2792,N_2872);
or U3270 (N_3270,N_2998,N_2974);
xnor U3271 (N_3271,N_2706,N_2986);
nor U3272 (N_3272,N_2911,N_2845);
or U3273 (N_3273,N_2701,N_2954);
nand U3274 (N_3274,N_2874,N_2706);
xor U3275 (N_3275,N_2826,N_2742);
or U3276 (N_3276,N_2842,N_2791);
or U3277 (N_3277,N_2875,N_2853);
nor U3278 (N_3278,N_2756,N_2700);
nand U3279 (N_3279,N_2707,N_2825);
and U3280 (N_3280,N_2964,N_2990);
or U3281 (N_3281,N_2816,N_2843);
and U3282 (N_3282,N_2881,N_2710);
nand U3283 (N_3283,N_2997,N_2972);
nand U3284 (N_3284,N_2918,N_2806);
nand U3285 (N_3285,N_2975,N_2922);
nor U3286 (N_3286,N_2804,N_2750);
nand U3287 (N_3287,N_2797,N_2825);
or U3288 (N_3288,N_2768,N_2717);
xnor U3289 (N_3289,N_2984,N_2897);
nor U3290 (N_3290,N_2792,N_2946);
and U3291 (N_3291,N_2825,N_2921);
xnor U3292 (N_3292,N_2832,N_2950);
and U3293 (N_3293,N_2851,N_2849);
xnor U3294 (N_3294,N_2899,N_2723);
or U3295 (N_3295,N_2719,N_2932);
nor U3296 (N_3296,N_2824,N_2862);
and U3297 (N_3297,N_2738,N_2805);
or U3298 (N_3298,N_2816,N_2819);
or U3299 (N_3299,N_2792,N_2715);
xor U3300 (N_3300,N_3257,N_3186);
nand U3301 (N_3301,N_3219,N_3125);
or U3302 (N_3302,N_3123,N_3046);
and U3303 (N_3303,N_3194,N_3025);
nand U3304 (N_3304,N_3007,N_3093);
xor U3305 (N_3305,N_3299,N_3058);
nor U3306 (N_3306,N_3107,N_3191);
xor U3307 (N_3307,N_3079,N_3032);
and U3308 (N_3308,N_3259,N_3020);
and U3309 (N_3309,N_3118,N_3236);
nor U3310 (N_3310,N_3222,N_3129);
nor U3311 (N_3311,N_3171,N_3014);
nand U3312 (N_3312,N_3266,N_3000);
nand U3313 (N_3313,N_3183,N_3089);
nand U3314 (N_3314,N_3182,N_3128);
nand U3315 (N_3315,N_3006,N_3174);
xor U3316 (N_3316,N_3167,N_3111);
xor U3317 (N_3317,N_3164,N_3292);
and U3318 (N_3318,N_3240,N_3022);
xor U3319 (N_3319,N_3094,N_3038);
xor U3320 (N_3320,N_3287,N_3012);
nand U3321 (N_3321,N_3075,N_3083);
nand U3322 (N_3322,N_3049,N_3248);
xor U3323 (N_3323,N_3192,N_3126);
or U3324 (N_3324,N_3003,N_3071);
and U3325 (N_3325,N_3291,N_3069);
and U3326 (N_3326,N_3055,N_3279);
and U3327 (N_3327,N_3253,N_3241);
xor U3328 (N_3328,N_3065,N_3036);
and U3329 (N_3329,N_3176,N_3010);
and U3330 (N_3330,N_3105,N_3269);
nor U3331 (N_3331,N_3024,N_3161);
and U3332 (N_3332,N_3189,N_3132);
nor U3333 (N_3333,N_3195,N_3286);
nand U3334 (N_3334,N_3138,N_3281);
nand U3335 (N_3335,N_3102,N_3116);
xor U3336 (N_3336,N_3270,N_3016);
or U3337 (N_3337,N_3205,N_3296);
nor U3338 (N_3338,N_3092,N_3288);
nor U3339 (N_3339,N_3005,N_3115);
or U3340 (N_3340,N_3229,N_3095);
nand U3341 (N_3341,N_3216,N_3066);
nor U3342 (N_3342,N_3117,N_3148);
xor U3343 (N_3343,N_3088,N_3063);
nor U3344 (N_3344,N_3218,N_3048);
xnor U3345 (N_3345,N_3208,N_3168);
nand U3346 (N_3346,N_3052,N_3059);
and U3347 (N_3347,N_3018,N_3134);
nand U3348 (N_3348,N_3173,N_3207);
and U3349 (N_3349,N_3251,N_3060);
or U3350 (N_3350,N_3143,N_3154);
nor U3351 (N_3351,N_3243,N_3033);
or U3352 (N_3352,N_3106,N_3230);
and U3353 (N_3353,N_3015,N_3085);
nor U3354 (N_3354,N_3001,N_3011);
nor U3355 (N_3355,N_3247,N_3004);
xor U3356 (N_3356,N_3170,N_3009);
or U3357 (N_3357,N_3023,N_3228);
and U3358 (N_3358,N_3097,N_3239);
or U3359 (N_3359,N_3262,N_3149);
xnor U3360 (N_3360,N_3080,N_3057);
nor U3361 (N_3361,N_3177,N_3213);
or U3362 (N_3362,N_3180,N_3068);
nor U3363 (N_3363,N_3050,N_3285);
or U3364 (N_3364,N_3127,N_3271);
nor U3365 (N_3365,N_3275,N_3045);
nand U3366 (N_3366,N_3153,N_3114);
and U3367 (N_3367,N_3233,N_3197);
nor U3368 (N_3368,N_3013,N_3273);
xor U3369 (N_3369,N_3072,N_3133);
xnor U3370 (N_3370,N_3254,N_3037);
or U3371 (N_3371,N_3157,N_3086);
or U3372 (N_3372,N_3031,N_3096);
nor U3373 (N_3373,N_3297,N_3258);
xor U3374 (N_3374,N_3109,N_3263);
or U3375 (N_3375,N_3108,N_3293);
nor U3376 (N_3376,N_3277,N_3224);
or U3377 (N_3377,N_3200,N_3294);
or U3378 (N_3378,N_3227,N_3193);
nor U3379 (N_3379,N_3112,N_3122);
nand U3380 (N_3380,N_3077,N_3017);
or U3381 (N_3381,N_3039,N_3130);
or U3382 (N_3382,N_3231,N_3078);
and U3383 (N_3383,N_3163,N_3204);
nor U3384 (N_3384,N_3196,N_3256);
or U3385 (N_3385,N_3245,N_3198);
xnor U3386 (N_3386,N_3220,N_3145);
or U3387 (N_3387,N_3042,N_3178);
xnor U3388 (N_3388,N_3061,N_3278);
nor U3389 (N_3389,N_3242,N_3087);
nor U3390 (N_3390,N_3158,N_3113);
nor U3391 (N_3391,N_3099,N_3289);
and U3392 (N_3392,N_3298,N_3203);
or U3393 (N_3393,N_3152,N_3265);
or U3394 (N_3394,N_3151,N_3104);
nand U3395 (N_3395,N_3201,N_3119);
nor U3396 (N_3396,N_3062,N_3249);
or U3397 (N_3397,N_3139,N_3255);
xnor U3398 (N_3398,N_3141,N_3043);
xnor U3399 (N_3399,N_3237,N_3206);
or U3400 (N_3400,N_3274,N_3029);
nor U3401 (N_3401,N_3047,N_3181);
xor U3402 (N_3402,N_3226,N_3051);
and U3403 (N_3403,N_3234,N_3188);
or U3404 (N_3404,N_3008,N_3054);
nand U3405 (N_3405,N_3140,N_3187);
and U3406 (N_3406,N_3210,N_3290);
and U3407 (N_3407,N_3067,N_3244);
nand U3408 (N_3408,N_3041,N_3150);
xor U3409 (N_3409,N_3053,N_3144);
or U3410 (N_3410,N_3267,N_3160);
nor U3411 (N_3411,N_3021,N_3030);
and U3412 (N_3412,N_3135,N_3044);
and U3413 (N_3413,N_3040,N_3162);
nor U3414 (N_3414,N_3002,N_3147);
xnor U3415 (N_3415,N_3137,N_3120);
and U3416 (N_3416,N_3246,N_3084);
and U3417 (N_3417,N_3110,N_3272);
xnor U3418 (N_3418,N_3172,N_3217);
or U3419 (N_3419,N_3250,N_3225);
xor U3420 (N_3420,N_3019,N_3261);
xnor U3421 (N_3421,N_3070,N_3284);
xnor U3422 (N_3422,N_3185,N_3121);
nor U3423 (N_3423,N_3260,N_3103);
or U3424 (N_3424,N_3136,N_3081);
nor U3425 (N_3425,N_3076,N_3142);
nor U3426 (N_3426,N_3166,N_3175);
and U3427 (N_3427,N_3026,N_3276);
and U3428 (N_3428,N_3264,N_3156);
nand U3429 (N_3429,N_3074,N_3202);
nor U3430 (N_3430,N_3235,N_3221);
xnor U3431 (N_3431,N_3280,N_3082);
nor U3432 (N_3432,N_3282,N_3064);
xnor U3433 (N_3433,N_3295,N_3268);
nand U3434 (N_3434,N_3027,N_3056);
or U3435 (N_3435,N_3124,N_3184);
nand U3436 (N_3436,N_3028,N_3101);
nor U3437 (N_3437,N_3131,N_3232);
and U3438 (N_3438,N_3214,N_3165);
nor U3439 (N_3439,N_3159,N_3283);
xnor U3440 (N_3440,N_3212,N_3169);
nand U3441 (N_3441,N_3146,N_3034);
nor U3442 (N_3442,N_3090,N_3211);
nand U3443 (N_3443,N_3091,N_3035);
or U3444 (N_3444,N_3100,N_3252);
nor U3445 (N_3445,N_3238,N_3155);
xor U3446 (N_3446,N_3199,N_3190);
nand U3447 (N_3447,N_3073,N_3179);
nand U3448 (N_3448,N_3215,N_3098);
or U3449 (N_3449,N_3209,N_3223);
and U3450 (N_3450,N_3125,N_3008);
nor U3451 (N_3451,N_3070,N_3001);
and U3452 (N_3452,N_3006,N_3098);
or U3453 (N_3453,N_3101,N_3255);
xor U3454 (N_3454,N_3291,N_3043);
xor U3455 (N_3455,N_3267,N_3253);
nand U3456 (N_3456,N_3213,N_3264);
and U3457 (N_3457,N_3241,N_3171);
xor U3458 (N_3458,N_3133,N_3010);
nand U3459 (N_3459,N_3014,N_3076);
nor U3460 (N_3460,N_3218,N_3101);
and U3461 (N_3461,N_3196,N_3109);
and U3462 (N_3462,N_3175,N_3246);
or U3463 (N_3463,N_3269,N_3286);
or U3464 (N_3464,N_3186,N_3264);
xor U3465 (N_3465,N_3042,N_3168);
or U3466 (N_3466,N_3075,N_3157);
and U3467 (N_3467,N_3210,N_3154);
nor U3468 (N_3468,N_3096,N_3297);
nor U3469 (N_3469,N_3100,N_3274);
and U3470 (N_3470,N_3207,N_3273);
nor U3471 (N_3471,N_3163,N_3243);
or U3472 (N_3472,N_3208,N_3289);
nor U3473 (N_3473,N_3223,N_3011);
nor U3474 (N_3474,N_3072,N_3065);
xor U3475 (N_3475,N_3060,N_3247);
nand U3476 (N_3476,N_3097,N_3096);
xnor U3477 (N_3477,N_3166,N_3298);
xor U3478 (N_3478,N_3152,N_3277);
nor U3479 (N_3479,N_3179,N_3268);
and U3480 (N_3480,N_3294,N_3224);
nand U3481 (N_3481,N_3257,N_3031);
nor U3482 (N_3482,N_3233,N_3024);
or U3483 (N_3483,N_3159,N_3130);
xor U3484 (N_3484,N_3160,N_3263);
xor U3485 (N_3485,N_3162,N_3240);
nor U3486 (N_3486,N_3051,N_3181);
nand U3487 (N_3487,N_3204,N_3108);
xor U3488 (N_3488,N_3000,N_3109);
nand U3489 (N_3489,N_3236,N_3096);
nand U3490 (N_3490,N_3106,N_3164);
or U3491 (N_3491,N_3010,N_3246);
nor U3492 (N_3492,N_3124,N_3032);
nor U3493 (N_3493,N_3152,N_3058);
nor U3494 (N_3494,N_3156,N_3263);
nor U3495 (N_3495,N_3040,N_3213);
nand U3496 (N_3496,N_3221,N_3216);
nand U3497 (N_3497,N_3119,N_3150);
xnor U3498 (N_3498,N_3217,N_3056);
nand U3499 (N_3499,N_3010,N_3271);
xnor U3500 (N_3500,N_3265,N_3278);
nor U3501 (N_3501,N_3017,N_3097);
nand U3502 (N_3502,N_3290,N_3198);
or U3503 (N_3503,N_3081,N_3159);
xor U3504 (N_3504,N_3241,N_3125);
xnor U3505 (N_3505,N_3252,N_3064);
xor U3506 (N_3506,N_3058,N_3075);
and U3507 (N_3507,N_3018,N_3053);
and U3508 (N_3508,N_3089,N_3026);
and U3509 (N_3509,N_3169,N_3204);
nor U3510 (N_3510,N_3138,N_3007);
nor U3511 (N_3511,N_3108,N_3259);
or U3512 (N_3512,N_3123,N_3110);
or U3513 (N_3513,N_3148,N_3295);
xor U3514 (N_3514,N_3105,N_3138);
nor U3515 (N_3515,N_3154,N_3193);
nand U3516 (N_3516,N_3092,N_3281);
xnor U3517 (N_3517,N_3056,N_3166);
nor U3518 (N_3518,N_3207,N_3005);
nand U3519 (N_3519,N_3254,N_3240);
or U3520 (N_3520,N_3103,N_3017);
nor U3521 (N_3521,N_3013,N_3147);
nor U3522 (N_3522,N_3099,N_3083);
or U3523 (N_3523,N_3001,N_3187);
xor U3524 (N_3524,N_3173,N_3234);
and U3525 (N_3525,N_3063,N_3276);
and U3526 (N_3526,N_3103,N_3165);
xor U3527 (N_3527,N_3166,N_3253);
and U3528 (N_3528,N_3178,N_3128);
xor U3529 (N_3529,N_3131,N_3262);
xnor U3530 (N_3530,N_3195,N_3219);
nand U3531 (N_3531,N_3224,N_3080);
or U3532 (N_3532,N_3153,N_3159);
nand U3533 (N_3533,N_3169,N_3065);
xnor U3534 (N_3534,N_3069,N_3063);
and U3535 (N_3535,N_3213,N_3101);
nand U3536 (N_3536,N_3098,N_3063);
nor U3537 (N_3537,N_3149,N_3025);
or U3538 (N_3538,N_3193,N_3290);
and U3539 (N_3539,N_3143,N_3277);
xnor U3540 (N_3540,N_3044,N_3002);
xnor U3541 (N_3541,N_3137,N_3101);
or U3542 (N_3542,N_3252,N_3098);
xnor U3543 (N_3543,N_3241,N_3126);
and U3544 (N_3544,N_3185,N_3110);
xnor U3545 (N_3545,N_3018,N_3157);
nand U3546 (N_3546,N_3037,N_3015);
xnor U3547 (N_3547,N_3021,N_3088);
nor U3548 (N_3548,N_3266,N_3015);
or U3549 (N_3549,N_3222,N_3297);
or U3550 (N_3550,N_3001,N_3006);
nand U3551 (N_3551,N_3263,N_3124);
nor U3552 (N_3552,N_3251,N_3165);
or U3553 (N_3553,N_3049,N_3222);
or U3554 (N_3554,N_3242,N_3166);
and U3555 (N_3555,N_3196,N_3122);
nand U3556 (N_3556,N_3028,N_3193);
or U3557 (N_3557,N_3030,N_3137);
or U3558 (N_3558,N_3212,N_3139);
xor U3559 (N_3559,N_3223,N_3137);
nand U3560 (N_3560,N_3240,N_3186);
xor U3561 (N_3561,N_3274,N_3193);
nor U3562 (N_3562,N_3177,N_3011);
or U3563 (N_3563,N_3185,N_3222);
nand U3564 (N_3564,N_3094,N_3078);
or U3565 (N_3565,N_3064,N_3246);
or U3566 (N_3566,N_3136,N_3182);
nor U3567 (N_3567,N_3018,N_3209);
nand U3568 (N_3568,N_3221,N_3167);
nor U3569 (N_3569,N_3194,N_3096);
and U3570 (N_3570,N_3170,N_3186);
xor U3571 (N_3571,N_3145,N_3080);
nor U3572 (N_3572,N_3075,N_3081);
or U3573 (N_3573,N_3153,N_3270);
and U3574 (N_3574,N_3248,N_3089);
nand U3575 (N_3575,N_3268,N_3132);
nand U3576 (N_3576,N_3078,N_3023);
nor U3577 (N_3577,N_3011,N_3034);
or U3578 (N_3578,N_3234,N_3042);
xnor U3579 (N_3579,N_3226,N_3281);
and U3580 (N_3580,N_3286,N_3016);
xnor U3581 (N_3581,N_3192,N_3229);
nand U3582 (N_3582,N_3003,N_3045);
nand U3583 (N_3583,N_3001,N_3125);
nor U3584 (N_3584,N_3112,N_3225);
nor U3585 (N_3585,N_3021,N_3090);
nor U3586 (N_3586,N_3072,N_3171);
xor U3587 (N_3587,N_3240,N_3229);
nand U3588 (N_3588,N_3028,N_3033);
and U3589 (N_3589,N_3115,N_3210);
or U3590 (N_3590,N_3291,N_3156);
nor U3591 (N_3591,N_3168,N_3181);
xor U3592 (N_3592,N_3251,N_3209);
or U3593 (N_3593,N_3065,N_3197);
nor U3594 (N_3594,N_3070,N_3171);
xor U3595 (N_3595,N_3226,N_3160);
xor U3596 (N_3596,N_3039,N_3188);
xnor U3597 (N_3597,N_3090,N_3180);
nand U3598 (N_3598,N_3205,N_3125);
nor U3599 (N_3599,N_3259,N_3072);
and U3600 (N_3600,N_3352,N_3327);
xnor U3601 (N_3601,N_3535,N_3350);
nor U3602 (N_3602,N_3317,N_3523);
or U3603 (N_3603,N_3530,N_3356);
xnor U3604 (N_3604,N_3384,N_3357);
or U3605 (N_3605,N_3441,N_3528);
nor U3606 (N_3606,N_3454,N_3568);
and U3607 (N_3607,N_3456,N_3566);
nand U3608 (N_3608,N_3449,N_3473);
or U3609 (N_3609,N_3544,N_3585);
or U3610 (N_3610,N_3436,N_3391);
nand U3611 (N_3611,N_3533,N_3539);
xnor U3612 (N_3612,N_3598,N_3513);
or U3613 (N_3613,N_3440,N_3435);
xnor U3614 (N_3614,N_3331,N_3442);
and U3615 (N_3615,N_3363,N_3467);
xnor U3616 (N_3616,N_3344,N_3531);
nor U3617 (N_3617,N_3348,N_3494);
nor U3618 (N_3618,N_3332,N_3583);
xnor U3619 (N_3619,N_3592,N_3377);
and U3620 (N_3620,N_3394,N_3323);
and U3621 (N_3621,N_3554,N_3489);
and U3622 (N_3622,N_3591,N_3371);
xor U3623 (N_3623,N_3461,N_3507);
nor U3624 (N_3624,N_3315,N_3556);
and U3625 (N_3625,N_3477,N_3532);
nand U3626 (N_3626,N_3309,N_3369);
nor U3627 (N_3627,N_3515,N_3355);
xor U3628 (N_3628,N_3445,N_3307);
or U3629 (N_3629,N_3413,N_3486);
and U3630 (N_3630,N_3433,N_3476);
nor U3631 (N_3631,N_3590,N_3395);
or U3632 (N_3632,N_3412,N_3541);
or U3633 (N_3633,N_3574,N_3506);
xor U3634 (N_3634,N_3399,N_3409);
nand U3635 (N_3635,N_3316,N_3347);
xnor U3636 (N_3636,N_3415,N_3500);
or U3637 (N_3637,N_3346,N_3563);
xnor U3638 (N_3638,N_3479,N_3520);
or U3639 (N_3639,N_3376,N_3587);
and U3640 (N_3640,N_3326,N_3542);
nor U3641 (N_3641,N_3322,N_3349);
nand U3642 (N_3642,N_3337,N_3559);
and U3643 (N_3643,N_3504,N_3519);
nand U3644 (N_3644,N_3543,N_3334);
nand U3645 (N_3645,N_3594,N_3397);
nand U3646 (N_3646,N_3368,N_3407);
nand U3647 (N_3647,N_3548,N_3458);
xor U3648 (N_3648,N_3573,N_3300);
and U3649 (N_3649,N_3429,N_3596);
xor U3650 (N_3650,N_3552,N_3342);
nand U3651 (N_3651,N_3540,N_3324);
and U3652 (N_3652,N_3450,N_3453);
or U3653 (N_3653,N_3372,N_3405);
and U3654 (N_3654,N_3571,N_3444);
nand U3655 (N_3655,N_3595,N_3546);
nor U3656 (N_3656,N_3373,N_3398);
nor U3657 (N_3657,N_3484,N_3538);
and U3658 (N_3658,N_3490,N_3560);
nor U3659 (N_3659,N_3330,N_3410);
or U3660 (N_3660,N_3553,N_3313);
xor U3661 (N_3661,N_3432,N_3304);
and U3662 (N_3662,N_3478,N_3509);
and U3663 (N_3663,N_3597,N_3392);
or U3664 (N_3664,N_3408,N_3565);
nor U3665 (N_3665,N_3516,N_3488);
and U3666 (N_3666,N_3406,N_3366);
xnor U3667 (N_3667,N_3501,N_3470);
nand U3668 (N_3668,N_3321,N_3562);
xnor U3669 (N_3669,N_3320,N_3498);
and U3670 (N_3670,N_3381,N_3517);
or U3671 (N_3671,N_3529,N_3588);
or U3672 (N_3672,N_3380,N_3522);
and U3673 (N_3673,N_3362,N_3459);
and U3674 (N_3674,N_3303,N_3464);
and U3675 (N_3675,N_3434,N_3510);
xor U3676 (N_3676,N_3319,N_3534);
nand U3677 (N_3677,N_3420,N_3555);
and U3678 (N_3678,N_3382,N_3425);
nand U3679 (N_3679,N_3580,N_3495);
xnor U3680 (N_3680,N_3482,N_3452);
or U3681 (N_3681,N_3389,N_3448);
and U3682 (N_3682,N_3387,N_3401);
xnor U3683 (N_3683,N_3483,N_3577);
xor U3684 (N_3684,N_3561,N_3423);
nor U3685 (N_3685,N_3526,N_3466);
xor U3686 (N_3686,N_3314,N_3469);
nand U3687 (N_3687,N_3505,N_3305);
and U3688 (N_3688,N_3474,N_3338);
nor U3689 (N_3689,N_3365,N_3567);
nand U3690 (N_3690,N_3599,N_3312);
or U3691 (N_3691,N_3447,N_3537);
xnor U3692 (N_3692,N_3462,N_3460);
nor U3693 (N_3693,N_3385,N_3302);
nand U3694 (N_3694,N_3421,N_3499);
xor U3695 (N_3695,N_3438,N_3388);
xnor U3696 (N_3696,N_3351,N_3339);
nor U3697 (N_3697,N_3343,N_3579);
and U3698 (N_3698,N_3481,N_3325);
and U3699 (N_3699,N_3443,N_3581);
xor U3700 (N_3700,N_3364,N_3578);
and U3701 (N_3701,N_3508,N_3422);
or U3702 (N_3702,N_3359,N_3393);
nor U3703 (N_3703,N_3518,N_3502);
nor U3704 (N_3704,N_3416,N_3572);
xor U3705 (N_3705,N_3301,N_3426);
nor U3706 (N_3706,N_3336,N_3335);
nand U3707 (N_3707,N_3471,N_3428);
xor U3708 (N_3708,N_3536,N_3485);
xnor U3709 (N_3709,N_3463,N_3524);
and U3710 (N_3710,N_3308,N_3512);
nor U3711 (N_3711,N_3589,N_3402);
or U3712 (N_3712,N_3427,N_3419);
nand U3713 (N_3713,N_3551,N_3378);
nor U3714 (N_3714,N_3493,N_3576);
nor U3715 (N_3715,N_3558,N_3549);
nand U3716 (N_3716,N_3403,N_3468);
nor U3717 (N_3717,N_3569,N_3545);
nor U3718 (N_3718,N_3390,N_3593);
or U3719 (N_3719,N_3367,N_3496);
xnor U3720 (N_3720,N_3311,N_3418);
nor U3721 (N_3721,N_3310,N_3455);
nor U3722 (N_3722,N_3437,N_3375);
and U3723 (N_3723,N_3396,N_3480);
xor U3724 (N_3724,N_3353,N_3527);
nor U3725 (N_3725,N_3345,N_3439);
and U3726 (N_3726,N_3329,N_3370);
and U3727 (N_3727,N_3451,N_3582);
or U3728 (N_3728,N_3411,N_3503);
nand U3729 (N_3729,N_3586,N_3491);
xnor U3730 (N_3730,N_3358,N_3521);
nand U3731 (N_3731,N_3400,N_3472);
or U3732 (N_3732,N_3570,N_3446);
nand U3733 (N_3733,N_3457,N_3333);
xor U3734 (N_3734,N_3383,N_3374);
or U3735 (N_3735,N_3525,N_3475);
nand U3736 (N_3736,N_3341,N_3306);
nand U3737 (N_3737,N_3547,N_3492);
xnor U3738 (N_3738,N_3354,N_3550);
nor U3739 (N_3739,N_3414,N_3404);
xor U3740 (N_3740,N_3417,N_3318);
xnor U3741 (N_3741,N_3557,N_3497);
or U3742 (N_3742,N_3575,N_3379);
or U3743 (N_3743,N_3386,N_3511);
xor U3744 (N_3744,N_3360,N_3487);
nor U3745 (N_3745,N_3424,N_3564);
or U3746 (N_3746,N_3514,N_3340);
or U3747 (N_3747,N_3584,N_3465);
and U3748 (N_3748,N_3430,N_3431);
nor U3749 (N_3749,N_3328,N_3361);
and U3750 (N_3750,N_3455,N_3545);
nand U3751 (N_3751,N_3457,N_3590);
xor U3752 (N_3752,N_3496,N_3516);
nor U3753 (N_3753,N_3471,N_3588);
nor U3754 (N_3754,N_3428,N_3303);
or U3755 (N_3755,N_3522,N_3535);
nand U3756 (N_3756,N_3583,N_3560);
nor U3757 (N_3757,N_3456,N_3426);
nand U3758 (N_3758,N_3379,N_3572);
or U3759 (N_3759,N_3485,N_3467);
nor U3760 (N_3760,N_3312,N_3440);
and U3761 (N_3761,N_3456,N_3553);
nor U3762 (N_3762,N_3338,N_3334);
nand U3763 (N_3763,N_3548,N_3569);
or U3764 (N_3764,N_3598,N_3356);
nor U3765 (N_3765,N_3397,N_3582);
nand U3766 (N_3766,N_3569,N_3317);
nor U3767 (N_3767,N_3335,N_3490);
nand U3768 (N_3768,N_3589,N_3573);
nand U3769 (N_3769,N_3573,N_3428);
and U3770 (N_3770,N_3512,N_3420);
nor U3771 (N_3771,N_3437,N_3405);
nor U3772 (N_3772,N_3484,N_3333);
or U3773 (N_3773,N_3315,N_3572);
and U3774 (N_3774,N_3440,N_3500);
xor U3775 (N_3775,N_3333,N_3316);
nor U3776 (N_3776,N_3424,N_3427);
and U3777 (N_3777,N_3327,N_3337);
and U3778 (N_3778,N_3325,N_3598);
nand U3779 (N_3779,N_3351,N_3368);
and U3780 (N_3780,N_3522,N_3497);
nor U3781 (N_3781,N_3462,N_3533);
and U3782 (N_3782,N_3302,N_3482);
or U3783 (N_3783,N_3454,N_3412);
or U3784 (N_3784,N_3369,N_3412);
and U3785 (N_3785,N_3343,N_3336);
nor U3786 (N_3786,N_3394,N_3478);
or U3787 (N_3787,N_3411,N_3404);
nor U3788 (N_3788,N_3401,N_3573);
nor U3789 (N_3789,N_3399,N_3415);
xnor U3790 (N_3790,N_3308,N_3412);
xnor U3791 (N_3791,N_3563,N_3352);
nand U3792 (N_3792,N_3487,N_3354);
or U3793 (N_3793,N_3580,N_3525);
nand U3794 (N_3794,N_3484,N_3454);
xnor U3795 (N_3795,N_3449,N_3533);
and U3796 (N_3796,N_3491,N_3434);
and U3797 (N_3797,N_3384,N_3505);
nor U3798 (N_3798,N_3440,N_3457);
xnor U3799 (N_3799,N_3543,N_3472);
nand U3800 (N_3800,N_3415,N_3352);
and U3801 (N_3801,N_3492,N_3316);
nor U3802 (N_3802,N_3524,N_3446);
or U3803 (N_3803,N_3361,N_3543);
and U3804 (N_3804,N_3517,N_3310);
xor U3805 (N_3805,N_3441,N_3511);
nand U3806 (N_3806,N_3545,N_3343);
xor U3807 (N_3807,N_3505,N_3570);
or U3808 (N_3808,N_3499,N_3378);
xnor U3809 (N_3809,N_3503,N_3444);
xor U3810 (N_3810,N_3417,N_3399);
nand U3811 (N_3811,N_3372,N_3341);
xnor U3812 (N_3812,N_3485,N_3521);
nand U3813 (N_3813,N_3377,N_3460);
nand U3814 (N_3814,N_3342,N_3333);
nand U3815 (N_3815,N_3378,N_3300);
nand U3816 (N_3816,N_3401,N_3513);
nand U3817 (N_3817,N_3527,N_3540);
nand U3818 (N_3818,N_3360,N_3321);
nor U3819 (N_3819,N_3504,N_3345);
xnor U3820 (N_3820,N_3405,N_3423);
nor U3821 (N_3821,N_3422,N_3323);
xor U3822 (N_3822,N_3401,N_3406);
or U3823 (N_3823,N_3363,N_3447);
or U3824 (N_3824,N_3436,N_3494);
and U3825 (N_3825,N_3323,N_3402);
and U3826 (N_3826,N_3542,N_3365);
nor U3827 (N_3827,N_3401,N_3503);
and U3828 (N_3828,N_3565,N_3368);
and U3829 (N_3829,N_3531,N_3468);
nor U3830 (N_3830,N_3567,N_3495);
or U3831 (N_3831,N_3340,N_3484);
nor U3832 (N_3832,N_3511,N_3440);
and U3833 (N_3833,N_3570,N_3530);
or U3834 (N_3834,N_3355,N_3528);
or U3835 (N_3835,N_3310,N_3503);
and U3836 (N_3836,N_3393,N_3547);
or U3837 (N_3837,N_3377,N_3447);
and U3838 (N_3838,N_3344,N_3493);
nor U3839 (N_3839,N_3354,N_3443);
and U3840 (N_3840,N_3438,N_3586);
or U3841 (N_3841,N_3564,N_3371);
nor U3842 (N_3842,N_3300,N_3563);
nand U3843 (N_3843,N_3314,N_3415);
xor U3844 (N_3844,N_3576,N_3458);
and U3845 (N_3845,N_3462,N_3409);
xor U3846 (N_3846,N_3559,N_3405);
and U3847 (N_3847,N_3416,N_3386);
nand U3848 (N_3848,N_3559,N_3328);
xor U3849 (N_3849,N_3574,N_3590);
and U3850 (N_3850,N_3436,N_3380);
xnor U3851 (N_3851,N_3568,N_3541);
or U3852 (N_3852,N_3452,N_3463);
xor U3853 (N_3853,N_3310,N_3507);
or U3854 (N_3854,N_3470,N_3459);
or U3855 (N_3855,N_3575,N_3311);
xor U3856 (N_3856,N_3450,N_3424);
nor U3857 (N_3857,N_3340,N_3472);
nor U3858 (N_3858,N_3510,N_3580);
nor U3859 (N_3859,N_3454,N_3322);
nor U3860 (N_3860,N_3355,N_3300);
and U3861 (N_3861,N_3530,N_3567);
xor U3862 (N_3862,N_3541,N_3551);
xor U3863 (N_3863,N_3476,N_3369);
or U3864 (N_3864,N_3441,N_3526);
and U3865 (N_3865,N_3569,N_3559);
nand U3866 (N_3866,N_3593,N_3397);
nand U3867 (N_3867,N_3599,N_3455);
nand U3868 (N_3868,N_3348,N_3353);
nand U3869 (N_3869,N_3361,N_3502);
nand U3870 (N_3870,N_3355,N_3404);
xnor U3871 (N_3871,N_3436,N_3510);
and U3872 (N_3872,N_3588,N_3568);
or U3873 (N_3873,N_3486,N_3548);
nand U3874 (N_3874,N_3341,N_3413);
nor U3875 (N_3875,N_3524,N_3570);
or U3876 (N_3876,N_3563,N_3439);
and U3877 (N_3877,N_3574,N_3526);
nand U3878 (N_3878,N_3373,N_3306);
and U3879 (N_3879,N_3535,N_3480);
and U3880 (N_3880,N_3510,N_3338);
nand U3881 (N_3881,N_3546,N_3332);
and U3882 (N_3882,N_3390,N_3508);
xnor U3883 (N_3883,N_3389,N_3417);
and U3884 (N_3884,N_3486,N_3524);
nand U3885 (N_3885,N_3356,N_3407);
nor U3886 (N_3886,N_3359,N_3406);
and U3887 (N_3887,N_3536,N_3521);
nor U3888 (N_3888,N_3403,N_3323);
nand U3889 (N_3889,N_3308,N_3397);
nor U3890 (N_3890,N_3400,N_3508);
and U3891 (N_3891,N_3335,N_3432);
nor U3892 (N_3892,N_3364,N_3466);
nor U3893 (N_3893,N_3414,N_3402);
or U3894 (N_3894,N_3386,N_3496);
and U3895 (N_3895,N_3571,N_3531);
xor U3896 (N_3896,N_3411,N_3336);
and U3897 (N_3897,N_3300,N_3368);
nor U3898 (N_3898,N_3304,N_3552);
and U3899 (N_3899,N_3502,N_3377);
xnor U3900 (N_3900,N_3813,N_3770);
or U3901 (N_3901,N_3837,N_3631);
xnor U3902 (N_3902,N_3853,N_3835);
and U3903 (N_3903,N_3693,N_3734);
nor U3904 (N_3904,N_3721,N_3867);
nor U3905 (N_3905,N_3619,N_3610);
or U3906 (N_3906,N_3681,N_3695);
nor U3907 (N_3907,N_3869,N_3609);
nor U3908 (N_3908,N_3843,N_3830);
xor U3909 (N_3909,N_3859,N_3738);
nor U3910 (N_3910,N_3688,N_3742);
and U3911 (N_3911,N_3884,N_3653);
nand U3912 (N_3912,N_3777,N_3698);
nand U3913 (N_3913,N_3745,N_3793);
and U3914 (N_3914,N_3800,N_3799);
xor U3915 (N_3915,N_3611,N_3879);
nor U3916 (N_3916,N_3739,N_3840);
xnor U3917 (N_3917,N_3749,N_3851);
or U3918 (N_3918,N_3862,N_3806);
nand U3919 (N_3919,N_3651,N_3877);
xor U3920 (N_3920,N_3831,N_3866);
and U3921 (N_3921,N_3684,N_3661);
xor U3922 (N_3922,N_3662,N_3704);
and U3923 (N_3923,N_3630,N_3640);
nor U3924 (N_3924,N_3743,N_3798);
or U3925 (N_3925,N_3679,N_3622);
nor U3926 (N_3926,N_3687,N_3827);
nor U3927 (N_3927,N_3892,N_3784);
xnor U3928 (N_3928,N_3621,N_3678);
xor U3929 (N_3929,N_3825,N_3861);
xor U3930 (N_3930,N_3846,N_3744);
and U3931 (N_3931,N_3849,N_3834);
nand U3932 (N_3932,N_3774,N_3768);
xnor U3933 (N_3933,N_3636,N_3603);
or U3934 (N_3934,N_3863,N_3880);
xnor U3935 (N_3935,N_3865,N_3864);
nand U3936 (N_3936,N_3785,N_3733);
nor U3937 (N_3937,N_3690,N_3729);
or U3938 (N_3938,N_3815,N_3606);
nor U3939 (N_3939,N_3665,N_3796);
or U3940 (N_3940,N_3847,N_3720);
nand U3941 (N_3941,N_3642,N_3699);
xnor U3942 (N_3942,N_3683,N_3635);
nor U3943 (N_3943,N_3760,N_3828);
xnor U3944 (N_3944,N_3714,N_3805);
nor U3945 (N_3945,N_3775,N_3794);
and U3946 (N_3946,N_3814,N_3791);
or U3947 (N_3947,N_3885,N_3882);
nor U3948 (N_3948,N_3645,N_3842);
and U3949 (N_3949,N_3829,N_3726);
xor U3950 (N_3950,N_3708,N_3624);
xor U3951 (N_3951,N_3649,N_3689);
and U3952 (N_3952,N_3823,N_3826);
or U3953 (N_3953,N_3607,N_3776);
or U3954 (N_3954,N_3747,N_3854);
nand U3955 (N_3955,N_3718,N_3618);
or U3956 (N_3956,N_3638,N_3613);
and U3957 (N_3957,N_3803,N_3601);
nand U3958 (N_3958,N_3767,N_3673);
xor U3959 (N_3959,N_3615,N_3870);
and U3960 (N_3960,N_3872,N_3762);
or U3961 (N_3961,N_3755,N_3629);
and U3962 (N_3962,N_3614,N_3632);
or U3963 (N_3963,N_3616,N_3797);
xnor U3964 (N_3964,N_3725,N_3858);
xor U3965 (N_3965,N_3833,N_3891);
nor U3966 (N_3966,N_3671,N_3628);
or U3967 (N_3967,N_3824,N_3752);
or U3968 (N_3968,N_3600,N_3735);
nor U3969 (N_3969,N_3652,N_3765);
nand U3970 (N_3970,N_3660,N_3746);
and U3971 (N_3971,N_3818,N_3778);
or U3972 (N_3972,N_3686,N_3789);
nor U3973 (N_3973,N_3772,N_3773);
or U3974 (N_3974,N_3667,N_3697);
and U3975 (N_3975,N_3832,N_3850);
nor U3976 (N_3976,N_3790,N_3875);
and U3977 (N_3977,N_3728,N_3612);
xor U3978 (N_3978,N_3702,N_3807);
nor U3979 (N_3979,N_3820,N_3672);
xnor U3980 (N_3980,N_3692,N_3899);
and U3981 (N_3981,N_3750,N_3656);
xor U3982 (N_3982,N_3766,N_3757);
or U3983 (N_3983,N_3719,N_3694);
nand U3984 (N_3984,N_3779,N_3771);
or U3985 (N_3985,N_3887,N_3896);
and U3986 (N_3986,N_3758,N_3644);
and U3987 (N_3987,N_3761,N_3881);
xor U3988 (N_3988,N_3647,N_3666);
nand U3989 (N_3989,N_3654,N_3731);
xnor U3990 (N_3990,N_3886,N_3871);
nand U3991 (N_3991,N_3633,N_3650);
nand U3992 (N_3992,N_3659,N_3626);
nand U3993 (N_3993,N_3878,N_3696);
nor U3994 (N_3994,N_3670,N_3819);
xor U3995 (N_3995,N_3602,N_3816);
xor U3996 (N_3996,N_3657,N_3677);
nand U3997 (N_3997,N_3634,N_3608);
or U3998 (N_3998,N_3643,N_3732);
and U3999 (N_3999,N_3857,N_3868);
nand U4000 (N_4000,N_3641,N_3706);
nand U4001 (N_4001,N_3883,N_3780);
and U4002 (N_4002,N_3736,N_3841);
nand U4003 (N_4003,N_3711,N_3783);
xor U4004 (N_4004,N_3860,N_3727);
nand U4005 (N_4005,N_3713,N_3845);
and U4006 (N_4006,N_3754,N_3741);
and U4007 (N_4007,N_3604,N_3811);
and U4008 (N_4008,N_3804,N_3876);
xor U4009 (N_4009,N_3821,N_3756);
or U4010 (N_4010,N_3623,N_3838);
nor U4011 (N_4011,N_3737,N_3810);
nand U4012 (N_4012,N_3707,N_3753);
nand U4013 (N_4013,N_3764,N_3795);
or U4014 (N_4014,N_3890,N_3844);
nor U4015 (N_4015,N_3605,N_3716);
xnor U4016 (N_4016,N_3893,N_3620);
nor U4017 (N_4017,N_3817,N_3724);
nand U4018 (N_4018,N_3751,N_3788);
or U4019 (N_4019,N_3680,N_3717);
nor U4020 (N_4020,N_3894,N_3782);
and U4021 (N_4021,N_3639,N_3898);
and U4022 (N_4022,N_3715,N_3655);
xnor U4023 (N_4023,N_3691,N_3787);
or U4024 (N_4024,N_3710,N_3664);
nor U4025 (N_4025,N_3700,N_3625);
xnor U4026 (N_4026,N_3701,N_3809);
xnor U4027 (N_4027,N_3812,N_3669);
xnor U4028 (N_4028,N_3802,N_3705);
xor U4029 (N_4029,N_3801,N_3740);
nand U4030 (N_4030,N_3888,N_3658);
xor U4031 (N_4031,N_3874,N_3709);
nor U4032 (N_4032,N_3748,N_3674);
nand U4033 (N_4033,N_3685,N_3637);
xor U4034 (N_4034,N_3703,N_3781);
xnor U4035 (N_4035,N_3856,N_3763);
nor U4036 (N_4036,N_3792,N_3769);
or U4037 (N_4037,N_3682,N_3895);
nor U4038 (N_4038,N_3730,N_3759);
nand U4039 (N_4039,N_3855,N_3889);
xnor U4040 (N_4040,N_3675,N_3663);
xnor U4041 (N_4041,N_3786,N_3627);
nand U4042 (N_4042,N_3648,N_3822);
xnor U4043 (N_4043,N_3897,N_3873);
xor U4044 (N_4044,N_3852,N_3839);
or U4045 (N_4045,N_3848,N_3712);
or U4046 (N_4046,N_3676,N_3808);
and U4047 (N_4047,N_3646,N_3617);
and U4048 (N_4048,N_3836,N_3723);
xor U4049 (N_4049,N_3722,N_3668);
and U4050 (N_4050,N_3666,N_3853);
and U4051 (N_4051,N_3742,N_3656);
nor U4052 (N_4052,N_3623,N_3808);
xnor U4053 (N_4053,N_3750,N_3603);
nand U4054 (N_4054,N_3602,N_3649);
or U4055 (N_4055,N_3872,N_3601);
nand U4056 (N_4056,N_3881,N_3804);
and U4057 (N_4057,N_3750,N_3667);
or U4058 (N_4058,N_3681,N_3606);
or U4059 (N_4059,N_3618,N_3610);
or U4060 (N_4060,N_3797,N_3734);
and U4061 (N_4061,N_3800,N_3754);
xnor U4062 (N_4062,N_3806,N_3678);
xnor U4063 (N_4063,N_3634,N_3607);
and U4064 (N_4064,N_3650,N_3644);
nand U4065 (N_4065,N_3721,N_3835);
or U4066 (N_4066,N_3622,N_3687);
or U4067 (N_4067,N_3671,N_3633);
nor U4068 (N_4068,N_3842,N_3677);
xnor U4069 (N_4069,N_3675,N_3827);
xor U4070 (N_4070,N_3888,N_3777);
xnor U4071 (N_4071,N_3864,N_3827);
xor U4072 (N_4072,N_3731,N_3810);
or U4073 (N_4073,N_3602,N_3651);
and U4074 (N_4074,N_3759,N_3650);
or U4075 (N_4075,N_3737,N_3632);
and U4076 (N_4076,N_3861,N_3690);
nand U4077 (N_4077,N_3663,N_3635);
xnor U4078 (N_4078,N_3633,N_3838);
and U4079 (N_4079,N_3854,N_3722);
or U4080 (N_4080,N_3827,N_3892);
nor U4081 (N_4081,N_3664,N_3728);
xnor U4082 (N_4082,N_3834,N_3674);
xnor U4083 (N_4083,N_3791,N_3708);
xor U4084 (N_4084,N_3731,N_3841);
or U4085 (N_4085,N_3707,N_3643);
or U4086 (N_4086,N_3752,N_3655);
xnor U4087 (N_4087,N_3713,N_3890);
and U4088 (N_4088,N_3776,N_3775);
xor U4089 (N_4089,N_3823,N_3618);
xnor U4090 (N_4090,N_3724,N_3893);
nor U4091 (N_4091,N_3836,N_3641);
nor U4092 (N_4092,N_3807,N_3835);
or U4093 (N_4093,N_3807,N_3726);
nand U4094 (N_4094,N_3873,N_3737);
nand U4095 (N_4095,N_3839,N_3858);
or U4096 (N_4096,N_3871,N_3672);
xor U4097 (N_4097,N_3646,N_3865);
nand U4098 (N_4098,N_3810,N_3827);
xnor U4099 (N_4099,N_3768,N_3707);
nand U4100 (N_4100,N_3845,N_3874);
nor U4101 (N_4101,N_3607,N_3807);
xnor U4102 (N_4102,N_3617,N_3657);
and U4103 (N_4103,N_3610,N_3649);
nand U4104 (N_4104,N_3751,N_3745);
xnor U4105 (N_4105,N_3653,N_3826);
or U4106 (N_4106,N_3886,N_3642);
nand U4107 (N_4107,N_3678,N_3712);
and U4108 (N_4108,N_3759,N_3747);
or U4109 (N_4109,N_3690,N_3882);
and U4110 (N_4110,N_3766,N_3833);
xnor U4111 (N_4111,N_3828,N_3792);
nand U4112 (N_4112,N_3827,N_3729);
or U4113 (N_4113,N_3680,N_3741);
nor U4114 (N_4114,N_3725,N_3843);
and U4115 (N_4115,N_3786,N_3642);
nand U4116 (N_4116,N_3843,N_3803);
xor U4117 (N_4117,N_3687,N_3822);
and U4118 (N_4118,N_3613,N_3682);
and U4119 (N_4119,N_3704,N_3746);
and U4120 (N_4120,N_3848,N_3871);
nor U4121 (N_4121,N_3889,N_3619);
xor U4122 (N_4122,N_3880,N_3815);
xnor U4123 (N_4123,N_3883,N_3604);
or U4124 (N_4124,N_3691,N_3760);
or U4125 (N_4125,N_3629,N_3783);
nand U4126 (N_4126,N_3721,N_3717);
nand U4127 (N_4127,N_3694,N_3817);
xor U4128 (N_4128,N_3650,N_3768);
or U4129 (N_4129,N_3609,N_3677);
or U4130 (N_4130,N_3774,N_3634);
nand U4131 (N_4131,N_3714,N_3626);
xor U4132 (N_4132,N_3743,N_3794);
nand U4133 (N_4133,N_3688,N_3777);
nand U4134 (N_4134,N_3751,N_3671);
and U4135 (N_4135,N_3691,N_3790);
nor U4136 (N_4136,N_3617,N_3700);
nor U4137 (N_4137,N_3860,N_3719);
xor U4138 (N_4138,N_3701,N_3733);
nand U4139 (N_4139,N_3895,N_3701);
nand U4140 (N_4140,N_3657,N_3805);
nand U4141 (N_4141,N_3645,N_3776);
nor U4142 (N_4142,N_3681,N_3730);
or U4143 (N_4143,N_3860,N_3889);
nor U4144 (N_4144,N_3846,N_3883);
nand U4145 (N_4145,N_3707,N_3701);
or U4146 (N_4146,N_3655,N_3769);
xor U4147 (N_4147,N_3776,N_3838);
nand U4148 (N_4148,N_3674,N_3806);
xor U4149 (N_4149,N_3671,N_3776);
nand U4150 (N_4150,N_3806,N_3668);
nor U4151 (N_4151,N_3690,N_3838);
nand U4152 (N_4152,N_3821,N_3705);
nand U4153 (N_4153,N_3875,N_3877);
or U4154 (N_4154,N_3866,N_3687);
xnor U4155 (N_4155,N_3871,N_3669);
or U4156 (N_4156,N_3605,N_3756);
and U4157 (N_4157,N_3727,N_3695);
nand U4158 (N_4158,N_3708,N_3600);
or U4159 (N_4159,N_3757,N_3864);
nand U4160 (N_4160,N_3749,N_3880);
xnor U4161 (N_4161,N_3745,N_3721);
or U4162 (N_4162,N_3798,N_3763);
or U4163 (N_4163,N_3746,N_3884);
or U4164 (N_4164,N_3844,N_3779);
nor U4165 (N_4165,N_3774,N_3833);
nor U4166 (N_4166,N_3732,N_3824);
nor U4167 (N_4167,N_3831,N_3855);
or U4168 (N_4168,N_3837,N_3745);
xor U4169 (N_4169,N_3850,N_3705);
nand U4170 (N_4170,N_3847,N_3803);
xor U4171 (N_4171,N_3871,N_3888);
nor U4172 (N_4172,N_3898,N_3605);
or U4173 (N_4173,N_3728,N_3671);
nand U4174 (N_4174,N_3816,N_3677);
nor U4175 (N_4175,N_3646,N_3772);
nand U4176 (N_4176,N_3870,N_3757);
or U4177 (N_4177,N_3886,N_3639);
nand U4178 (N_4178,N_3828,N_3845);
and U4179 (N_4179,N_3813,N_3748);
xor U4180 (N_4180,N_3668,N_3739);
nor U4181 (N_4181,N_3869,N_3721);
nand U4182 (N_4182,N_3752,N_3839);
and U4183 (N_4183,N_3625,N_3805);
nand U4184 (N_4184,N_3784,N_3732);
xor U4185 (N_4185,N_3722,N_3850);
xnor U4186 (N_4186,N_3860,N_3802);
and U4187 (N_4187,N_3682,N_3837);
nand U4188 (N_4188,N_3639,N_3810);
xnor U4189 (N_4189,N_3878,N_3677);
xor U4190 (N_4190,N_3602,N_3851);
and U4191 (N_4191,N_3660,N_3616);
nor U4192 (N_4192,N_3631,N_3736);
and U4193 (N_4193,N_3609,N_3639);
nand U4194 (N_4194,N_3740,N_3891);
and U4195 (N_4195,N_3743,N_3842);
nand U4196 (N_4196,N_3668,N_3737);
and U4197 (N_4197,N_3811,N_3752);
and U4198 (N_4198,N_3623,N_3654);
or U4199 (N_4199,N_3859,N_3626);
and U4200 (N_4200,N_4085,N_4025);
or U4201 (N_4201,N_4178,N_4000);
and U4202 (N_4202,N_4096,N_4036);
nor U4203 (N_4203,N_4084,N_4071);
nand U4204 (N_4204,N_4080,N_3927);
nand U4205 (N_4205,N_4127,N_4068);
xor U4206 (N_4206,N_4179,N_4171);
or U4207 (N_4207,N_4141,N_4134);
or U4208 (N_4208,N_3999,N_4184);
or U4209 (N_4209,N_4046,N_4119);
and U4210 (N_4210,N_4149,N_4114);
nor U4211 (N_4211,N_4072,N_3964);
nor U4212 (N_4212,N_4166,N_4194);
or U4213 (N_4213,N_4031,N_4122);
nor U4214 (N_4214,N_4100,N_4181);
and U4215 (N_4215,N_4143,N_4117);
and U4216 (N_4216,N_3976,N_4125);
and U4217 (N_4217,N_4169,N_4094);
nor U4218 (N_4218,N_4073,N_4187);
or U4219 (N_4219,N_3955,N_4182);
nand U4220 (N_4220,N_4106,N_4019);
or U4221 (N_4221,N_4111,N_4067);
nor U4222 (N_4222,N_3941,N_3994);
nand U4223 (N_4223,N_3931,N_4093);
or U4224 (N_4224,N_4066,N_4157);
or U4225 (N_4225,N_3990,N_3909);
and U4226 (N_4226,N_4062,N_4042);
xnor U4227 (N_4227,N_4097,N_4156);
and U4228 (N_4228,N_4189,N_4022);
or U4229 (N_4229,N_4057,N_3950);
or U4230 (N_4230,N_3973,N_3956);
or U4231 (N_4231,N_4091,N_4095);
and U4232 (N_4232,N_4192,N_3977);
nor U4233 (N_4233,N_4045,N_3929);
and U4234 (N_4234,N_4105,N_4001);
nand U4235 (N_4235,N_3998,N_3922);
nand U4236 (N_4236,N_4015,N_3930);
xnor U4237 (N_4237,N_4152,N_4083);
xnor U4238 (N_4238,N_3982,N_4188);
xor U4239 (N_4239,N_4172,N_3985);
or U4240 (N_4240,N_4150,N_4033);
nor U4241 (N_4241,N_4089,N_4087);
nor U4242 (N_4242,N_4163,N_4136);
nand U4243 (N_4243,N_3932,N_4041);
or U4244 (N_4244,N_4060,N_4116);
xor U4245 (N_4245,N_3916,N_3901);
nand U4246 (N_4246,N_4173,N_4026);
nor U4247 (N_4247,N_4098,N_4162);
and U4248 (N_4248,N_4112,N_3962);
xor U4249 (N_4249,N_4047,N_3997);
and U4250 (N_4250,N_4040,N_3989);
and U4251 (N_4251,N_3900,N_3969);
nor U4252 (N_4252,N_4024,N_3904);
or U4253 (N_4253,N_4107,N_3960);
xnor U4254 (N_4254,N_4065,N_3942);
nor U4255 (N_4255,N_3965,N_4147);
and U4256 (N_4256,N_3943,N_4012);
nand U4257 (N_4257,N_4195,N_3970);
nor U4258 (N_4258,N_3972,N_4058);
and U4259 (N_4259,N_4014,N_4138);
or U4260 (N_4260,N_3984,N_4023);
nand U4261 (N_4261,N_4129,N_4011);
or U4262 (N_4262,N_4161,N_3907);
and U4263 (N_4263,N_4092,N_4109);
or U4264 (N_4264,N_3939,N_3987);
xnor U4265 (N_4265,N_4160,N_4034);
xor U4266 (N_4266,N_4153,N_4115);
or U4267 (N_4267,N_4020,N_3946);
and U4268 (N_4268,N_4102,N_3995);
and U4269 (N_4269,N_4076,N_4061);
nand U4270 (N_4270,N_3953,N_3958);
xnor U4271 (N_4271,N_3902,N_3938);
xor U4272 (N_4272,N_3912,N_3906);
nand U4273 (N_4273,N_4039,N_3934);
nand U4274 (N_4274,N_4177,N_3951);
nor U4275 (N_4275,N_4048,N_4159);
nand U4276 (N_4276,N_4032,N_3966);
xnor U4277 (N_4277,N_4104,N_3911);
or U4278 (N_4278,N_4035,N_4165);
xor U4279 (N_4279,N_3993,N_4146);
nand U4280 (N_4280,N_3979,N_4069);
or U4281 (N_4281,N_4140,N_3923);
xor U4282 (N_4282,N_4130,N_4135);
nor U4283 (N_4283,N_4082,N_3954);
nand U4284 (N_4284,N_4174,N_4155);
nor U4285 (N_4285,N_3991,N_4151);
nor U4286 (N_4286,N_4079,N_3986);
and U4287 (N_4287,N_3947,N_3957);
and U4288 (N_4288,N_4103,N_4144);
or U4289 (N_4289,N_3936,N_4108);
and U4290 (N_4290,N_4131,N_4145);
and U4291 (N_4291,N_4120,N_4081);
or U4292 (N_4292,N_3959,N_3915);
nand U4293 (N_4293,N_4123,N_4044);
or U4294 (N_4294,N_4137,N_4009);
xor U4295 (N_4295,N_4002,N_3980);
nand U4296 (N_4296,N_4049,N_4154);
nor U4297 (N_4297,N_3975,N_4043);
and U4298 (N_4298,N_4176,N_3918);
nand U4299 (N_4299,N_4168,N_3935);
or U4300 (N_4300,N_3952,N_4027);
or U4301 (N_4301,N_4158,N_3937);
and U4302 (N_4302,N_4050,N_4142);
and U4303 (N_4303,N_3945,N_4064);
and U4304 (N_4304,N_4053,N_4077);
nor U4305 (N_4305,N_4059,N_4010);
or U4306 (N_4306,N_3905,N_4196);
or U4307 (N_4307,N_4021,N_4055);
and U4308 (N_4308,N_4110,N_4126);
nor U4309 (N_4309,N_4075,N_4038);
nor U4310 (N_4310,N_4029,N_4088);
nor U4311 (N_4311,N_3961,N_4004);
and U4312 (N_4312,N_4132,N_3992);
and U4313 (N_4313,N_3971,N_3908);
and U4314 (N_4314,N_3917,N_3940);
and U4315 (N_4315,N_4052,N_3903);
and U4316 (N_4316,N_3920,N_4051);
xnor U4317 (N_4317,N_4028,N_3968);
nand U4318 (N_4318,N_3914,N_4128);
nand U4319 (N_4319,N_4005,N_4074);
nor U4320 (N_4320,N_3925,N_3926);
and U4321 (N_4321,N_3933,N_4164);
or U4322 (N_4322,N_4113,N_3967);
or U4323 (N_4323,N_4018,N_4078);
nor U4324 (N_4324,N_4006,N_3910);
xor U4325 (N_4325,N_4170,N_4118);
xnor U4326 (N_4326,N_4193,N_4199);
or U4327 (N_4327,N_4063,N_4016);
xor U4328 (N_4328,N_4090,N_4180);
xor U4329 (N_4329,N_3913,N_4124);
nand U4330 (N_4330,N_4007,N_3974);
xnor U4331 (N_4331,N_3988,N_4054);
xnor U4332 (N_4332,N_4185,N_4186);
or U4333 (N_4333,N_4175,N_4167);
xor U4334 (N_4334,N_4086,N_4037);
or U4335 (N_4335,N_4198,N_3983);
nand U4336 (N_4336,N_4121,N_4003);
xor U4337 (N_4337,N_3978,N_4030);
nor U4338 (N_4338,N_3928,N_4008);
and U4339 (N_4339,N_4017,N_4056);
nand U4340 (N_4340,N_4013,N_4101);
or U4341 (N_4341,N_4099,N_3944);
and U4342 (N_4342,N_4070,N_4183);
and U4343 (N_4343,N_3921,N_3981);
or U4344 (N_4344,N_3949,N_3996);
nor U4345 (N_4345,N_4139,N_3963);
xnor U4346 (N_4346,N_4197,N_4133);
or U4347 (N_4347,N_4191,N_4190);
xnor U4348 (N_4348,N_4148,N_3924);
xnor U4349 (N_4349,N_3948,N_3919);
xor U4350 (N_4350,N_4052,N_3988);
nor U4351 (N_4351,N_3985,N_3973);
and U4352 (N_4352,N_3960,N_3908);
nor U4353 (N_4353,N_3932,N_4147);
nand U4354 (N_4354,N_4144,N_3992);
nand U4355 (N_4355,N_4036,N_4103);
nor U4356 (N_4356,N_4136,N_4101);
nor U4357 (N_4357,N_3982,N_4167);
nand U4358 (N_4358,N_4022,N_4143);
or U4359 (N_4359,N_3947,N_3972);
or U4360 (N_4360,N_4084,N_3928);
nand U4361 (N_4361,N_4178,N_4134);
nor U4362 (N_4362,N_4101,N_3926);
xor U4363 (N_4363,N_4070,N_4153);
and U4364 (N_4364,N_3953,N_4141);
xor U4365 (N_4365,N_4059,N_4061);
and U4366 (N_4366,N_3990,N_3983);
nor U4367 (N_4367,N_4033,N_4040);
nand U4368 (N_4368,N_4031,N_4163);
nand U4369 (N_4369,N_3998,N_4020);
nand U4370 (N_4370,N_4015,N_3957);
and U4371 (N_4371,N_3920,N_4105);
nand U4372 (N_4372,N_4117,N_4071);
nand U4373 (N_4373,N_4000,N_4017);
nand U4374 (N_4374,N_3920,N_3957);
or U4375 (N_4375,N_4177,N_4030);
nand U4376 (N_4376,N_3987,N_4136);
nor U4377 (N_4377,N_4024,N_4020);
and U4378 (N_4378,N_3942,N_3954);
xor U4379 (N_4379,N_3905,N_4191);
nand U4380 (N_4380,N_4162,N_4027);
nor U4381 (N_4381,N_4160,N_4135);
or U4382 (N_4382,N_4111,N_4016);
and U4383 (N_4383,N_4038,N_4096);
nand U4384 (N_4384,N_4047,N_4198);
nand U4385 (N_4385,N_3940,N_3903);
or U4386 (N_4386,N_4020,N_4040);
or U4387 (N_4387,N_3942,N_4089);
and U4388 (N_4388,N_3965,N_4045);
or U4389 (N_4389,N_4105,N_4161);
or U4390 (N_4390,N_4138,N_3925);
nor U4391 (N_4391,N_4026,N_3906);
and U4392 (N_4392,N_4126,N_3947);
nor U4393 (N_4393,N_4023,N_4009);
or U4394 (N_4394,N_4072,N_4192);
and U4395 (N_4395,N_4158,N_3953);
and U4396 (N_4396,N_4001,N_4159);
xnor U4397 (N_4397,N_4047,N_3969);
nor U4398 (N_4398,N_4018,N_3976);
nor U4399 (N_4399,N_3997,N_4086);
or U4400 (N_4400,N_4125,N_3938);
nand U4401 (N_4401,N_4067,N_4116);
nand U4402 (N_4402,N_4162,N_4061);
xnor U4403 (N_4403,N_4063,N_4171);
nor U4404 (N_4404,N_4120,N_3925);
xnor U4405 (N_4405,N_4098,N_4171);
and U4406 (N_4406,N_4157,N_4112);
nand U4407 (N_4407,N_4009,N_3930);
xor U4408 (N_4408,N_4005,N_4040);
and U4409 (N_4409,N_4048,N_4042);
and U4410 (N_4410,N_3925,N_3987);
and U4411 (N_4411,N_4167,N_4126);
nand U4412 (N_4412,N_4029,N_4007);
nand U4413 (N_4413,N_3907,N_3922);
or U4414 (N_4414,N_3981,N_4182);
xor U4415 (N_4415,N_3912,N_4037);
and U4416 (N_4416,N_3922,N_4131);
nor U4417 (N_4417,N_4146,N_4110);
nand U4418 (N_4418,N_3925,N_4117);
or U4419 (N_4419,N_3912,N_3900);
xnor U4420 (N_4420,N_4062,N_4152);
nand U4421 (N_4421,N_4036,N_4089);
xor U4422 (N_4422,N_4079,N_4082);
nand U4423 (N_4423,N_3909,N_4129);
or U4424 (N_4424,N_3973,N_3976);
nand U4425 (N_4425,N_4113,N_3963);
and U4426 (N_4426,N_3990,N_3969);
and U4427 (N_4427,N_4020,N_3997);
nand U4428 (N_4428,N_4000,N_4072);
xor U4429 (N_4429,N_4077,N_4105);
nand U4430 (N_4430,N_4173,N_3923);
nor U4431 (N_4431,N_4033,N_3968);
and U4432 (N_4432,N_4159,N_4056);
nand U4433 (N_4433,N_4088,N_4114);
or U4434 (N_4434,N_4139,N_4002);
xnor U4435 (N_4435,N_3912,N_4081);
nor U4436 (N_4436,N_4117,N_4106);
and U4437 (N_4437,N_4193,N_4186);
nor U4438 (N_4438,N_4116,N_3939);
nand U4439 (N_4439,N_3968,N_4098);
and U4440 (N_4440,N_4046,N_3908);
and U4441 (N_4441,N_4082,N_3953);
nor U4442 (N_4442,N_3962,N_4080);
xor U4443 (N_4443,N_3905,N_4146);
nand U4444 (N_4444,N_4171,N_3999);
xor U4445 (N_4445,N_4081,N_4174);
nand U4446 (N_4446,N_4104,N_4119);
and U4447 (N_4447,N_4133,N_4043);
nand U4448 (N_4448,N_3970,N_4126);
or U4449 (N_4449,N_4125,N_3968);
and U4450 (N_4450,N_4060,N_4170);
and U4451 (N_4451,N_3921,N_3964);
nor U4452 (N_4452,N_3923,N_4109);
nand U4453 (N_4453,N_4119,N_4062);
and U4454 (N_4454,N_4015,N_4079);
or U4455 (N_4455,N_4067,N_4119);
nand U4456 (N_4456,N_3976,N_3938);
or U4457 (N_4457,N_3994,N_3937);
nand U4458 (N_4458,N_3936,N_4138);
or U4459 (N_4459,N_4088,N_4164);
xor U4460 (N_4460,N_4051,N_4069);
or U4461 (N_4461,N_4033,N_3995);
xor U4462 (N_4462,N_3974,N_4194);
nand U4463 (N_4463,N_3921,N_4194);
nand U4464 (N_4464,N_3986,N_4112);
nor U4465 (N_4465,N_4016,N_4056);
xnor U4466 (N_4466,N_4106,N_4015);
xor U4467 (N_4467,N_3945,N_3984);
nand U4468 (N_4468,N_3995,N_4120);
and U4469 (N_4469,N_4079,N_4004);
or U4470 (N_4470,N_4031,N_3947);
nor U4471 (N_4471,N_4036,N_4068);
and U4472 (N_4472,N_3969,N_4090);
xor U4473 (N_4473,N_4096,N_4016);
xnor U4474 (N_4474,N_4172,N_4178);
or U4475 (N_4475,N_4181,N_4143);
xor U4476 (N_4476,N_3940,N_4149);
nor U4477 (N_4477,N_4118,N_3974);
nand U4478 (N_4478,N_4027,N_4062);
xnor U4479 (N_4479,N_3967,N_4121);
xor U4480 (N_4480,N_4188,N_3917);
xnor U4481 (N_4481,N_4006,N_4031);
and U4482 (N_4482,N_3969,N_4018);
and U4483 (N_4483,N_4117,N_4042);
and U4484 (N_4484,N_3926,N_4026);
or U4485 (N_4485,N_4124,N_4069);
nor U4486 (N_4486,N_4161,N_4115);
xnor U4487 (N_4487,N_4190,N_4111);
nor U4488 (N_4488,N_4126,N_3986);
or U4489 (N_4489,N_4029,N_4167);
and U4490 (N_4490,N_4128,N_4146);
xnor U4491 (N_4491,N_4110,N_4025);
xnor U4492 (N_4492,N_4082,N_4095);
and U4493 (N_4493,N_4197,N_4128);
or U4494 (N_4494,N_4046,N_4129);
and U4495 (N_4495,N_4095,N_4003);
or U4496 (N_4496,N_4173,N_4175);
nor U4497 (N_4497,N_4115,N_4111);
or U4498 (N_4498,N_3927,N_4125);
xnor U4499 (N_4499,N_4144,N_4029);
nand U4500 (N_4500,N_4364,N_4307);
nor U4501 (N_4501,N_4204,N_4429);
xnor U4502 (N_4502,N_4409,N_4406);
and U4503 (N_4503,N_4487,N_4303);
xor U4504 (N_4504,N_4237,N_4338);
xor U4505 (N_4505,N_4371,N_4356);
and U4506 (N_4506,N_4256,N_4498);
and U4507 (N_4507,N_4434,N_4301);
and U4508 (N_4508,N_4347,N_4424);
nand U4509 (N_4509,N_4208,N_4431);
and U4510 (N_4510,N_4414,N_4390);
and U4511 (N_4511,N_4304,N_4355);
or U4512 (N_4512,N_4335,N_4393);
and U4513 (N_4513,N_4318,N_4278);
or U4514 (N_4514,N_4377,N_4324);
nand U4515 (N_4515,N_4437,N_4352);
nor U4516 (N_4516,N_4284,N_4286);
and U4517 (N_4517,N_4253,N_4398);
nor U4518 (N_4518,N_4403,N_4361);
and U4519 (N_4519,N_4485,N_4211);
and U4520 (N_4520,N_4354,N_4474);
or U4521 (N_4521,N_4220,N_4490);
and U4522 (N_4522,N_4225,N_4380);
and U4523 (N_4523,N_4357,N_4353);
and U4524 (N_4524,N_4410,N_4287);
nor U4525 (N_4525,N_4358,N_4374);
nand U4526 (N_4526,N_4486,N_4482);
nand U4527 (N_4527,N_4423,N_4389);
and U4528 (N_4528,N_4332,N_4293);
nand U4529 (N_4529,N_4362,N_4435);
nand U4530 (N_4530,N_4483,N_4239);
and U4531 (N_4531,N_4451,N_4306);
or U4532 (N_4532,N_4473,N_4452);
nand U4533 (N_4533,N_4213,N_4309);
nor U4534 (N_4534,N_4450,N_4396);
xor U4535 (N_4535,N_4432,N_4343);
nor U4536 (N_4536,N_4480,N_4238);
and U4537 (N_4537,N_4369,N_4310);
nand U4538 (N_4538,N_4242,N_4263);
xnor U4539 (N_4539,N_4367,N_4400);
or U4540 (N_4540,N_4265,N_4472);
nand U4541 (N_4541,N_4317,N_4234);
and U4542 (N_4542,N_4259,N_4210);
xnor U4543 (N_4543,N_4257,N_4385);
or U4544 (N_4544,N_4449,N_4202);
nor U4545 (N_4545,N_4228,N_4489);
nand U4546 (N_4546,N_4248,N_4296);
nor U4547 (N_4547,N_4288,N_4311);
and U4548 (N_4548,N_4496,N_4252);
nor U4549 (N_4549,N_4407,N_4333);
or U4550 (N_4550,N_4264,N_4408);
or U4551 (N_4551,N_4484,N_4391);
nand U4552 (N_4552,N_4281,N_4376);
nor U4553 (N_4553,N_4413,N_4491);
xor U4554 (N_4554,N_4440,N_4420);
or U4555 (N_4555,N_4471,N_4351);
nor U4556 (N_4556,N_4349,N_4241);
nand U4557 (N_4557,N_4326,N_4456);
xnor U4558 (N_4558,N_4399,N_4319);
or U4559 (N_4559,N_4282,N_4279);
xnor U4560 (N_4560,N_4442,N_4388);
nor U4561 (N_4561,N_4387,N_4422);
xnor U4562 (N_4562,N_4243,N_4274);
xor U4563 (N_4563,N_4383,N_4277);
or U4564 (N_4564,N_4322,N_4245);
nand U4565 (N_4565,N_4469,N_4497);
nor U4566 (N_4566,N_4478,N_4488);
nor U4567 (N_4567,N_4302,N_4395);
nor U4568 (N_4568,N_4365,N_4464);
nor U4569 (N_4569,N_4315,N_4381);
nor U4570 (N_4570,N_4405,N_4271);
xnor U4571 (N_4571,N_4305,N_4421);
nor U4572 (N_4572,N_4339,N_4350);
nor U4573 (N_4573,N_4217,N_4209);
xnor U4574 (N_4574,N_4240,N_4360);
nand U4575 (N_4575,N_4323,N_4341);
nor U4576 (N_4576,N_4227,N_4272);
nand U4577 (N_4577,N_4499,N_4261);
nor U4578 (N_4578,N_4445,N_4430);
and U4579 (N_4579,N_4379,N_4280);
and U4580 (N_4580,N_4222,N_4224);
xor U4581 (N_4581,N_4444,N_4461);
nor U4582 (N_4582,N_4329,N_4249);
nor U4583 (N_4583,N_4463,N_4330);
xnor U4584 (N_4584,N_4229,N_4459);
and U4585 (N_4585,N_4299,N_4251);
xor U4586 (N_4586,N_4466,N_4412);
nor U4587 (N_4587,N_4441,N_4223);
nor U4588 (N_4588,N_4453,N_4382);
nand U4589 (N_4589,N_4216,N_4266);
and U4590 (N_4590,N_4402,N_4269);
nand U4591 (N_4591,N_4260,N_4295);
xnor U4592 (N_4592,N_4439,N_4255);
or U4593 (N_4593,N_4460,N_4316);
and U4594 (N_4594,N_4207,N_4268);
xnor U4595 (N_4595,N_4425,N_4290);
and U4596 (N_4596,N_4378,N_4258);
xor U4597 (N_4597,N_4455,N_4447);
nand U4598 (N_4598,N_4458,N_4366);
nand U4599 (N_4599,N_4345,N_4344);
xor U4600 (N_4600,N_4298,N_4436);
xnor U4601 (N_4601,N_4334,N_4401);
nor U4602 (N_4602,N_4337,N_4415);
or U4603 (N_4603,N_4465,N_4203);
xnor U4604 (N_4604,N_4373,N_4416);
nand U4605 (N_4605,N_4419,N_4244);
and U4606 (N_4606,N_4481,N_4494);
or U4607 (N_4607,N_4200,N_4283);
xor U4608 (N_4608,N_4294,N_4340);
xnor U4609 (N_4609,N_4363,N_4325);
and U4610 (N_4610,N_4492,N_4384);
xor U4611 (N_4611,N_4254,N_4218);
nand U4612 (N_4612,N_4457,N_4433);
nand U4613 (N_4613,N_4285,N_4328);
nand U4614 (N_4614,N_4327,N_4336);
or U4615 (N_4615,N_4386,N_4411);
nor U4616 (N_4616,N_4308,N_4348);
xor U4617 (N_4617,N_4233,N_4443);
and U4618 (N_4618,N_4270,N_4292);
or U4619 (N_4619,N_4236,N_4477);
nor U4620 (N_4620,N_4428,N_4297);
or U4621 (N_4621,N_4247,N_4454);
nand U4622 (N_4622,N_4346,N_4314);
xnor U4623 (N_4623,N_4404,N_4215);
nor U4624 (N_4624,N_4375,N_4370);
or U4625 (N_4625,N_4462,N_4475);
or U4626 (N_4626,N_4418,N_4246);
nand U4627 (N_4627,N_4275,N_4392);
or U4628 (N_4628,N_4262,N_4212);
nor U4629 (N_4629,N_4493,N_4446);
and U4630 (N_4630,N_4470,N_4467);
nor U4631 (N_4631,N_4313,N_4267);
nand U4632 (N_4632,N_4226,N_4479);
or U4633 (N_4633,N_4201,N_4331);
nor U4634 (N_4634,N_4219,N_4232);
nor U4635 (N_4635,N_4438,N_4320);
xor U4636 (N_4636,N_4426,N_4231);
xnor U4637 (N_4637,N_4476,N_4250);
nand U4638 (N_4638,N_4394,N_4289);
xor U4639 (N_4639,N_4417,N_4427);
nor U4640 (N_4640,N_4291,N_4359);
nand U4641 (N_4641,N_4312,N_4495);
or U4642 (N_4642,N_4321,N_4230);
nor U4643 (N_4643,N_4342,N_4448);
and U4644 (N_4644,N_4273,N_4205);
and U4645 (N_4645,N_4221,N_4214);
or U4646 (N_4646,N_4300,N_4206);
or U4647 (N_4647,N_4397,N_4276);
nand U4648 (N_4648,N_4372,N_4368);
nand U4649 (N_4649,N_4235,N_4468);
nor U4650 (N_4650,N_4441,N_4318);
and U4651 (N_4651,N_4308,N_4438);
xor U4652 (N_4652,N_4436,N_4472);
nor U4653 (N_4653,N_4425,N_4223);
nand U4654 (N_4654,N_4388,N_4218);
or U4655 (N_4655,N_4219,N_4285);
xor U4656 (N_4656,N_4486,N_4329);
or U4657 (N_4657,N_4468,N_4367);
and U4658 (N_4658,N_4481,N_4476);
nor U4659 (N_4659,N_4304,N_4279);
nand U4660 (N_4660,N_4424,N_4287);
xor U4661 (N_4661,N_4272,N_4309);
nand U4662 (N_4662,N_4297,N_4471);
nand U4663 (N_4663,N_4219,N_4307);
and U4664 (N_4664,N_4226,N_4311);
xnor U4665 (N_4665,N_4241,N_4239);
xnor U4666 (N_4666,N_4375,N_4450);
nand U4667 (N_4667,N_4490,N_4463);
or U4668 (N_4668,N_4286,N_4320);
or U4669 (N_4669,N_4415,N_4335);
nand U4670 (N_4670,N_4378,N_4364);
and U4671 (N_4671,N_4475,N_4348);
nand U4672 (N_4672,N_4217,N_4299);
nand U4673 (N_4673,N_4239,N_4463);
or U4674 (N_4674,N_4319,N_4246);
nor U4675 (N_4675,N_4345,N_4355);
and U4676 (N_4676,N_4242,N_4365);
nor U4677 (N_4677,N_4475,N_4332);
nand U4678 (N_4678,N_4375,N_4386);
nand U4679 (N_4679,N_4349,N_4441);
nand U4680 (N_4680,N_4252,N_4281);
xnor U4681 (N_4681,N_4425,N_4267);
or U4682 (N_4682,N_4346,N_4273);
and U4683 (N_4683,N_4467,N_4320);
xnor U4684 (N_4684,N_4365,N_4496);
and U4685 (N_4685,N_4299,N_4467);
or U4686 (N_4686,N_4261,N_4388);
or U4687 (N_4687,N_4322,N_4304);
xnor U4688 (N_4688,N_4257,N_4375);
or U4689 (N_4689,N_4465,N_4282);
or U4690 (N_4690,N_4446,N_4273);
nor U4691 (N_4691,N_4240,N_4320);
nand U4692 (N_4692,N_4234,N_4348);
nand U4693 (N_4693,N_4272,N_4422);
xor U4694 (N_4694,N_4231,N_4311);
or U4695 (N_4695,N_4264,N_4328);
xnor U4696 (N_4696,N_4458,N_4494);
and U4697 (N_4697,N_4273,N_4429);
nor U4698 (N_4698,N_4274,N_4235);
or U4699 (N_4699,N_4466,N_4202);
or U4700 (N_4700,N_4333,N_4238);
or U4701 (N_4701,N_4255,N_4355);
nor U4702 (N_4702,N_4387,N_4390);
xnor U4703 (N_4703,N_4362,N_4476);
or U4704 (N_4704,N_4357,N_4317);
and U4705 (N_4705,N_4257,N_4245);
and U4706 (N_4706,N_4307,N_4420);
or U4707 (N_4707,N_4404,N_4339);
or U4708 (N_4708,N_4461,N_4394);
nand U4709 (N_4709,N_4354,N_4488);
or U4710 (N_4710,N_4339,N_4211);
and U4711 (N_4711,N_4415,N_4329);
nor U4712 (N_4712,N_4204,N_4416);
and U4713 (N_4713,N_4276,N_4444);
nor U4714 (N_4714,N_4430,N_4298);
or U4715 (N_4715,N_4271,N_4227);
nor U4716 (N_4716,N_4232,N_4223);
or U4717 (N_4717,N_4201,N_4490);
nand U4718 (N_4718,N_4250,N_4375);
or U4719 (N_4719,N_4252,N_4310);
xnor U4720 (N_4720,N_4228,N_4255);
nor U4721 (N_4721,N_4463,N_4337);
nand U4722 (N_4722,N_4369,N_4284);
nor U4723 (N_4723,N_4482,N_4282);
and U4724 (N_4724,N_4360,N_4238);
nor U4725 (N_4725,N_4401,N_4262);
and U4726 (N_4726,N_4376,N_4458);
nand U4727 (N_4727,N_4401,N_4359);
or U4728 (N_4728,N_4390,N_4393);
xor U4729 (N_4729,N_4490,N_4477);
nand U4730 (N_4730,N_4305,N_4253);
and U4731 (N_4731,N_4241,N_4403);
and U4732 (N_4732,N_4485,N_4288);
and U4733 (N_4733,N_4283,N_4408);
xnor U4734 (N_4734,N_4246,N_4317);
and U4735 (N_4735,N_4266,N_4433);
xor U4736 (N_4736,N_4367,N_4309);
nor U4737 (N_4737,N_4318,N_4455);
nand U4738 (N_4738,N_4291,N_4234);
nand U4739 (N_4739,N_4403,N_4233);
nand U4740 (N_4740,N_4473,N_4234);
nand U4741 (N_4741,N_4484,N_4329);
and U4742 (N_4742,N_4294,N_4227);
or U4743 (N_4743,N_4233,N_4358);
and U4744 (N_4744,N_4366,N_4290);
and U4745 (N_4745,N_4414,N_4233);
nand U4746 (N_4746,N_4497,N_4454);
nor U4747 (N_4747,N_4364,N_4499);
xor U4748 (N_4748,N_4261,N_4418);
or U4749 (N_4749,N_4202,N_4298);
and U4750 (N_4750,N_4305,N_4440);
nand U4751 (N_4751,N_4356,N_4283);
nor U4752 (N_4752,N_4342,N_4439);
or U4753 (N_4753,N_4297,N_4294);
nor U4754 (N_4754,N_4369,N_4308);
and U4755 (N_4755,N_4481,N_4245);
nand U4756 (N_4756,N_4371,N_4219);
nand U4757 (N_4757,N_4440,N_4433);
or U4758 (N_4758,N_4350,N_4361);
or U4759 (N_4759,N_4433,N_4248);
or U4760 (N_4760,N_4322,N_4218);
xor U4761 (N_4761,N_4260,N_4479);
nand U4762 (N_4762,N_4359,N_4271);
and U4763 (N_4763,N_4420,N_4497);
nor U4764 (N_4764,N_4267,N_4391);
nand U4765 (N_4765,N_4319,N_4455);
nor U4766 (N_4766,N_4417,N_4405);
or U4767 (N_4767,N_4399,N_4253);
or U4768 (N_4768,N_4333,N_4403);
nand U4769 (N_4769,N_4347,N_4258);
nand U4770 (N_4770,N_4315,N_4386);
nor U4771 (N_4771,N_4310,N_4269);
or U4772 (N_4772,N_4326,N_4337);
xor U4773 (N_4773,N_4341,N_4254);
xor U4774 (N_4774,N_4443,N_4276);
and U4775 (N_4775,N_4224,N_4341);
xnor U4776 (N_4776,N_4442,N_4334);
and U4777 (N_4777,N_4384,N_4396);
nor U4778 (N_4778,N_4317,N_4443);
nor U4779 (N_4779,N_4343,N_4356);
nand U4780 (N_4780,N_4496,N_4316);
nand U4781 (N_4781,N_4380,N_4406);
nand U4782 (N_4782,N_4411,N_4395);
nor U4783 (N_4783,N_4302,N_4388);
xor U4784 (N_4784,N_4302,N_4366);
or U4785 (N_4785,N_4404,N_4383);
nand U4786 (N_4786,N_4307,N_4335);
or U4787 (N_4787,N_4201,N_4431);
and U4788 (N_4788,N_4343,N_4315);
and U4789 (N_4789,N_4439,N_4413);
and U4790 (N_4790,N_4496,N_4319);
or U4791 (N_4791,N_4313,N_4264);
or U4792 (N_4792,N_4221,N_4417);
and U4793 (N_4793,N_4423,N_4495);
xnor U4794 (N_4794,N_4443,N_4231);
and U4795 (N_4795,N_4466,N_4305);
or U4796 (N_4796,N_4266,N_4380);
and U4797 (N_4797,N_4294,N_4496);
and U4798 (N_4798,N_4384,N_4436);
and U4799 (N_4799,N_4280,N_4378);
xor U4800 (N_4800,N_4699,N_4715);
and U4801 (N_4801,N_4544,N_4705);
or U4802 (N_4802,N_4640,N_4508);
or U4803 (N_4803,N_4737,N_4696);
and U4804 (N_4804,N_4525,N_4761);
nor U4805 (N_4805,N_4746,N_4659);
or U4806 (N_4806,N_4764,N_4643);
nor U4807 (N_4807,N_4636,N_4686);
and U4808 (N_4808,N_4721,N_4528);
nand U4809 (N_4809,N_4533,N_4654);
and U4810 (N_4810,N_4778,N_4688);
and U4811 (N_4811,N_4673,N_4552);
and U4812 (N_4812,N_4790,N_4542);
nand U4813 (N_4813,N_4700,N_4719);
nand U4814 (N_4814,N_4671,N_4617);
nor U4815 (N_4815,N_4515,N_4590);
xnor U4816 (N_4816,N_4510,N_4585);
xor U4817 (N_4817,N_4720,N_4663);
nor U4818 (N_4818,N_4537,N_4651);
nand U4819 (N_4819,N_4685,N_4546);
nand U4820 (N_4820,N_4511,N_4574);
and U4821 (N_4821,N_4777,N_4607);
and U4822 (N_4822,N_4750,N_4539);
nor U4823 (N_4823,N_4763,N_4577);
or U4824 (N_4824,N_4524,N_4744);
nor U4825 (N_4825,N_4759,N_4770);
xnor U4826 (N_4826,N_4691,N_4677);
and U4827 (N_4827,N_4587,N_4704);
xnor U4828 (N_4828,N_4765,N_4712);
or U4829 (N_4829,N_4598,N_4603);
xnor U4830 (N_4830,N_4583,N_4683);
or U4831 (N_4831,N_4772,N_4707);
xor U4832 (N_4832,N_4516,N_4664);
or U4833 (N_4833,N_4675,N_4788);
xor U4834 (N_4834,N_4612,N_4754);
nor U4835 (N_4835,N_4626,N_4566);
nor U4836 (N_4836,N_4655,N_4536);
nand U4837 (N_4837,N_4735,N_4678);
and U4838 (N_4838,N_4624,N_4580);
or U4839 (N_4839,N_4798,N_4676);
nand U4840 (N_4840,N_4782,N_4710);
xor U4841 (N_4841,N_4596,N_4581);
or U4842 (N_4842,N_4733,N_4632);
or U4843 (N_4843,N_4792,N_4668);
and U4844 (N_4844,N_4775,N_4556);
xnor U4845 (N_4845,N_4523,N_4797);
and U4846 (N_4846,N_4535,N_4589);
or U4847 (N_4847,N_4698,N_4512);
nor U4848 (N_4848,N_4505,N_4785);
and U4849 (N_4849,N_4743,N_4689);
xnor U4850 (N_4850,N_4711,N_4600);
xor U4851 (N_4851,N_4760,N_4594);
xor U4852 (N_4852,N_4681,N_4554);
nor U4853 (N_4853,N_4749,N_4724);
nand U4854 (N_4854,N_4503,N_4540);
and U4855 (N_4855,N_4783,N_4672);
nor U4856 (N_4856,N_4570,N_4674);
nand U4857 (N_4857,N_4709,N_4627);
nand U4858 (N_4858,N_4738,N_4670);
or U4859 (N_4859,N_4758,N_4684);
nand U4860 (N_4860,N_4679,N_4722);
xnor U4861 (N_4861,N_4747,N_4530);
nor U4862 (N_4862,N_4693,N_4717);
nand U4863 (N_4863,N_4774,N_4543);
nand U4864 (N_4864,N_4648,N_4652);
xor U4865 (N_4865,N_4610,N_4776);
and U4866 (N_4866,N_4514,N_4784);
xnor U4867 (N_4867,N_4517,N_4615);
nor U4868 (N_4868,N_4661,N_4755);
xor U4869 (N_4869,N_4529,N_4628);
nand U4870 (N_4870,N_4527,N_4729);
and U4871 (N_4871,N_4616,N_4572);
nand U4872 (N_4872,N_4713,N_4584);
nand U4873 (N_4873,N_4504,N_4521);
and U4874 (N_4874,N_4740,N_4642);
and U4875 (N_4875,N_4682,N_4562);
xor U4876 (N_4876,N_4519,N_4762);
and U4877 (N_4877,N_4773,N_4509);
nand U4878 (N_4878,N_4622,N_4706);
or U4879 (N_4879,N_4561,N_4791);
nand U4880 (N_4880,N_4796,N_4518);
or U4881 (N_4881,N_4752,N_4701);
nor U4882 (N_4882,N_4520,N_4599);
or U4883 (N_4883,N_4500,N_4613);
nand U4884 (N_4884,N_4633,N_4656);
and U4885 (N_4885,N_4732,N_4559);
nor U4886 (N_4886,N_4578,N_4526);
xnor U4887 (N_4887,N_4799,N_4634);
nand U4888 (N_4888,N_4601,N_4767);
xnor U4889 (N_4889,N_4639,N_4629);
nor U4890 (N_4890,N_4567,N_4553);
xnor U4891 (N_4891,N_4786,N_4619);
nor U4892 (N_4892,N_4502,N_4532);
xnor U4893 (N_4893,N_4669,N_4573);
nand U4894 (N_4894,N_4662,N_4625);
and U4895 (N_4895,N_4692,N_4565);
nor U4896 (N_4896,N_4702,N_4728);
and U4897 (N_4897,N_4793,N_4649);
or U4898 (N_4898,N_4576,N_4555);
nor U4899 (N_4899,N_4522,N_4769);
and U4900 (N_4900,N_4575,N_4795);
nor U4901 (N_4901,N_4725,N_4507);
nor U4902 (N_4902,N_4534,N_4551);
and U4903 (N_4903,N_4731,N_4726);
nand U4904 (N_4904,N_4779,N_4660);
and U4905 (N_4905,N_4501,N_4736);
nor U4906 (N_4906,N_4653,N_4579);
xor U4907 (N_4907,N_4637,N_4694);
or U4908 (N_4908,N_4753,N_4739);
or U4909 (N_4909,N_4650,N_4593);
xnor U4910 (N_4910,N_4716,N_4586);
or U4911 (N_4911,N_4563,N_4568);
nand U4912 (N_4912,N_4560,N_4550);
and U4913 (N_4913,N_4794,N_4757);
nand U4914 (N_4914,N_4549,N_4611);
or U4915 (N_4915,N_4620,N_4766);
xor U4916 (N_4916,N_4741,N_4771);
and U4917 (N_4917,N_4690,N_4582);
xnor U4918 (N_4918,N_4703,N_4609);
nor U4919 (N_4919,N_4789,N_4548);
and U4920 (N_4920,N_4768,N_4606);
and U4921 (N_4921,N_4571,N_4541);
xor U4922 (N_4922,N_4621,N_4695);
nor U4923 (N_4923,N_4730,N_4645);
nand U4924 (N_4924,N_4602,N_4742);
nand U4925 (N_4925,N_4646,N_4748);
xnor U4926 (N_4926,N_4513,N_4638);
and U4927 (N_4927,N_4605,N_4635);
and U4928 (N_4928,N_4745,N_4708);
and U4929 (N_4929,N_4564,N_4595);
nand U4930 (N_4930,N_4658,N_4734);
xnor U4931 (N_4931,N_4618,N_4588);
and U4932 (N_4932,N_4641,N_4697);
xnor U4933 (N_4933,N_4647,N_4558);
nand U4934 (N_4934,N_4667,N_4718);
and U4935 (N_4935,N_4557,N_4756);
and U4936 (N_4936,N_4591,N_4657);
nand U4937 (N_4937,N_4723,N_4630);
or U4938 (N_4938,N_4608,N_4751);
xnor U4939 (N_4939,N_4592,N_4644);
or U4940 (N_4940,N_4780,N_4547);
and U4941 (N_4941,N_4614,N_4631);
xnor U4942 (N_4942,N_4538,N_4665);
xor U4943 (N_4943,N_4781,N_4727);
and U4944 (N_4944,N_4680,N_4506);
and U4945 (N_4945,N_4569,N_4545);
xor U4946 (N_4946,N_4666,N_4787);
or U4947 (N_4947,N_4623,N_4597);
and U4948 (N_4948,N_4687,N_4714);
xnor U4949 (N_4949,N_4531,N_4604);
or U4950 (N_4950,N_4691,N_4588);
xnor U4951 (N_4951,N_4742,N_4604);
nor U4952 (N_4952,N_4643,N_4502);
xnor U4953 (N_4953,N_4589,N_4752);
or U4954 (N_4954,N_4736,N_4614);
or U4955 (N_4955,N_4735,N_4756);
xnor U4956 (N_4956,N_4520,N_4501);
xor U4957 (N_4957,N_4748,N_4627);
or U4958 (N_4958,N_4748,N_4707);
and U4959 (N_4959,N_4733,N_4594);
xnor U4960 (N_4960,N_4555,N_4754);
nor U4961 (N_4961,N_4700,N_4784);
xnor U4962 (N_4962,N_4573,N_4783);
xor U4963 (N_4963,N_4614,N_4564);
xor U4964 (N_4964,N_4733,N_4527);
nor U4965 (N_4965,N_4742,N_4504);
and U4966 (N_4966,N_4761,N_4512);
xnor U4967 (N_4967,N_4714,N_4590);
xnor U4968 (N_4968,N_4517,N_4634);
and U4969 (N_4969,N_4607,N_4685);
xor U4970 (N_4970,N_4718,N_4635);
xnor U4971 (N_4971,N_4748,N_4559);
nand U4972 (N_4972,N_4614,N_4629);
nor U4973 (N_4973,N_4784,N_4512);
or U4974 (N_4974,N_4749,N_4799);
and U4975 (N_4975,N_4615,N_4770);
or U4976 (N_4976,N_4663,N_4666);
or U4977 (N_4977,N_4578,N_4507);
xor U4978 (N_4978,N_4612,N_4650);
and U4979 (N_4979,N_4600,N_4773);
nor U4980 (N_4980,N_4540,N_4721);
and U4981 (N_4981,N_4572,N_4700);
nor U4982 (N_4982,N_4668,N_4635);
or U4983 (N_4983,N_4793,N_4597);
and U4984 (N_4984,N_4623,N_4585);
nand U4985 (N_4985,N_4794,N_4691);
xor U4986 (N_4986,N_4677,N_4553);
nor U4987 (N_4987,N_4728,N_4621);
nand U4988 (N_4988,N_4547,N_4647);
xor U4989 (N_4989,N_4583,N_4736);
xor U4990 (N_4990,N_4737,N_4505);
nand U4991 (N_4991,N_4567,N_4562);
nand U4992 (N_4992,N_4662,N_4697);
and U4993 (N_4993,N_4541,N_4791);
nand U4994 (N_4994,N_4532,N_4530);
and U4995 (N_4995,N_4791,N_4669);
nor U4996 (N_4996,N_4690,N_4503);
and U4997 (N_4997,N_4624,N_4646);
xnor U4998 (N_4998,N_4735,N_4646);
xor U4999 (N_4999,N_4572,N_4766);
or U5000 (N_5000,N_4712,N_4608);
and U5001 (N_5001,N_4512,N_4751);
nor U5002 (N_5002,N_4657,N_4768);
nand U5003 (N_5003,N_4735,N_4786);
nand U5004 (N_5004,N_4667,N_4769);
xnor U5005 (N_5005,N_4674,N_4684);
and U5006 (N_5006,N_4756,N_4653);
xnor U5007 (N_5007,N_4617,N_4501);
nand U5008 (N_5008,N_4597,N_4756);
nand U5009 (N_5009,N_4797,N_4507);
xor U5010 (N_5010,N_4513,N_4659);
or U5011 (N_5011,N_4799,N_4727);
xor U5012 (N_5012,N_4729,N_4598);
and U5013 (N_5013,N_4796,N_4564);
or U5014 (N_5014,N_4649,N_4755);
and U5015 (N_5015,N_4704,N_4567);
nand U5016 (N_5016,N_4708,N_4633);
or U5017 (N_5017,N_4750,N_4764);
nor U5018 (N_5018,N_4550,N_4688);
nor U5019 (N_5019,N_4662,N_4562);
and U5020 (N_5020,N_4683,N_4532);
or U5021 (N_5021,N_4681,N_4515);
or U5022 (N_5022,N_4538,N_4638);
nor U5023 (N_5023,N_4775,N_4725);
and U5024 (N_5024,N_4774,N_4708);
and U5025 (N_5025,N_4594,N_4677);
xor U5026 (N_5026,N_4657,N_4580);
or U5027 (N_5027,N_4600,N_4725);
xnor U5028 (N_5028,N_4714,N_4692);
or U5029 (N_5029,N_4735,N_4576);
nand U5030 (N_5030,N_4687,N_4731);
nand U5031 (N_5031,N_4747,N_4562);
and U5032 (N_5032,N_4709,N_4510);
nor U5033 (N_5033,N_4731,N_4655);
and U5034 (N_5034,N_4512,N_4745);
xnor U5035 (N_5035,N_4529,N_4755);
and U5036 (N_5036,N_4730,N_4650);
nor U5037 (N_5037,N_4710,N_4704);
or U5038 (N_5038,N_4766,N_4559);
xnor U5039 (N_5039,N_4504,N_4711);
nor U5040 (N_5040,N_4590,N_4587);
xnor U5041 (N_5041,N_4642,N_4684);
nand U5042 (N_5042,N_4717,N_4638);
nand U5043 (N_5043,N_4689,N_4742);
nand U5044 (N_5044,N_4675,N_4568);
or U5045 (N_5045,N_4687,N_4735);
or U5046 (N_5046,N_4560,N_4593);
xnor U5047 (N_5047,N_4710,N_4712);
and U5048 (N_5048,N_4508,N_4701);
and U5049 (N_5049,N_4763,N_4541);
or U5050 (N_5050,N_4641,N_4632);
or U5051 (N_5051,N_4738,N_4736);
xnor U5052 (N_5052,N_4581,N_4646);
xnor U5053 (N_5053,N_4626,N_4690);
xor U5054 (N_5054,N_4530,N_4579);
and U5055 (N_5055,N_4551,N_4664);
nand U5056 (N_5056,N_4778,N_4550);
nor U5057 (N_5057,N_4608,N_4643);
xnor U5058 (N_5058,N_4750,N_4642);
nand U5059 (N_5059,N_4609,N_4599);
nand U5060 (N_5060,N_4663,N_4556);
nor U5061 (N_5061,N_4686,N_4570);
and U5062 (N_5062,N_4552,N_4628);
nand U5063 (N_5063,N_4678,N_4552);
nor U5064 (N_5064,N_4690,N_4557);
or U5065 (N_5065,N_4607,N_4761);
and U5066 (N_5066,N_4795,N_4748);
and U5067 (N_5067,N_4626,N_4561);
and U5068 (N_5068,N_4719,N_4588);
or U5069 (N_5069,N_4778,N_4558);
nor U5070 (N_5070,N_4707,N_4768);
xnor U5071 (N_5071,N_4556,N_4649);
xor U5072 (N_5072,N_4670,N_4751);
nand U5073 (N_5073,N_4529,N_4636);
and U5074 (N_5074,N_4519,N_4671);
nor U5075 (N_5075,N_4694,N_4664);
nor U5076 (N_5076,N_4662,N_4517);
xnor U5077 (N_5077,N_4531,N_4586);
and U5078 (N_5078,N_4524,N_4574);
or U5079 (N_5079,N_4765,N_4778);
nor U5080 (N_5080,N_4731,N_4554);
xor U5081 (N_5081,N_4784,N_4528);
nor U5082 (N_5082,N_4611,N_4702);
or U5083 (N_5083,N_4517,N_4632);
or U5084 (N_5084,N_4744,N_4569);
and U5085 (N_5085,N_4616,N_4584);
xor U5086 (N_5086,N_4509,N_4785);
nand U5087 (N_5087,N_4713,N_4615);
nor U5088 (N_5088,N_4644,N_4796);
nand U5089 (N_5089,N_4724,N_4707);
xnor U5090 (N_5090,N_4739,N_4656);
and U5091 (N_5091,N_4584,N_4746);
xnor U5092 (N_5092,N_4665,N_4655);
nand U5093 (N_5093,N_4714,N_4655);
or U5094 (N_5094,N_4529,N_4505);
nor U5095 (N_5095,N_4560,N_4611);
or U5096 (N_5096,N_4541,N_4614);
nor U5097 (N_5097,N_4556,N_4786);
xnor U5098 (N_5098,N_4753,N_4573);
nor U5099 (N_5099,N_4658,N_4567);
or U5100 (N_5100,N_5029,N_5023);
nor U5101 (N_5101,N_4862,N_4841);
nand U5102 (N_5102,N_5008,N_5077);
nand U5103 (N_5103,N_5045,N_4812);
and U5104 (N_5104,N_4849,N_4840);
or U5105 (N_5105,N_4961,N_4853);
or U5106 (N_5106,N_4984,N_5080);
nor U5107 (N_5107,N_4877,N_5047);
nand U5108 (N_5108,N_5020,N_4960);
nor U5109 (N_5109,N_4972,N_4871);
nor U5110 (N_5110,N_5078,N_4934);
nor U5111 (N_5111,N_4810,N_4935);
nand U5112 (N_5112,N_4887,N_4855);
and U5113 (N_5113,N_4918,N_4832);
or U5114 (N_5114,N_4967,N_4857);
and U5115 (N_5115,N_4833,N_4915);
or U5116 (N_5116,N_4842,N_4808);
or U5117 (N_5117,N_5017,N_5057);
nor U5118 (N_5118,N_4920,N_4912);
nand U5119 (N_5119,N_4968,N_5025);
nand U5120 (N_5120,N_5084,N_4979);
and U5121 (N_5121,N_4991,N_5031);
nand U5122 (N_5122,N_4989,N_4927);
and U5123 (N_5123,N_4928,N_4925);
xor U5124 (N_5124,N_5033,N_4802);
nor U5125 (N_5125,N_4894,N_4942);
and U5126 (N_5126,N_5085,N_4873);
and U5127 (N_5127,N_5083,N_5000);
nor U5128 (N_5128,N_5005,N_4936);
nor U5129 (N_5129,N_4924,N_4962);
and U5130 (N_5130,N_4910,N_5019);
xor U5131 (N_5131,N_4969,N_5087);
xor U5132 (N_5132,N_4819,N_4868);
xor U5133 (N_5133,N_4815,N_5004);
and U5134 (N_5134,N_4801,N_5046);
and U5135 (N_5135,N_5093,N_4823);
or U5136 (N_5136,N_5054,N_4870);
xnor U5137 (N_5137,N_4803,N_5011);
xor U5138 (N_5138,N_4839,N_4957);
xnor U5139 (N_5139,N_4985,N_4933);
nand U5140 (N_5140,N_4838,N_4986);
and U5141 (N_5141,N_5039,N_4913);
and U5142 (N_5142,N_5060,N_5079);
xor U5143 (N_5143,N_4916,N_4847);
and U5144 (N_5144,N_4923,N_5052);
xnor U5145 (N_5145,N_4947,N_4848);
nor U5146 (N_5146,N_4906,N_4882);
nor U5147 (N_5147,N_4902,N_5071);
nor U5148 (N_5148,N_5050,N_4948);
xor U5149 (N_5149,N_4945,N_4814);
and U5150 (N_5150,N_4834,N_5044);
xnor U5151 (N_5151,N_5055,N_4858);
xnor U5152 (N_5152,N_4951,N_4852);
and U5153 (N_5153,N_4930,N_5028);
nand U5154 (N_5154,N_5049,N_4931);
or U5155 (N_5155,N_4982,N_5068);
nand U5156 (N_5156,N_5073,N_4946);
nor U5157 (N_5157,N_4828,N_5099);
nand U5158 (N_5158,N_5014,N_4876);
nor U5159 (N_5159,N_5059,N_5081);
and U5160 (N_5160,N_4922,N_5074);
xnor U5161 (N_5161,N_4835,N_4896);
or U5162 (N_5162,N_4900,N_4937);
nor U5163 (N_5163,N_4864,N_5037);
nor U5164 (N_5164,N_4919,N_5036);
nor U5165 (N_5165,N_4890,N_4996);
nor U5166 (N_5166,N_4820,N_4859);
xnor U5167 (N_5167,N_5026,N_4867);
or U5168 (N_5168,N_4953,N_5065);
or U5169 (N_5169,N_4821,N_4895);
xnor U5170 (N_5170,N_4880,N_4813);
nor U5171 (N_5171,N_4949,N_4939);
nor U5172 (N_5172,N_5058,N_4805);
nor U5173 (N_5173,N_4964,N_4863);
and U5174 (N_5174,N_4889,N_5072);
xor U5175 (N_5175,N_5034,N_4917);
and U5176 (N_5176,N_5013,N_4909);
or U5177 (N_5177,N_4892,N_4943);
nand U5178 (N_5178,N_5091,N_4999);
and U5179 (N_5179,N_5003,N_4975);
nand U5180 (N_5180,N_4845,N_4811);
nor U5181 (N_5181,N_4959,N_4884);
nor U5182 (N_5182,N_5062,N_4965);
nor U5183 (N_5183,N_4977,N_4897);
nor U5184 (N_5184,N_4970,N_5086);
nand U5185 (N_5185,N_5043,N_4978);
or U5186 (N_5186,N_5067,N_4854);
xnor U5187 (N_5187,N_4874,N_4866);
or U5188 (N_5188,N_5010,N_4872);
and U5189 (N_5189,N_4994,N_4893);
nor U5190 (N_5190,N_4908,N_4954);
or U5191 (N_5191,N_4829,N_5092);
and U5192 (N_5192,N_4851,N_5040);
or U5193 (N_5193,N_5070,N_4941);
or U5194 (N_5194,N_5030,N_5076);
or U5195 (N_5195,N_4888,N_5096);
xnor U5196 (N_5196,N_4983,N_4881);
and U5197 (N_5197,N_4886,N_5056);
xnor U5198 (N_5198,N_4990,N_5038);
nand U5199 (N_5199,N_5098,N_4879);
nor U5200 (N_5200,N_5018,N_4827);
or U5201 (N_5201,N_5035,N_4804);
nor U5202 (N_5202,N_4809,N_4997);
nand U5203 (N_5203,N_4825,N_4966);
nor U5204 (N_5204,N_5094,N_4800);
nor U5205 (N_5205,N_5082,N_4891);
xnor U5206 (N_5206,N_4958,N_4806);
nand U5207 (N_5207,N_4903,N_5088);
nor U5208 (N_5208,N_4911,N_4818);
or U5209 (N_5209,N_5090,N_5007);
nand U5210 (N_5210,N_4981,N_4831);
xnor U5211 (N_5211,N_4846,N_4861);
nor U5212 (N_5212,N_4901,N_4971);
xor U5213 (N_5213,N_4869,N_4988);
or U5214 (N_5214,N_4952,N_4944);
xnor U5215 (N_5215,N_4998,N_4976);
nand U5216 (N_5216,N_5027,N_4907);
or U5217 (N_5217,N_5006,N_4899);
xor U5218 (N_5218,N_4824,N_4837);
or U5219 (N_5219,N_4843,N_5015);
xnor U5220 (N_5220,N_4844,N_4940);
and U5221 (N_5221,N_4932,N_4905);
xnor U5222 (N_5222,N_5022,N_4875);
and U5223 (N_5223,N_5061,N_5095);
and U5224 (N_5224,N_5016,N_5021);
or U5225 (N_5225,N_5012,N_5075);
or U5226 (N_5226,N_4987,N_5053);
nor U5227 (N_5227,N_5069,N_5002);
xor U5228 (N_5228,N_5051,N_4980);
or U5229 (N_5229,N_4865,N_5032);
nor U5230 (N_5230,N_4878,N_4830);
or U5231 (N_5231,N_4995,N_4914);
nand U5232 (N_5232,N_4836,N_4974);
nand U5233 (N_5233,N_4883,N_5048);
nand U5234 (N_5234,N_4822,N_4807);
or U5235 (N_5235,N_4950,N_5063);
nand U5236 (N_5236,N_4898,N_4963);
nand U5237 (N_5237,N_5009,N_5001);
nor U5238 (N_5238,N_4816,N_4929);
nand U5239 (N_5239,N_5089,N_5024);
xor U5240 (N_5240,N_4885,N_5066);
nand U5241 (N_5241,N_4850,N_5064);
nor U5242 (N_5242,N_4993,N_4992);
and U5243 (N_5243,N_4955,N_4904);
and U5244 (N_5244,N_5041,N_4817);
xor U5245 (N_5245,N_4926,N_5097);
and U5246 (N_5246,N_4973,N_4856);
or U5247 (N_5247,N_4860,N_4921);
or U5248 (N_5248,N_4956,N_4938);
and U5249 (N_5249,N_4826,N_5042);
and U5250 (N_5250,N_5065,N_5053);
or U5251 (N_5251,N_4952,N_4923);
xnor U5252 (N_5252,N_5024,N_5018);
and U5253 (N_5253,N_4814,N_5065);
xor U5254 (N_5254,N_5060,N_4881);
xor U5255 (N_5255,N_5000,N_4862);
xor U5256 (N_5256,N_4973,N_4855);
or U5257 (N_5257,N_5015,N_5092);
or U5258 (N_5258,N_4915,N_4836);
nand U5259 (N_5259,N_4866,N_5044);
or U5260 (N_5260,N_4940,N_4831);
nand U5261 (N_5261,N_4831,N_4851);
nor U5262 (N_5262,N_4835,N_5030);
or U5263 (N_5263,N_4983,N_4848);
nor U5264 (N_5264,N_4848,N_5061);
nand U5265 (N_5265,N_4838,N_4839);
nor U5266 (N_5266,N_4868,N_4967);
xnor U5267 (N_5267,N_4855,N_4935);
or U5268 (N_5268,N_4992,N_4818);
nand U5269 (N_5269,N_5072,N_4837);
nand U5270 (N_5270,N_4943,N_4926);
xnor U5271 (N_5271,N_4993,N_4931);
or U5272 (N_5272,N_4921,N_4850);
nor U5273 (N_5273,N_5044,N_4922);
nor U5274 (N_5274,N_4843,N_4826);
xnor U5275 (N_5275,N_4865,N_5064);
xor U5276 (N_5276,N_5028,N_4985);
or U5277 (N_5277,N_5020,N_4946);
nand U5278 (N_5278,N_4860,N_5066);
xnor U5279 (N_5279,N_5008,N_4815);
nand U5280 (N_5280,N_4837,N_5076);
xor U5281 (N_5281,N_5092,N_4856);
and U5282 (N_5282,N_4804,N_4869);
and U5283 (N_5283,N_4854,N_4832);
nand U5284 (N_5284,N_4810,N_4846);
nand U5285 (N_5285,N_4965,N_4828);
nor U5286 (N_5286,N_4886,N_4934);
nand U5287 (N_5287,N_4860,N_4917);
or U5288 (N_5288,N_4933,N_4858);
or U5289 (N_5289,N_4809,N_5031);
nor U5290 (N_5290,N_4959,N_4868);
nor U5291 (N_5291,N_4835,N_4946);
nand U5292 (N_5292,N_4833,N_5069);
or U5293 (N_5293,N_4871,N_4912);
or U5294 (N_5294,N_4946,N_5013);
nand U5295 (N_5295,N_4989,N_5047);
and U5296 (N_5296,N_4842,N_4802);
nand U5297 (N_5297,N_4949,N_4980);
nand U5298 (N_5298,N_4909,N_4815);
and U5299 (N_5299,N_5026,N_5034);
or U5300 (N_5300,N_4911,N_5041);
and U5301 (N_5301,N_4975,N_5019);
nand U5302 (N_5302,N_4928,N_4836);
xor U5303 (N_5303,N_5009,N_4958);
and U5304 (N_5304,N_4850,N_4879);
xnor U5305 (N_5305,N_4899,N_5078);
xnor U5306 (N_5306,N_4867,N_5017);
xnor U5307 (N_5307,N_4830,N_4870);
or U5308 (N_5308,N_4822,N_4970);
nand U5309 (N_5309,N_4892,N_5083);
nor U5310 (N_5310,N_5042,N_4810);
or U5311 (N_5311,N_5045,N_4929);
and U5312 (N_5312,N_5046,N_4829);
nand U5313 (N_5313,N_5012,N_5027);
nor U5314 (N_5314,N_5068,N_4952);
and U5315 (N_5315,N_5087,N_4881);
xor U5316 (N_5316,N_4928,N_4972);
and U5317 (N_5317,N_4943,N_5036);
and U5318 (N_5318,N_5082,N_4888);
nor U5319 (N_5319,N_4833,N_4842);
nor U5320 (N_5320,N_4918,N_4962);
nand U5321 (N_5321,N_4907,N_5014);
nor U5322 (N_5322,N_4879,N_4950);
and U5323 (N_5323,N_5027,N_5026);
and U5324 (N_5324,N_4873,N_5013);
nor U5325 (N_5325,N_4993,N_5077);
and U5326 (N_5326,N_5070,N_4894);
nand U5327 (N_5327,N_5046,N_5042);
nor U5328 (N_5328,N_4942,N_4838);
or U5329 (N_5329,N_5046,N_4845);
and U5330 (N_5330,N_5061,N_5094);
nor U5331 (N_5331,N_4928,N_4961);
and U5332 (N_5332,N_4924,N_4896);
xnor U5333 (N_5333,N_4861,N_5044);
nor U5334 (N_5334,N_4825,N_5088);
or U5335 (N_5335,N_4874,N_5087);
and U5336 (N_5336,N_4885,N_4810);
or U5337 (N_5337,N_5052,N_5069);
xor U5338 (N_5338,N_4837,N_4968);
nor U5339 (N_5339,N_4855,N_4989);
nor U5340 (N_5340,N_4927,N_4954);
or U5341 (N_5341,N_4951,N_4860);
nor U5342 (N_5342,N_5075,N_4813);
and U5343 (N_5343,N_4971,N_4816);
xnor U5344 (N_5344,N_5018,N_4933);
nor U5345 (N_5345,N_4891,N_4997);
or U5346 (N_5346,N_5069,N_4849);
xor U5347 (N_5347,N_5012,N_4899);
and U5348 (N_5348,N_4945,N_5003);
xor U5349 (N_5349,N_5071,N_5011);
or U5350 (N_5350,N_4910,N_4944);
and U5351 (N_5351,N_4910,N_4848);
xor U5352 (N_5352,N_4814,N_4892);
xnor U5353 (N_5353,N_4876,N_4941);
or U5354 (N_5354,N_4950,N_4981);
nor U5355 (N_5355,N_4925,N_4901);
xnor U5356 (N_5356,N_5057,N_4890);
xnor U5357 (N_5357,N_4853,N_4897);
and U5358 (N_5358,N_4893,N_5062);
xnor U5359 (N_5359,N_4861,N_5001);
xor U5360 (N_5360,N_4885,N_5039);
or U5361 (N_5361,N_4961,N_5045);
nand U5362 (N_5362,N_5015,N_4864);
nand U5363 (N_5363,N_5013,N_4843);
xor U5364 (N_5364,N_4912,N_5061);
or U5365 (N_5365,N_4860,N_4960);
or U5366 (N_5366,N_4949,N_4826);
and U5367 (N_5367,N_4929,N_5005);
and U5368 (N_5368,N_4883,N_4941);
and U5369 (N_5369,N_5010,N_4954);
or U5370 (N_5370,N_4807,N_4963);
xor U5371 (N_5371,N_4808,N_4995);
and U5372 (N_5372,N_4887,N_4950);
nor U5373 (N_5373,N_4806,N_5031);
nor U5374 (N_5374,N_4949,N_4811);
and U5375 (N_5375,N_5077,N_4949);
xnor U5376 (N_5376,N_5013,N_5085);
xnor U5377 (N_5377,N_5099,N_4931);
and U5378 (N_5378,N_5006,N_5095);
xnor U5379 (N_5379,N_4984,N_5006);
and U5380 (N_5380,N_5081,N_4855);
nand U5381 (N_5381,N_4903,N_5031);
nand U5382 (N_5382,N_4910,N_4985);
nor U5383 (N_5383,N_4973,N_4851);
and U5384 (N_5384,N_4858,N_4932);
xnor U5385 (N_5385,N_4917,N_4985);
or U5386 (N_5386,N_5072,N_5028);
xnor U5387 (N_5387,N_4991,N_5038);
nand U5388 (N_5388,N_5080,N_5076);
or U5389 (N_5389,N_4958,N_5031);
xnor U5390 (N_5390,N_5099,N_5071);
xnor U5391 (N_5391,N_4895,N_4862);
nor U5392 (N_5392,N_4849,N_4926);
xor U5393 (N_5393,N_4962,N_5035);
nor U5394 (N_5394,N_4902,N_5002);
xor U5395 (N_5395,N_4803,N_4913);
nand U5396 (N_5396,N_5032,N_4867);
nor U5397 (N_5397,N_4862,N_5095);
and U5398 (N_5398,N_4977,N_5078);
and U5399 (N_5399,N_4926,N_5002);
nor U5400 (N_5400,N_5364,N_5367);
xnor U5401 (N_5401,N_5337,N_5100);
xnor U5402 (N_5402,N_5300,N_5108);
or U5403 (N_5403,N_5395,N_5210);
and U5404 (N_5404,N_5199,N_5320);
xnor U5405 (N_5405,N_5250,N_5135);
xnor U5406 (N_5406,N_5336,N_5278);
xnor U5407 (N_5407,N_5370,N_5277);
or U5408 (N_5408,N_5228,N_5276);
nand U5409 (N_5409,N_5376,N_5114);
xnor U5410 (N_5410,N_5350,N_5357);
xnor U5411 (N_5411,N_5154,N_5251);
xor U5412 (N_5412,N_5183,N_5379);
nor U5413 (N_5413,N_5227,N_5174);
xnor U5414 (N_5414,N_5230,N_5391);
nand U5415 (N_5415,N_5241,N_5368);
and U5416 (N_5416,N_5188,N_5116);
xor U5417 (N_5417,N_5329,N_5328);
xnor U5418 (N_5418,N_5206,N_5127);
and U5419 (N_5419,N_5349,N_5198);
nand U5420 (N_5420,N_5211,N_5342);
nor U5421 (N_5421,N_5104,N_5148);
and U5422 (N_5422,N_5190,N_5345);
nor U5423 (N_5423,N_5222,N_5132);
nor U5424 (N_5424,N_5352,N_5255);
nor U5425 (N_5425,N_5217,N_5141);
nand U5426 (N_5426,N_5205,N_5166);
or U5427 (N_5427,N_5207,N_5121);
xnor U5428 (N_5428,N_5363,N_5149);
nor U5429 (N_5429,N_5196,N_5373);
nor U5430 (N_5430,N_5134,N_5112);
and U5431 (N_5431,N_5189,N_5312);
nand U5432 (N_5432,N_5371,N_5197);
nor U5433 (N_5433,N_5351,N_5202);
or U5434 (N_5434,N_5283,N_5332);
nor U5435 (N_5435,N_5101,N_5378);
xnor U5436 (N_5436,N_5284,N_5331);
nand U5437 (N_5437,N_5225,N_5268);
nand U5438 (N_5438,N_5272,N_5171);
nand U5439 (N_5439,N_5327,N_5374);
xor U5440 (N_5440,N_5263,N_5247);
and U5441 (N_5441,N_5167,N_5309);
nand U5442 (N_5442,N_5246,N_5296);
or U5443 (N_5443,N_5220,N_5229);
xnor U5444 (N_5444,N_5181,N_5308);
nor U5445 (N_5445,N_5216,N_5117);
xor U5446 (N_5446,N_5269,N_5209);
xnor U5447 (N_5447,N_5143,N_5281);
and U5448 (N_5448,N_5297,N_5318);
and U5449 (N_5449,N_5129,N_5261);
nand U5450 (N_5450,N_5338,N_5260);
or U5451 (N_5451,N_5393,N_5356);
and U5452 (N_5452,N_5285,N_5106);
or U5453 (N_5453,N_5124,N_5287);
nand U5454 (N_5454,N_5194,N_5235);
nand U5455 (N_5455,N_5324,N_5311);
nor U5456 (N_5456,N_5214,N_5282);
or U5457 (N_5457,N_5265,N_5257);
or U5458 (N_5458,N_5170,N_5301);
and U5459 (N_5459,N_5271,N_5240);
nor U5460 (N_5460,N_5314,N_5133);
or U5461 (N_5461,N_5292,N_5145);
and U5462 (N_5462,N_5245,N_5153);
or U5463 (N_5463,N_5142,N_5102);
or U5464 (N_5464,N_5361,N_5175);
or U5465 (N_5465,N_5258,N_5299);
xnor U5466 (N_5466,N_5270,N_5128);
xnor U5467 (N_5467,N_5172,N_5176);
or U5468 (N_5468,N_5192,N_5321);
xnor U5469 (N_5469,N_5182,N_5138);
and U5470 (N_5470,N_5390,N_5253);
or U5471 (N_5471,N_5146,N_5115);
nand U5472 (N_5472,N_5159,N_5111);
and U5473 (N_5473,N_5291,N_5103);
xnor U5474 (N_5474,N_5243,N_5305);
nor U5475 (N_5475,N_5160,N_5215);
nand U5476 (N_5476,N_5262,N_5334);
nand U5477 (N_5477,N_5392,N_5204);
and U5478 (N_5478,N_5226,N_5218);
nand U5479 (N_5479,N_5120,N_5273);
and U5480 (N_5480,N_5274,N_5335);
and U5481 (N_5481,N_5286,N_5168);
nand U5482 (N_5482,N_5213,N_5252);
nor U5483 (N_5483,N_5122,N_5293);
nand U5484 (N_5484,N_5303,N_5231);
nor U5485 (N_5485,N_5169,N_5396);
and U5486 (N_5486,N_5399,N_5372);
nand U5487 (N_5487,N_5178,N_5302);
or U5488 (N_5488,N_5359,N_5158);
nor U5489 (N_5489,N_5144,N_5185);
xor U5490 (N_5490,N_5389,N_5341);
xor U5491 (N_5491,N_5137,N_5326);
and U5492 (N_5492,N_5295,N_5173);
or U5493 (N_5493,N_5307,N_5223);
nand U5494 (N_5494,N_5152,N_5256);
or U5495 (N_5495,N_5203,N_5369);
and U5496 (N_5496,N_5343,N_5346);
or U5497 (N_5497,N_5384,N_5164);
nand U5498 (N_5498,N_5322,N_5239);
and U5499 (N_5499,N_5306,N_5360);
xor U5500 (N_5500,N_5304,N_5165);
nand U5501 (N_5501,N_5157,N_5386);
xor U5502 (N_5502,N_5219,N_5348);
xor U5503 (N_5503,N_5130,N_5319);
nor U5504 (N_5504,N_5366,N_5248);
xor U5505 (N_5505,N_5186,N_5313);
and U5506 (N_5506,N_5195,N_5325);
and U5507 (N_5507,N_5234,N_5200);
or U5508 (N_5508,N_5344,N_5381);
xnor U5509 (N_5509,N_5236,N_5151);
or U5510 (N_5510,N_5394,N_5289);
nand U5511 (N_5511,N_5290,N_5275);
and U5512 (N_5512,N_5347,N_5339);
xor U5513 (N_5513,N_5315,N_5310);
xor U5514 (N_5514,N_5125,N_5237);
and U5515 (N_5515,N_5212,N_5266);
xnor U5516 (N_5516,N_5377,N_5398);
nand U5517 (N_5517,N_5267,N_5387);
nor U5518 (N_5518,N_5340,N_5354);
xor U5519 (N_5519,N_5233,N_5288);
and U5520 (N_5520,N_5208,N_5232);
nand U5521 (N_5521,N_5110,N_5259);
xor U5522 (N_5522,N_5355,N_5221);
and U5523 (N_5523,N_5358,N_5107);
or U5524 (N_5524,N_5383,N_5123);
nor U5525 (N_5525,N_5244,N_5388);
and U5526 (N_5526,N_5380,N_5375);
nor U5527 (N_5527,N_5242,N_5140);
nor U5528 (N_5528,N_5254,N_5298);
nor U5529 (N_5529,N_5113,N_5131);
nand U5530 (N_5530,N_5179,N_5353);
nand U5531 (N_5531,N_5119,N_5316);
or U5532 (N_5532,N_5184,N_5264);
nand U5533 (N_5533,N_5162,N_5155);
xor U5534 (N_5534,N_5330,N_5280);
and U5535 (N_5535,N_5294,N_5150);
nor U5536 (N_5536,N_5187,N_5397);
nor U5537 (N_5537,N_5191,N_5362);
xor U5538 (N_5538,N_5163,N_5333);
xnor U5539 (N_5539,N_5224,N_5382);
nor U5540 (N_5540,N_5118,N_5109);
nand U5541 (N_5541,N_5139,N_5156);
and U5542 (N_5542,N_5201,N_5177);
xnor U5543 (N_5543,N_5279,N_5105);
nor U5544 (N_5544,N_5249,N_5385);
or U5545 (N_5545,N_5323,N_5136);
or U5546 (N_5546,N_5238,N_5365);
nor U5547 (N_5547,N_5193,N_5147);
nand U5548 (N_5548,N_5180,N_5126);
or U5549 (N_5549,N_5317,N_5161);
nor U5550 (N_5550,N_5299,N_5135);
nand U5551 (N_5551,N_5368,N_5324);
nand U5552 (N_5552,N_5238,N_5309);
nand U5553 (N_5553,N_5330,N_5292);
nand U5554 (N_5554,N_5390,N_5281);
and U5555 (N_5555,N_5268,N_5377);
xor U5556 (N_5556,N_5320,N_5107);
nand U5557 (N_5557,N_5390,N_5166);
xnor U5558 (N_5558,N_5325,N_5155);
xor U5559 (N_5559,N_5226,N_5148);
nor U5560 (N_5560,N_5356,N_5220);
or U5561 (N_5561,N_5116,N_5245);
nor U5562 (N_5562,N_5338,N_5103);
xnor U5563 (N_5563,N_5236,N_5385);
nor U5564 (N_5564,N_5163,N_5387);
or U5565 (N_5565,N_5119,N_5229);
or U5566 (N_5566,N_5230,N_5197);
nor U5567 (N_5567,N_5233,N_5394);
nand U5568 (N_5568,N_5369,N_5158);
xnor U5569 (N_5569,N_5367,N_5308);
nand U5570 (N_5570,N_5103,N_5223);
nand U5571 (N_5571,N_5104,N_5276);
or U5572 (N_5572,N_5204,N_5368);
or U5573 (N_5573,N_5334,N_5291);
nand U5574 (N_5574,N_5360,N_5373);
nand U5575 (N_5575,N_5179,N_5396);
nand U5576 (N_5576,N_5143,N_5248);
nor U5577 (N_5577,N_5181,N_5275);
nand U5578 (N_5578,N_5171,N_5250);
nor U5579 (N_5579,N_5276,N_5336);
xor U5580 (N_5580,N_5324,N_5298);
nand U5581 (N_5581,N_5221,N_5333);
xor U5582 (N_5582,N_5201,N_5233);
xnor U5583 (N_5583,N_5381,N_5383);
xor U5584 (N_5584,N_5184,N_5171);
nor U5585 (N_5585,N_5283,N_5398);
and U5586 (N_5586,N_5341,N_5224);
or U5587 (N_5587,N_5179,N_5286);
xor U5588 (N_5588,N_5382,N_5118);
or U5589 (N_5589,N_5176,N_5134);
nor U5590 (N_5590,N_5390,N_5329);
and U5591 (N_5591,N_5283,N_5180);
xnor U5592 (N_5592,N_5147,N_5227);
xnor U5593 (N_5593,N_5340,N_5129);
or U5594 (N_5594,N_5133,N_5168);
xor U5595 (N_5595,N_5301,N_5204);
or U5596 (N_5596,N_5329,N_5122);
nand U5597 (N_5597,N_5351,N_5184);
xor U5598 (N_5598,N_5288,N_5360);
and U5599 (N_5599,N_5111,N_5258);
xnor U5600 (N_5600,N_5195,N_5282);
or U5601 (N_5601,N_5231,N_5369);
xor U5602 (N_5602,N_5114,N_5124);
or U5603 (N_5603,N_5248,N_5317);
or U5604 (N_5604,N_5120,N_5141);
nand U5605 (N_5605,N_5197,N_5185);
and U5606 (N_5606,N_5135,N_5268);
or U5607 (N_5607,N_5385,N_5367);
nor U5608 (N_5608,N_5150,N_5159);
nand U5609 (N_5609,N_5382,N_5174);
or U5610 (N_5610,N_5115,N_5202);
or U5611 (N_5611,N_5395,N_5365);
nor U5612 (N_5612,N_5329,N_5194);
nand U5613 (N_5613,N_5386,N_5154);
xnor U5614 (N_5614,N_5171,N_5202);
nand U5615 (N_5615,N_5275,N_5217);
or U5616 (N_5616,N_5169,N_5193);
nand U5617 (N_5617,N_5352,N_5277);
and U5618 (N_5618,N_5318,N_5235);
nand U5619 (N_5619,N_5141,N_5290);
nand U5620 (N_5620,N_5325,N_5341);
nand U5621 (N_5621,N_5352,N_5212);
nand U5622 (N_5622,N_5206,N_5399);
nand U5623 (N_5623,N_5287,N_5104);
and U5624 (N_5624,N_5221,N_5155);
or U5625 (N_5625,N_5110,N_5303);
nor U5626 (N_5626,N_5274,N_5105);
xnor U5627 (N_5627,N_5373,N_5399);
and U5628 (N_5628,N_5132,N_5300);
and U5629 (N_5629,N_5299,N_5267);
xor U5630 (N_5630,N_5352,N_5282);
and U5631 (N_5631,N_5194,N_5133);
nor U5632 (N_5632,N_5176,N_5237);
nand U5633 (N_5633,N_5232,N_5340);
nand U5634 (N_5634,N_5258,N_5202);
nand U5635 (N_5635,N_5368,N_5375);
nor U5636 (N_5636,N_5315,N_5279);
and U5637 (N_5637,N_5180,N_5115);
or U5638 (N_5638,N_5152,N_5156);
or U5639 (N_5639,N_5254,N_5204);
or U5640 (N_5640,N_5150,N_5181);
nand U5641 (N_5641,N_5266,N_5293);
and U5642 (N_5642,N_5329,N_5316);
xor U5643 (N_5643,N_5350,N_5249);
and U5644 (N_5644,N_5116,N_5266);
and U5645 (N_5645,N_5189,N_5393);
nand U5646 (N_5646,N_5159,N_5290);
nor U5647 (N_5647,N_5341,N_5309);
or U5648 (N_5648,N_5175,N_5380);
and U5649 (N_5649,N_5184,N_5303);
nor U5650 (N_5650,N_5315,N_5294);
or U5651 (N_5651,N_5118,N_5339);
or U5652 (N_5652,N_5291,N_5185);
nand U5653 (N_5653,N_5345,N_5350);
or U5654 (N_5654,N_5331,N_5273);
and U5655 (N_5655,N_5145,N_5345);
nand U5656 (N_5656,N_5339,N_5233);
or U5657 (N_5657,N_5389,N_5368);
xor U5658 (N_5658,N_5114,N_5394);
nor U5659 (N_5659,N_5247,N_5297);
xnor U5660 (N_5660,N_5145,N_5190);
and U5661 (N_5661,N_5384,N_5168);
nand U5662 (N_5662,N_5350,N_5145);
nor U5663 (N_5663,N_5350,N_5110);
nand U5664 (N_5664,N_5235,N_5122);
and U5665 (N_5665,N_5171,N_5121);
and U5666 (N_5666,N_5367,N_5207);
nor U5667 (N_5667,N_5238,N_5130);
or U5668 (N_5668,N_5106,N_5261);
xnor U5669 (N_5669,N_5196,N_5399);
xor U5670 (N_5670,N_5199,N_5345);
or U5671 (N_5671,N_5207,N_5240);
xnor U5672 (N_5672,N_5331,N_5138);
nand U5673 (N_5673,N_5382,N_5214);
nor U5674 (N_5674,N_5313,N_5306);
and U5675 (N_5675,N_5312,N_5134);
nor U5676 (N_5676,N_5195,N_5308);
nor U5677 (N_5677,N_5236,N_5253);
and U5678 (N_5678,N_5279,N_5213);
nand U5679 (N_5679,N_5242,N_5151);
xnor U5680 (N_5680,N_5140,N_5224);
nor U5681 (N_5681,N_5187,N_5341);
or U5682 (N_5682,N_5275,N_5236);
xor U5683 (N_5683,N_5223,N_5283);
or U5684 (N_5684,N_5399,N_5232);
and U5685 (N_5685,N_5230,N_5148);
nor U5686 (N_5686,N_5230,N_5116);
xnor U5687 (N_5687,N_5192,N_5143);
nand U5688 (N_5688,N_5175,N_5281);
and U5689 (N_5689,N_5199,N_5230);
or U5690 (N_5690,N_5121,N_5313);
xor U5691 (N_5691,N_5282,N_5151);
or U5692 (N_5692,N_5162,N_5267);
or U5693 (N_5693,N_5367,N_5265);
nor U5694 (N_5694,N_5292,N_5109);
and U5695 (N_5695,N_5181,N_5210);
nor U5696 (N_5696,N_5363,N_5380);
nor U5697 (N_5697,N_5133,N_5213);
nor U5698 (N_5698,N_5386,N_5236);
nand U5699 (N_5699,N_5317,N_5141);
and U5700 (N_5700,N_5450,N_5686);
or U5701 (N_5701,N_5586,N_5648);
or U5702 (N_5702,N_5410,N_5479);
nor U5703 (N_5703,N_5453,N_5423);
xor U5704 (N_5704,N_5670,N_5432);
or U5705 (N_5705,N_5455,N_5692);
xor U5706 (N_5706,N_5641,N_5654);
or U5707 (N_5707,N_5611,N_5445);
or U5708 (N_5708,N_5467,N_5605);
and U5709 (N_5709,N_5638,N_5663);
or U5710 (N_5710,N_5464,N_5606);
and U5711 (N_5711,N_5409,N_5458);
xnor U5712 (N_5712,N_5540,N_5497);
or U5713 (N_5713,N_5647,N_5521);
xnor U5714 (N_5714,N_5619,N_5678);
or U5715 (N_5715,N_5646,N_5413);
nor U5716 (N_5716,N_5463,N_5472);
and U5717 (N_5717,N_5543,N_5471);
xor U5718 (N_5718,N_5695,N_5486);
or U5719 (N_5719,N_5673,N_5633);
xor U5720 (N_5720,N_5443,N_5515);
xnor U5721 (N_5721,N_5563,N_5542);
nor U5722 (N_5722,N_5579,N_5444);
or U5723 (N_5723,N_5532,N_5434);
xnor U5724 (N_5724,N_5545,N_5672);
and U5725 (N_5725,N_5671,N_5488);
nand U5726 (N_5726,N_5635,N_5621);
nand U5727 (N_5727,N_5603,N_5448);
nor U5728 (N_5728,N_5554,N_5562);
nor U5729 (N_5729,N_5602,N_5574);
nand U5730 (N_5730,N_5408,N_5680);
xnor U5731 (N_5731,N_5662,N_5481);
nand U5732 (N_5732,N_5430,N_5642);
xor U5733 (N_5733,N_5523,N_5512);
and U5734 (N_5734,N_5502,N_5496);
and U5735 (N_5735,N_5414,N_5473);
or U5736 (N_5736,N_5539,N_5524);
nand U5737 (N_5737,N_5519,N_5651);
nand U5738 (N_5738,N_5616,N_5557);
nand U5739 (N_5739,N_5507,N_5652);
xnor U5740 (N_5740,N_5427,N_5591);
and U5741 (N_5741,N_5428,N_5531);
nor U5742 (N_5742,N_5608,N_5565);
and U5743 (N_5743,N_5576,N_5613);
xnor U5744 (N_5744,N_5457,N_5696);
nand U5745 (N_5745,N_5598,N_5689);
nor U5746 (N_5746,N_5513,N_5510);
nand U5747 (N_5747,N_5607,N_5449);
xnor U5748 (N_5748,N_5679,N_5601);
nor U5749 (N_5749,N_5571,N_5547);
xor U5750 (N_5750,N_5477,N_5506);
nor U5751 (N_5751,N_5583,N_5657);
and U5752 (N_5752,N_5517,N_5442);
nor U5753 (N_5753,N_5402,N_5528);
or U5754 (N_5754,N_5491,N_5552);
or U5755 (N_5755,N_5569,N_5509);
xnor U5756 (N_5756,N_5431,N_5439);
nor U5757 (N_5757,N_5687,N_5536);
nand U5758 (N_5758,N_5677,N_5694);
and U5759 (N_5759,N_5661,N_5446);
nand U5760 (N_5760,N_5600,N_5452);
nor U5761 (N_5761,N_5643,N_5482);
nand U5762 (N_5762,N_5666,N_5584);
xnor U5763 (N_5763,N_5594,N_5614);
and U5764 (N_5764,N_5631,N_5630);
nand U5765 (N_5765,N_5566,N_5592);
nand U5766 (N_5766,N_5644,N_5675);
or U5767 (N_5767,N_5550,N_5549);
nand U5768 (N_5768,N_5535,N_5625);
nand U5769 (N_5769,N_5660,N_5440);
nand U5770 (N_5770,N_5418,N_5555);
xor U5771 (N_5771,N_5698,N_5438);
nor U5772 (N_5772,N_5508,N_5623);
or U5773 (N_5773,N_5494,N_5699);
or U5774 (N_5774,N_5470,N_5570);
xnor U5775 (N_5775,N_5604,N_5588);
xor U5776 (N_5776,N_5674,N_5465);
nand U5777 (N_5777,N_5454,N_5628);
xnor U5778 (N_5778,N_5505,N_5558);
xnor U5779 (N_5779,N_5411,N_5437);
or U5780 (N_5780,N_5475,N_5511);
or U5781 (N_5781,N_5469,N_5466);
and U5782 (N_5782,N_5518,N_5567);
and U5783 (N_5783,N_5632,N_5495);
or U5784 (N_5784,N_5492,N_5564);
nand U5785 (N_5785,N_5429,N_5615);
nand U5786 (N_5786,N_5541,N_5653);
and U5787 (N_5787,N_5587,N_5561);
nand U5788 (N_5788,N_5612,N_5530);
nor U5789 (N_5789,N_5656,N_5476);
and U5790 (N_5790,N_5640,N_5456);
nor U5791 (N_5791,N_5676,N_5667);
and U5792 (N_5792,N_5412,N_5575);
nor U5793 (N_5793,N_5420,N_5544);
nand U5794 (N_5794,N_5500,N_5415);
or U5795 (N_5795,N_5609,N_5682);
xor U5796 (N_5796,N_5596,N_5425);
or U5797 (N_5797,N_5669,N_5650);
or U5798 (N_5798,N_5527,N_5533);
xor U5799 (N_5799,N_5582,N_5480);
and U5800 (N_5800,N_5610,N_5634);
or U5801 (N_5801,N_5426,N_5489);
nor U5802 (N_5802,N_5424,N_5520);
and U5803 (N_5803,N_5441,N_5684);
or U5804 (N_5804,N_5577,N_5685);
and U5805 (N_5805,N_5435,N_5461);
and U5806 (N_5806,N_5559,N_5617);
or U5807 (N_5807,N_5406,N_5416);
and U5808 (N_5808,N_5516,N_5407);
xnor U5809 (N_5809,N_5404,N_5659);
and U5810 (N_5810,N_5537,N_5487);
xor U5811 (N_5811,N_5451,N_5645);
nand U5812 (N_5812,N_5589,N_5525);
or U5813 (N_5813,N_5581,N_5538);
nand U5814 (N_5814,N_5683,N_5629);
or U5815 (N_5815,N_5526,N_5405);
nand U5816 (N_5816,N_5401,N_5503);
nand U5817 (N_5817,N_5655,N_5499);
nor U5818 (N_5818,N_5419,N_5636);
nand U5819 (N_5819,N_5556,N_5590);
xor U5820 (N_5820,N_5658,N_5620);
nand U5821 (N_5821,N_5485,N_5553);
and U5822 (N_5822,N_5447,N_5422);
and U5823 (N_5823,N_5637,N_5462);
and U5824 (N_5824,N_5483,N_5572);
xor U5825 (N_5825,N_5436,N_5459);
xor U5826 (N_5826,N_5568,N_5622);
nor U5827 (N_5827,N_5691,N_5490);
nor U5828 (N_5828,N_5400,N_5460);
nor U5829 (N_5829,N_5649,N_5474);
xor U5830 (N_5830,N_5580,N_5693);
nand U5831 (N_5831,N_5560,N_5627);
and U5832 (N_5832,N_5573,N_5664);
nor U5833 (N_5833,N_5639,N_5514);
nor U5834 (N_5834,N_5498,N_5433);
nand U5835 (N_5835,N_5597,N_5668);
xor U5836 (N_5836,N_5618,N_5599);
and U5837 (N_5837,N_5551,N_5690);
nor U5838 (N_5838,N_5484,N_5665);
or U5839 (N_5839,N_5478,N_5697);
xnor U5840 (N_5840,N_5595,N_5626);
nor U5841 (N_5841,N_5681,N_5522);
nand U5842 (N_5842,N_5504,N_5493);
nor U5843 (N_5843,N_5624,N_5534);
and U5844 (N_5844,N_5403,N_5421);
or U5845 (N_5845,N_5546,N_5578);
and U5846 (N_5846,N_5548,N_5593);
nor U5847 (N_5847,N_5501,N_5417);
or U5848 (N_5848,N_5585,N_5468);
nor U5849 (N_5849,N_5529,N_5688);
nand U5850 (N_5850,N_5486,N_5556);
or U5851 (N_5851,N_5507,N_5519);
nor U5852 (N_5852,N_5492,N_5448);
nand U5853 (N_5853,N_5552,N_5440);
xor U5854 (N_5854,N_5622,N_5550);
or U5855 (N_5855,N_5698,N_5418);
and U5856 (N_5856,N_5482,N_5662);
and U5857 (N_5857,N_5561,N_5473);
xnor U5858 (N_5858,N_5437,N_5664);
and U5859 (N_5859,N_5419,N_5522);
nor U5860 (N_5860,N_5516,N_5424);
nor U5861 (N_5861,N_5420,N_5474);
or U5862 (N_5862,N_5613,N_5561);
nand U5863 (N_5863,N_5456,N_5543);
xnor U5864 (N_5864,N_5657,N_5630);
and U5865 (N_5865,N_5498,N_5634);
or U5866 (N_5866,N_5505,N_5660);
or U5867 (N_5867,N_5405,N_5485);
or U5868 (N_5868,N_5624,N_5519);
xor U5869 (N_5869,N_5588,N_5442);
or U5870 (N_5870,N_5494,N_5648);
and U5871 (N_5871,N_5563,N_5485);
or U5872 (N_5872,N_5503,N_5613);
xnor U5873 (N_5873,N_5645,N_5495);
or U5874 (N_5874,N_5670,N_5688);
nand U5875 (N_5875,N_5474,N_5660);
or U5876 (N_5876,N_5417,N_5422);
or U5877 (N_5877,N_5517,N_5404);
xnor U5878 (N_5878,N_5481,N_5655);
or U5879 (N_5879,N_5437,N_5504);
and U5880 (N_5880,N_5493,N_5545);
and U5881 (N_5881,N_5486,N_5471);
xor U5882 (N_5882,N_5603,N_5438);
nand U5883 (N_5883,N_5503,N_5638);
and U5884 (N_5884,N_5414,N_5590);
xor U5885 (N_5885,N_5569,N_5608);
xnor U5886 (N_5886,N_5474,N_5522);
and U5887 (N_5887,N_5489,N_5576);
or U5888 (N_5888,N_5574,N_5495);
nand U5889 (N_5889,N_5510,N_5668);
nor U5890 (N_5890,N_5461,N_5673);
nand U5891 (N_5891,N_5514,N_5670);
and U5892 (N_5892,N_5682,N_5513);
nor U5893 (N_5893,N_5564,N_5594);
and U5894 (N_5894,N_5473,N_5531);
or U5895 (N_5895,N_5627,N_5548);
xor U5896 (N_5896,N_5569,N_5498);
nand U5897 (N_5897,N_5438,N_5630);
nor U5898 (N_5898,N_5559,N_5691);
nand U5899 (N_5899,N_5401,N_5499);
xnor U5900 (N_5900,N_5437,N_5476);
nor U5901 (N_5901,N_5487,N_5528);
xor U5902 (N_5902,N_5611,N_5402);
nand U5903 (N_5903,N_5587,N_5556);
and U5904 (N_5904,N_5611,N_5573);
nor U5905 (N_5905,N_5565,N_5591);
xor U5906 (N_5906,N_5530,N_5614);
nand U5907 (N_5907,N_5481,N_5558);
xnor U5908 (N_5908,N_5438,N_5491);
and U5909 (N_5909,N_5536,N_5578);
or U5910 (N_5910,N_5581,N_5694);
or U5911 (N_5911,N_5461,N_5416);
and U5912 (N_5912,N_5578,N_5685);
nand U5913 (N_5913,N_5546,N_5504);
nor U5914 (N_5914,N_5627,N_5679);
xor U5915 (N_5915,N_5620,N_5442);
or U5916 (N_5916,N_5421,N_5517);
nand U5917 (N_5917,N_5615,N_5697);
xor U5918 (N_5918,N_5429,N_5560);
xor U5919 (N_5919,N_5614,N_5479);
or U5920 (N_5920,N_5556,N_5690);
and U5921 (N_5921,N_5454,N_5608);
xnor U5922 (N_5922,N_5435,N_5669);
nand U5923 (N_5923,N_5452,N_5619);
or U5924 (N_5924,N_5656,N_5588);
or U5925 (N_5925,N_5507,N_5624);
nor U5926 (N_5926,N_5557,N_5641);
and U5927 (N_5927,N_5435,N_5657);
and U5928 (N_5928,N_5522,N_5466);
and U5929 (N_5929,N_5647,N_5611);
xor U5930 (N_5930,N_5417,N_5418);
xor U5931 (N_5931,N_5610,N_5582);
or U5932 (N_5932,N_5639,N_5548);
nand U5933 (N_5933,N_5629,N_5543);
nand U5934 (N_5934,N_5401,N_5414);
and U5935 (N_5935,N_5606,N_5591);
and U5936 (N_5936,N_5539,N_5589);
or U5937 (N_5937,N_5656,N_5643);
nor U5938 (N_5938,N_5575,N_5521);
nand U5939 (N_5939,N_5489,N_5672);
or U5940 (N_5940,N_5593,N_5590);
nand U5941 (N_5941,N_5671,N_5697);
xnor U5942 (N_5942,N_5542,N_5539);
nand U5943 (N_5943,N_5656,N_5657);
nor U5944 (N_5944,N_5599,N_5474);
nand U5945 (N_5945,N_5402,N_5694);
nor U5946 (N_5946,N_5547,N_5634);
and U5947 (N_5947,N_5625,N_5549);
nor U5948 (N_5948,N_5401,N_5621);
xor U5949 (N_5949,N_5506,N_5516);
and U5950 (N_5950,N_5657,N_5636);
and U5951 (N_5951,N_5687,N_5491);
xnor U5952 (N_5952,N_5414,N_5488);
or U5953 (N_5953,N_5643,N_5520);
nand U5954 (N_5954,N_5476,N_5688);
xnor U5955 (N_5955,N_5650,N_5533);
nor U5956 (N_5956,N_5615,N_5519);
or U5957 (N_5957,N_5652,N_5490);
xnor U5958 (N_5958,N_5533,N_5540);
nand U5959 (N_5959,N_5550,N_5472);
nand U5960 (N_5960,N_5444,N_5572);
nor U5961 (N_5961,N_5570,N_5648);
xor U5962 (N_5962,N_5478,N_5401);
or U5963 (N_5963,N_5544,N_5542);
and U5964 (N_5964,N_5489,N_5490);
xor U5965 (N_5965,N_5458,N_5520);
xor U5966 (N_5966,N_5690,N_5692);
and U5967 (N_5967,N_5648,N_5432);
xnor U5968 (N_5968,N_5505,N_5546);
nor U5969 (N_5969,N_5519,N_5485);
nor U5970 (N_5970,N_5578,N_5623);
nand U5971 (N_5971,N_5452,N_5609);
nand U5972 (N_5972,N_5506,N_5414);
and U5973 (N_5973,N_5576,N_5694);
or U5974 (N_5974,N_5479,N_5630);
and U5975 (N_5975,N_5576,N_5662);
nor U5976 (N_5976,N_5411,N_5477);
nor U5977 (N_5977,N_5444,N_5534);
xor U5978 (N_5978,N_5675,N_5402);
xnor U5979 (N_5979,N_5650,N_5474);
and U5980 (N_5980,N_5646,N_5404);
or U5981 (N_5981,N_5602,N_5671);
nor U5982 (N_5982,N_5572,N_5656);
and U5983 (N_5983,N_5619,N_5419);
xnor U5984 (N_5984,N_5558,N_5624);
xor U5985 (N_5985,N_5551,N_5667);
nor U5986 (N_5986,N_5625,N_5512);
xor U5987 (N_5987,N_5679,N_5464);
nand U5988 (N_5988,N_5419,N_5422);
and U5989 (N_5989,N_5635,N_5657);
xor U5990 (N_5990,N_5633,N_5553);
or U5991 (N_5991,N_5456,N_5440);
and U5992 (N_5992,N_5562,N_5400);
or U5993 (N_5993,N_5497,N_5441);
nand U5994 (N_5994,N_5400,N_5454);
xor U5995 (N_5995,N_5450,N_5580);
and U5996 (N_5996,N_5684,N_5578);
nand U5997 (N_5997,N_5457,N_5569);
or U5998 (N_5998,N_5560,N_5619);
and U5999 (N_5999,N_5400,N_5561);
nand U6000 (N_6000,N_5839,N_5854);
nand U6001 (N_6001,N_5941,N_5730);
or U6002 (N_6002,N_5747,N_5804);
and U6003 (N_6003,N_5852,N_5889);
nor U6004 (N_6004,N_5760,N_5923);
nor U6005 (N_6005,N_5936,N_5811);
and U6006 (N_6006,N_5962,N_5703);
nand U6007 (N_6007,N_5818,N_5711);
xnor U6008 (N_6008,N_5914,N_5769);
and U6009 (N_6009,N_5900,N_5890);
nor U6010 (N_6010,N_5754,N_5779);
or U6011 (N_6011,N_5857,N_5996);
or U6012 (N_6012,N_5847,N_5888);
or U6013 (N_6013,N_5970,N_5834);
and U6014 (N_6014,N_5731,N_5904);
nor U6015 (N_6015,N_5708,N_5757);
nand U6016 (N_6016,N_5773,N_5901);
nand U6017 (N_6017,N_5792,N_5809);
nand U6018 (N_6018,N_5785,N_5894);
xnor U6019 (N_6019,N_5994,N_5802);
nor U6020 (N_6020,N_5915,N_5828);
nor U6021 (N_6021,N_5976,N_5748);
xnor U6022 (N_6022,N_5930,N_5728);
nand U6023 (N_6023,N_5943,N_5856);
xnor U6024 (N_6024,N_5766,N_5750);
nor U6025 (N_6025,N_5843,N_5998);
and U6026 (N_6026,N_5793,N_5895);
nand U6027 (N_6027,N_5937,N_5922);
and U6028 (N_6028,N_5831,N_5739);
and U6029 (N_6029,N_5830,N_5737);
nand U6030 (N_6030,N_5898,N_5704);
xor U6031 (N_6031,N_5720,N_5876);
or U6032 (N_6032,N_5745,N_5826);
nand U6033 (N_6033,N_5764,N_5710);
xnor U6034 (N_6034,N_5806,N_5963);
nand U6035 (N_6035,N_5893,N_5749);
nand U6036 (N_6036,N_5794,N_5928);
or U6037 (N_6037,N_5991,N_5925);
nor U6038 (N_6038,N_5807,N_5988);
and U6039 (N_6039,N_5722,N_5741);
xor U6040 (N_6040,N_5944,N_5872);
and U6041 (N_6041,N_5887,N_5907);
nor U6042 (N_6042,N_5786,N_5924);
xor U6043 (N_6043,N_5926,N_5761);
nand U6044 (N_6044,N_5956,N_5995);
and U6045 (N_6045,N_5961,N_5712);
or U6046 (N_6046,N_5756,N_5951);
nor U6047 (N_6047,N_5734,N_5906);
nand U6048 (N_6048,N_5784,N_5952);
and U6049 (N_6049,N_5871,N_5860);
nor U6050 (N_6050,N_5935,N_5875);
and U6051 (N_6051,N_5724,N_5873);
nor U6052 (N_6052,N_5844,N_5767);
or U6053 (N_6053,N_5974,N_5788);
xor U6054 (N_6054,N_5886,N_5732);
xor U6055 (N_6055,N_5990,N_5978);
nor U6056 (N_6056,N_5816,N_5735);
nand U6057 (N_6057,N_5848,N_5950);
nor U6058 (N_6058,N_5927,N_5966);
xor U6059 (N_6059,N_5981,N_5780);
xnor U6060 (N_6060,N_5837,N_5993);
and U6061 (N_6061,N_5940,N_5999);
xnor U6062 (N_6062,N_5973,N_5789);
xor U6063 (N_6063,N_5706,N_5771);
xor U6064 (N_6064,N_5835,N_5972);
xor U6065 (N_6065,N_5954,N_5822);
or U6066 (N_6066,N_5958,N_5759);
nand U6067 (N_6067,N_5984,N_5909);
or U6068 (N_6068,N_5808,N_5862);
xor U6069 (N_6069,N_5989,N_5714);
nand U6070 (N_6070,N_5934,N_5740);
and U6071 (N_6071,N_5982,N_5823);
nor U6072 (N_6072,N_5920,N_5883);
and U6073 (N_6073,N_5846,N_5881);
and U6074 (N_6074,N_5772,N_5736);
nor U6075 (N_6075,N_5700,N_5803);
or U6076 (N_6076,N_5945,N_5863);
and U6077 (N_6077,N_5905,N_5902);
nand U6078 (N_6078,N_5752,N_5916);
nand U6079 (N_6079,N_5838,N_5791);
nor U6080 (N_6080,N_5949,N_5777);
nand U6081 (N_6081,N_5824,N_5762);
xor U6082 (N_6082,N_5866,N_5765);
nand U6083 (N_6083,N_5948,N_5727);
nand U6084 (N_6084,N_5778,N_5874);
nor U6085 (N_6085,N_5709,N_5983);
or U6086 (N_6086,N_5836,N_5965);
nor U6087 (N_6087,N_5885,N_5865);
and U6088 (N_6088,N_5742,N_5774);
and U6089 (N_6089,N_5849,N_5878);
or U6090 (N_6090,N_5845,N_5917);
nand U6091 (N_6091,N_5933,N_5971);
and U6092 (N_6092,N_5987,N_5858);
and U6093 (N_6093,N_5701,N_5851);
and U6094 (N_6094,N_5841,N_5781);
or U6095 (N_6095,N_5850,N_5790);
nor U6096 (N_6096,N_5912,N_5719);
and U6097 (N_6097,N_5763,N_5755);
nand U6098 (N_6098,N_5861,N_5795);
nor U6099 (N_6099,N_5725,N_5896);
xnor U6100 (N_6100,N_5827,N_5832);
xor U6101 (N_6101,N_5744,N_5979);
or U6102 (N_6102,N_5913,N_5814);
or U6103 (N_6103,N_5817,N_5867);
xnor U6104 (N_6104,N_5969,N_5942);
xor U6105 (N_6105,N_5733,N_5776);
and U6106 (N_6106,N_5967,N_5903);
and U6107 (N_6107,N_5947,N_5738);
or U6108 (N_6108,N_5820,N_5798);
nor U6109 (N_6109,N_5980,N_5829);
and U6110 (N_6110,N_5855,N_5997);
xor U6111 (N_6111,N_5892,N_5721);
nand U6112 (N_6112,N_5953,N_5833);
nand U6113 (N_6113,N_5812,N_5985);
xnor U6114 (N_6114,N_5910,N_5718);
or U6115 (N_6115,N_5751,N_5702);
and U6116 (N_6116,N_5783,N_5717);
and U6117 (N_6117,N_5840,N_5932);
xor U6118 (N_6118,N_5770,N_5929);
xor U6119 (N_6119,N_5815,N_5782);
nand U6120 (N_6120,N_5879,N_5884);
nor U6121 (N_6121,N_5964,N_5758);
and U6122 (N_6122,N_5869,N_5918);
xor U6123 (N_6123,N_5768,N_5715);
or U6124 (N_6124,N_5799,N_5746);
nand U6125 (N_6125,N_5716,N_5796);
or U6126 (N_6126,N_5797,N_5713);
nand U6127 (N_6127,N_5805,N_5931);
nand U6128 (N_6128,N_5938,N_5897);
nor U6129 (N_6129,N_5864,N_5743);
and U6130 (N_6130,N_5821,N_5959);
nor U6131 (N_6131,N_5975,N_5877);
nand U6132 (N_6132,N_5868,N_5753);
nor U6133 (N_6133,N_5729,N_5992);
nor U6134 (N_6134,N_5957,N_5853);
or U6135 (N_6135,N_5810,N_5946);
nand U6136 (N_6136,N_5968,N_5919);
xnor U6137 (N_6137,N_5921,N_5800);
nor U6138 (N_6138,N_5859,N_5819);
or U6139 (N_6139,N_5880,N_5726);
and U6140 (N_6140,N_5882,N_5825);
nor U6141 (N_6141,N_5775,N_5787);
nor U6142 (N_6142,N_5955,N_5899);
nand U6143 (N_6143,N_5960,N_5939);
nor U6144 (N_6144,N_5801,N_5908);
nor U6145 (N_6145,N_5870,N_5707);
nor U6146 (N_6146,N_5911,N_5891);
nor U6147 (N_6147,N_5705,N_5813);
or U6148 (N_6148,N_5842,N_5977);
or U6149 (N_6149,N_5986,N_5723);
nor U6150 (N_6150,N_5922,N_5796);
or U6151 (N_6151,N_5974,N_5766);
nor U6152 (N_6152,N_5987,N_5938);
nor U6153 (N_6153,N_5945,N_5806);
or U6154 (N_6154,N_5736,N_5850);
or U6155 (N_6155,N_5749,N_5836);
xnor U6156 (N_6156,N_5758,N_5724);
nor U6157 (N_6157,N_5866,N_5702);
and U6158 (N_6158,N_5884,N_5700);
nand U6159 (N_6159,N_5803,N_5732);
nor U6160 (N_6160,N_5822,N_5963);
xnor U6161 (N_6161,N_5919,N_5996);
xnor U6162 (N_6162,N_5919,N_5767);
nand U6163 (N_6163,N_5842,N_5847);
nor U6164 (N_6164,N_5832,N_5719);
xor U6165 (N_6165,N_5775,N_5896);
xnor U6166 (N_6166,N_5714,N_5946);
and U6167 (N_6167,N_5761,N_5710);
nor U6168 (N_6168,N_5860,N_5973);
xnor U6169 (N_6169,N_5905,N_5922);
and U6170 (N_6170,N_5801,N_5798);
nand U6171 (N_6171,N_5974,N_5765);
nor U6172 (N_6172,N_5878,N_5943);
and U6173 (N_6173,N_5744,N_5859);
nor U6174 (N_6174,N_5850,N_5928);
and U6175 (N_6175,N_5743,N_5710);
nand U6176 (N_6176,N_5973,N_5728);
and U6177 (N_6177,N_5815,N_5941);
and U6178 (N_6178,N_5887,N_5800);
xor U6179 (N_6179,N_5957,N_5723);
and U6180 (N_6180,N_5948,N_5960);
nand U6181 (N_6181,N_5765,N_5785);
xor U6182 (N_6182,N_5737,N_5798);
or U6183 (N_6183,N_5914,N_5852);
xor U6184 (N_6184,N_5773,N_5725);
xnor U6185 (N_6185,N_5779,N_5930);
nand U6186 (N_6186,N_5790,N_5974);
xor U6187 (N_6187,N_5822,N_5735);
or U6188 (N_6188,N_5987,N_5877);
and U6189 (N_6189,N_5941,N_5932);
and U6190 (N_6190,N_5873,N_5841);
and U6191 (N_6191,N_5739,N_5925);
nor U6192 (N_6192,N_5724,N_5948);
and U6193 (N_6193,N_5946,N_5792);
nor U6194 (N_6194,N_5833,N_5860);
and U6195 (N_6195,N_5750,N_5789);
or U6196 (N_6196,N_5959,N_5745);
or U6197 (N_6197,N_5976,N_5900);
nor U6198 (N_6198,N_5839,N_5972);
nor U6199 (N_6199,N_5930,N_5890);
and U6200 (N_6200,N_5856,N_5719);
nor U6201 (N_6201,N_5973,N_5755);
nand U6202 (N_6202,N_5845,N_5873);
nor U6203 (N_6203,N_5991,N_5989);
and U6204 (N_6204,N_5787,N_5926);
and U6205 (N_6205,N_5745,N_5836);
xor U6206 (N_6206,N_5916,N_5839);
nor U6207 (N_6207,N_5889,N_5880);
xnor U6208 (N_6208,N_5959,N_5889);
nor U6209 (N_6209,N_5937,N_5854);
and U6210 (N_6210,N_5970,N_5725);
nor U6211 (N_6211,N_5910,N_5948);
nor U6212 (N_6212,N_5915,N_5733);
or U6213 (N_6213,N_5739,N_5761);
and U6214 (N_6214,N_5990,N_5712);
or U6215 (N_6215,N_5922,N_5885);
or U6216 (N_6216,N_5739,N_5836);
nand U6217 (N_6217,N_5725,N_5737);
or U6218 (N_6218,N_5706,N_5893);
nor U6219 (N_6219,N_5875,N_5907);
nor U6220 (N_6220,N_5831,N_5860);
nand U6221 (N_6221,N_5748,N_5866);
nand U6222 (N_6222,N_5704,N_5890);
nor U6223 (N_6223,N_5775,N_5800);
and U6224 (N_6224,N_5987,N_5765);
or U6225 (N_6225,N_5875,N_5937);
nand U6226 (N_6226,N_5955,N_5898);
or U6227 (N_6227,N_5960,N_5840);
nand U6228 (N_6228,N_5918,N_5866);
nor U6229 (N_6229,N_5915,N_5811);
and U6230 (N_6230,N_5930,N_5804);
xor U6231 (N_6231,N_5857,N_5910);
and U6232 (N_6232,N_5985,N_5913);
xor U6233 (N_6233,N_5871,N_5768);
and U6234 (N_6234,N_5880,N_5882);
or U6235 (N_6235,N_5703,N_5933);
or U6236 (N_6236,N_5830,N_5859);
xor U6237 (N_6237,N_5937,N_5843);
and U6238 (N_6238,N_5941,N_5945);
xor U6239 (N_6239,N_5754,N_5873);
nand U6240 (N_6240,N_5898,N_5730);
xnor U6241 (N_6241,N_5817,N_5949);
or U6242 (N_6242,N_5816,N_5869);
or U6243 (N_6243,N_5995,N_5990);
or U6244 (N_6244,N_5752,N_5734);
xnor U6245 (N_6245,N_5773,N_5958);
nor U6246 (N_6246,N_5845,N_5880);
or U6247 (N_6247,N_5818,N_5755);
nor U6248 (N_6248,N_5822,N_5845);
xor U6249 (N_6249,N_5921,N_5843);
and U6250 (N_6250,N_5728,N_5786);
nor U6251 (N_6251,N_5945,N_5943);
xnor U6252 (N_6252,N_5718,N_5781);
xnor U6253 (N_6253,N_5842,N_5907);
xnor U6254 (N_6254,N_5818,N_5826);
and U6255 (N_6255,N_5798,N_5812);
nor U6256 (N_6256,N_5879,N_5740);
or U6257 (N_6257,N_5945,N_5942);
nor U6258 (N_6258,N_5932,N_5894);
or U6259 (N_6259,N_5981,N_5843);
nor U6260 (N_6260,N_5987,N_5907);
nor U6261 (N_6261,N_5974,N_5750);
nor U6262 (N_6262,N_5985,N_5924);
xnor U6263 (N_6263,N_5970,N_5942);
nor U6264 (N_6264,N_5782,N_5911);
nor U6265 (N_6265,N_5992,N_5943);
or U6266 (N_6266,N_5983,N_5896);
xor U6267 (N_6267,N_5831,N_5853);
nand U6268 (N_6268,N_5804,N_5711);
xnor U6269 (N_6269,N_5968,N_5924);
xnor U6270 (N_6270,N_5970,N_5747);
xnor U6271 (N_6271,N_5933,N_5977);
and U6272 (N_6272,N_5860,N_5845);
or U6273 (N_6273,N_5917,N_5851);
nand U6274 (N_6274,N_5726,N_5915);
or U6275 (N_6275,N_5938,N_5811);
xor U6276 (N_6276,N_5966,N_5834);
xor U6277 (N_6277,N_5868,N_5726);
or U6278 (N_6278,N_5895,N_5975);
xor U6279 (N_6279,N_5818,N_5861);
xor U6280 (N_6280,N_5751,N_5827);
and U6281 (N_6281,N_5889,N_5731);
xor U6282 (N_6282,N_5856,N_5879);
nor U6283 (N_6283,N_5910,N_5993);
xor U6284 (N_6284,N_5898,N_5885);
nand U6285 (N_6285,N_5817,N_5760);
or U6286 (N_6286,N_5779,N_5977);
xor U6287 (N_6287,N_5802,N_5914);
and U6288 (N_6288,N_5810,N_5970);
or U6289 (N_6289,N_5975,N_5885);
xnor U6290 (N_6290,N_5763,N_5970);
nand U6291 (N_6291,N_5753,N_5995);
xnor U6292 (N_6292,N_5779,N_5967);
xnor U6293 (N_6293,N_5827,N_5779);
nor U6294 (N_6294,N_5833,N_5938);
nor U6295 (N_6295,N_5796,N_5831);
xor U6296 (N_6296,N_5892,N_5982);
nor U6297 (N_6297,N_5986,N_5854);
and U6298 (N_6298,N_5851,N_5813);
or U6299 (N_6299,N_5973,N_5766);
and U6300 (N_6300,N_6068,N_6001);
nor U6301 (N_6301,N_6047,N_6230);
and U6302 (N_6302,N_6182,N_6150);
xnor U6303 (N_6303,N_6238,N_6133);
nand U6304 (N_6304,N_6161,N_6052);
xor U6305 (N_6305,N_6167,N_6169);
nor U6306 (N_6306,N_6264,N_6080);
xnor U6307 (N_6307,N_6060,N_6130);
xnor U6308 (N_6308,N_6078,N_6241);
nor U6309 (N_6309,N_6132,N_6252);
xnor U6310 (N_6310,N_6156,N_6114);
and U6311 (N_6311,N_6208,N_6269);
xor U6312 (N_6312,N_6012,N_6065);
xor U6313 (N_6313,N_6261,N_6263);
nor U6314 (N_6314,N_6103,N_6192);
xnor U6315 (N_6315,N_6274,N_6246);
xor U6316 (N_6316,N_6070,N_6044);
xnor U6317 (N_6317,N_6179,N_6104);
or U6318 (N_6318,N_6101,N_6049);
nor U6319 (N_6319,N_6096,N_6011);
xor U6320 (N_6320,N_6088,N_6066);
or U6321 (N_6321,N_6211,N_6021);
nor U6322 (N_6322,N_6216,N_6102);
or U6323 (N_6323,N_6034,N_6260);
and U6324 (N_6324,N_6199,N_6018);
xnor U6325 (N_6325,N_6178,N_6267);
and U6326 (N_6326,N_6069,N_6147);
nand U6327 (N_6327,N_6220,N_6146);
xnor U6328 (N_6328,N_6235,N_6038);
nor U6329 (N_6329,N_6223,N_6091);
and U6330 (N_6330,N_6154,N_6090);
nor U6331 (N_6331,N_6053,N_6042);
or U6332 (N_6332,N_6284,N_6159);
nand U6333 (N_6333,N_6128,N_6055);
xnor U6334 (N_6334,N_6099,N_6119);
nand U6335 (N_6335,N_6287,N_6174);
nand U6336 (N_6336,N_6243,N_6033);
nand U6337 (N_6337,N_6163,N_6266);
and U6338 (N_6338,N_6073,N_6109);
nor U6339 (N_6339,N_6257,N_6024);
xor U6340 (N_6340,N_6196,N_6268);
or U6341 (N_6341,N_6084,N_6108);
nand U6342 (N_6342,N_6014,N_6278);
nor U6343 (N_6343,N_6265,N_6105);
xnor U6344 (N_6344,N_6253,N_6095);
xnor U6345 (N_6345,N_6189,N_6110);
xnor U6346 (N_6346,N_6219,N_6258);
or U6347 (N_6347,N_6239,N_6272);
xnor U6348 (N_6348,N_6005,N_6125);
nor U6349 (N_6349,N_6247,N_6037);
nor U6350 (N_6350,N_6059,N_6111);
nand U6351 (N_6351,N_6008,N_6112);
and U6352 (N_6352,N_6067,N_6072);
or U6353 (N_6353,N_6200,N_6181);
nor U6354 (N_6354,N_6164,N_6116);
nand U6355 (N_6355,N_6143,N_6175);
nand U6356 (N_6356,N_6135,N_6121);
and U6357 (N_6357,N_6085,N_6298);
xor U6358 (N_6358,N_6195,N_6213);
nor U6359 (N_6359,N_6045,N_6023);
nor U6360 (N_6360,N_6129,N_6282);
or U6361 (N_6361,N_6134,N_6187);
nor U6362 (N_6362,N_6122,N_6126);
xor U6363 (N_6363,N_6145,N_6288);
or U6364 (N_6364,N_6294,N_6207);
xor U6365 (N_6365,N_6276,N_6249);
nor U6366 (N_6366,N_6149,N_6283);
nand U6367 (N_6367,N_6290,N_6003);
and U6368 (N_6368,N_6035,N_6215);
and U6369 (N_6369,N_6074,N_6032);
or U6370 (N_6370,N_6291,N_6270);
nand U6371 (N_6371,N_6089,N_6227);
or U6372 (N_6372,N_6240,N_6214);
nor U6373 (N_6373,N_6019,N_6170);
nand U6374 (N_6374,N_6212,N_6117);
nor U6375 (N_6375,N_6141,N_6275);
xor U6376 (N_6376,N_6234,N_6098);
or U6377 (N_6377,N_6262,N_6115);
xnor U6378 (N_6378,N_6177,N_6118);
nand U6379 (N_6379,N_6009,N_6222);
xor U6380 (N_6380,N_6006,N_6079);
nand U6381 (N_6381,N_6093,N_6013);
and U6382 (N_6382,N_6016,N_6131);
nand U6383 (N_6383,N_6158,N_6277);
nand U6384 (N_6384,N_6190,N_6194);
nand U6385 (N_6385,N_6236,N_6046);
nand U6386 (N_6386,N_6092,N_6279);
and U6387 (N_6387,N_6124,N_6025);
nor U6388 (N_6388,N_6086,N_6048);
nand U6389 (N_6389,N_6289,N_6157);
nor U6390 (N_6390,N_6259,N_6028);
xor U6391 (N_6391,N_6136,N_6206);
xor U6392 (N_6392,N_6137,N_6286);
nor U6393 (N_6393,N_6029,N_6063);
nand U6394 (N_6394,N_6077,N_6030);
nor U6395 (N_6395,N_6043,N_6185);
or U6396 (N_6396,N_6142,N_6296);
and U6397 (N_6397,N_6062,N_6094);
xor U6398 (N_6398,N_6224,N_6297);
xor U6399 (N_6399,N_6271,N_6209);
and U6400 (N_6400,N_6002,N_6000);
xnor U6401 (N_6401,N_6040,N_6076);
nor U6402 (N_6402,N_6285,N_6039);
nand U6403 (N_6403,N_6244,N_6015);
and U6404 (N_6404,N_6054,N_6248);
xnor U6405 (N_6405,N_6255,N_6056);
nor U6406 (N_6406,N_6250,N_6233);
and U6407 (N_6407,N_6191,N_6186);
and U6408 (N_6408,N_6188,N_6251);
nand U6409 (N_6409,N_6237,N_6201);
and U6410 (N_6410,N_6113,N_6075);
or U6411 (N_6411,N_6081,N_6058);
nor U6412 (N_6412,N_6082,N_6010);
and U6413 (N_6413,N_6097,N_6281);
and U6414 (N_6414,N_6183,N_6100);
nor U6415 (N_6415,N_6245,N_6151);
or U6416 (N_6416,N_6184,N_6221);
or U6417 (N_6417,N_6232,N_6026);
and U6418 (N_6418,N_6280,N_6210);
nor U6419 (N_6419,N_6138,N_6180);
and U6420 (N_6420,N_6036,N_6299);
nor U6421 (N_6421,N_6051,N_6166);
and U6422 (N_6422,N_6050,N_6273);
or U6423 (N_6423,N_6017,N_6172);
or U6424 (N_6424,N_6160,N_6231);
xor U6425 (N_6425,N_6020,N_6165);
nand U6426 (N_6426,N_6173,N_6155);
nor U6427 (N_6427,N_6152,N_6004);
nor U6428 (N_6428,N_6197,N_6107);
xor U6429 (N_6429,N_6242,N_6123);
or U6430 (N_6430,N_6202,N_6162);
nand U6431 (N_6431,N_6140,N_6027);
and U6432 (N_6432,N_6171,N_6087);
nor U6433 (N_6433,N_6106,N_6127);
or U6434 (N_6434,N_6057,N_6064);
xnor U6435 (N_6435,N_6031,N_6041);
nand U6436 (N_6436,N_6193,N_6198);
nand U6437 (N_6437,N_6007,N_6254);
and U6438 (N_6438,N_6293,N_6144);
and U6439 (N_6439,N_6204,N_6225);
or U6440 (N_6440,N_6083,N_6022);
nor U6441 (N_6441,N_6139,N_6176);
xor U6442 (N_6442,N_6203,N_6217);
and U6443 (N_6443,N_6295,N_6120);
and U6444 (N_6444,N_6168,N_6229);
nand U6445 (N_6445,N_6228,N_6061);
nor U6446 (N_6446,N_6226,N_6205);
nor U6447 (N_6447,N_6292,N_6148);
nand U6448 (N_6448,N_6153,N_6218);
or U6449 (N_6449,N_6256,N_6071);
xnor U6450 (N_6450,N_6293,N_6018);
nor U6451 (N_6451,N_6157,N_6171);
nand U6452 (N_6452,N_6194,N_6286);
nor U6453 (N_6453,N_6167,N_6102);
and U6454 (N_6454,N_6280,N_6269);
xor U6455 (N_6455,N_6005,N_6019);
nor U6456 (N_6456,N_6030,N_6138);
and U6457 (N_6457,N_6238,N_6248);
xnor U6458 (N_6458,N_6232,N_6262);
and U6459 (N_6459,N_6202,N_6046);
xnor U6460 (N_6460,N_6029,N_6009);
xor U6461 (N_6461,N_6243,N_6262);
or U6462 (N_6462,N_6034,N_6184);
and U6463 (N_6463,N_6249,N_6104);
nand U6464 (N_6464,N_6167,N_6164);
or U6465 (N_6465,N_6064,N_6293);
nor U6466 (N_6466,N_6262,N_6216);
xnor U6467 (N_6467,N_6110,N_6009);
xor U6468 (N_6468,N_6110,N_6054);
or U6469 (N_6469,N_6103,N_6158);
and U6470 (N_6470,N_6272,N_6237);
and U6471 (N_6471,N_6047,N_6069);
and U6472 (N_6472,N_6034,N_6047);
xor U6473 (N_6473,N_6259,N_6208);
nand U6474 (N_6474,N_6161,N_6095);
nand U6475 (N_6475,N_6179,N_6008);
xor U6476 (N_6476,N_6221,N_6249);
or U6477 (N_6477,N_6015,N_6112);
nand U6478 (N_6478,N_6021,N_6030);
nor U6479 (N_6479,N_6002,N_6043);
and U6480 (N_6480,N_6266,N_6178);
xnor U6481 (N_6481,N_6063,N_6132);
xor U6482 (N_6482,N_6053,N_6037);
or U6483 (N_6483,N_6275,N_6085);
or U6484 (N_6484,N_6134,N_6043);
and U6485 (N_6485,N_6265,N_6039);
nor U6486 (N_6486,N_6033,N_6020);
nor U6487 (N_6487,N_6260,N_6157);
xnor U6488 (N_6488,N_6154,N_6061);
or U6489 (N_6489,N_6254,N_6237);
and U6490 (N_6490,N_6201,N_6135);
and U6491 (N_6491,N_6021,N_6172);
nand U6492 (N_6492,N_6220,N_6021);
and U6493 (N_6493,N_6177,N_6126);
and U6494 (N_6494,N_6184,N_6278);
nand U6495 (N_6495,N_6000,N_6052);
nor U6496 (N_6496,N_6279,N_6077);
or U6497 (N_6497,N_6177,N_6014);
nor U6498 (N_6498,N_6257,N_6099);
nor U6499 (N_6499,N_6207,N_6165);
and U6500 (N_6500,N_6202,N_6052);
nand U6501 (N_6501,N_6100,N_6281);
xor U6502 (N_6502,N_6020,N_6139);
and U6503 (N_6503,N_6275,N_6066);
xnor U6504 (N_6504,N_6143,N_6103);
xnor U6505 (N_6505,N_6044,N_6243);
xor U6506 (N_6506,N_6056,N_6012);
and U6507 (N_6507,N_6088,N_6160);
or U6508 (N_6508,N_6196,N_6221);
nor U6509 (N_6509,N_6272,N_6248);
nor U6510 (N_6510,N_6277,N_6236);
or U6511 (N_6511,N_6016,N_6173);
nand U6512 (N_6512,N_6110,N_6039);
or U6513 (N_6513,N_6141,N_6017);
or U6514 (N_6514,N_6158,N_6180);
and U6515 (N_6515,N_6168,N_6100);
nor U6516 (N_6516,N_6016,N_6278);
or U6517 (N_6517,N_6122,N_6187);
or U6518 (N_6518,N_6205,N_6179);
and U6519 (N_6519,N_6012,N_6109);
xor U6520 (N_6520,N_6134,N_6051);
or U6521 (N_6521,N_6063,N_6119);
and U6522 (N_6522,N_6030,N_6057);
xnor U6523 (N_6523,N_6123,N_6003);
nor U6524 (N_6524,N_6051,N_6121);
and U6525 (N_6525,N_6145,N_6270);
or U6526 (N_6526,N_6211,N_6285);
and U6527 (N_6527,N_6022,N_6246);
and U6528 (N_6528,N_6239,N_6184);
and U6529 (N_6529,N_6126,N_6118);
nand U6530 (N_6530,N_6170,N_6149);
nor U6531 (N_6531,N_6177,N_6275);
nand U6532 (N_6532,N_6252,N_6091);
and U6533 (N_6533,N_6103,N_6048);
nand U6534 (N_6534,N_6114,N_6120);
xor U6535 (N_6535,N_6082,N_6001);
nand U6536 (N_6536,N_6259,N_6162);
xor U6537 (N_6537,N_6084,N_6271);
and U6538 (N_6538,N_6077,N_6053);
or U6539 (N_6539,N_6226,N_6225);
and U6540 (N_6540,N_6269,N_6249);
nor U6541 (N_6541,N_6117,N_6222);
nand U6542 (N_6542,N_6031,N_6106);
xor U6543 (N_6543,N_6227,N_6255);
xnor U6544 (N_6544,N_6219,N_6205);
or U6545 (N_6545,N_6238,N_6260);
nand U6546 (N_6546,N_6223,N_6296);
and U6547 (N_6547,N_6134,N_6084);
xnor U6548 (N_6548,N_6234,N_6275);
and U6549 (N_6549,N_6205,N_6099);
or U6550 (N_6550,N_6275,N_6133);
or U6551 (N_6551,N_6145,N_6250);
xnor U6552 (N_6552,N_6191,N_6197);
and U6553 (N_6553,N_6011,N_6215);
nand U6554 (N_6554,N_6017,N_6067);
and U6555 (N_6555,N_6299,N_6064);
nor U6556 (N_6556,N_6105,N_6054);
nor U6557 (N_6557,N_6050,N_6101);
or U6558 (N_6558,N_6248,N_6296);
xnor U6559 (N_6559,N_6096,N_6211);
xor U6560 (N_6560,N_6010,N_6139);
xnor U6561 (N_6561,N_6187,N_6251);
nor U6562 (N_6562,N_6238,N_6070);
or U6563 (N_6563,N_6067,N_6080);
xnor U6564 (N_6564,N_6223,N_6073);
nor U6565 (N_6565,N_6252,N_6181);
and U6566 (N_6566,N_6048,N_6139);
and U6567 (N_6567,N_6006,N_6018);
and U6568 (N_6568,N_6065,N_6155);
nand U6569 (N_6569,N_6116,N_6260);
or U6570 (N_6570,N_6131,N_6132);
and U6571 (N_6571,N_6006,N_6293);
or U6572 (N_6572,N_6060,N_6166);
or U6573 (N_6573,N_6105,N_6191);
nand U6574 (N_6574,N_6167,N_6220);
or U6575 (N_6575,N_6235,N_6229);
nand U6576 (N_6576,N_6156,N_6263);
nor U6577 (N_6577,N_6198,N_6091);
or U6578 (N_6578,N_6273,N_6119);
nand U6579 (N_6579,N_6237,N_6097);
xnor U6580 (N_6580,N_6161,N_6045);
and U6581 (N_6581,N_6277,N_6246);
nand U6582 (N_6582,N_6249,N_6089);
or U6583 (N_6583,N_6184,N_6010);
nand U6584 (N_6584,N_6039,N_6060);
nand U6585 (N_6585,N_6036,N_6194);
nor U6586 (N_6586,N_6153,N_6237);
and U6587 (N_6587,N_6235,N_6158);
and U6588 (N_6588,N_6047,N_6236);
nand U6589 (N_6589,N_6109,N_6182);
nor U6590 (N_6590,N_6116,N_6020);
nand U6591 (N_6591,N_6277,N_6212);
xnor U6592 (N_6592,N_6161,N_6186);
nor U6593 (N_6593,N_6168,N_6010);
nor U6594 (N_6594,N_6037,N_6127);
nand U6595 (N_6595,N_6025,N_6276);
or U6596 (N_6596,N_6212,N_6091);
nand U6597 (N_6597,N_6137,N_6074);
xor U6598 (N_6598,N_6116,N_6288);
nand U6599 (N_6599,N_6020,N_6140);
nor U6600 (N_6600,N_6347,N_6489);
and U6601 (N_6601,N_6394,N_6430);
nand U6602 (N_6602,N_6551,N_6423);
and U6603 (N_6603,N_6594,N_6416);
xor U6604 (N_6604,N_6498,N_6371);
and U6605 (N_6605,N_6348,N_6384);
nand U6606 (N_6606,N_6346,N_6548);
or U6607 (N_6607,N_6533,N_6504);
nor U6608 (N_6608,N_6494,N_6380);
nor U6609 (N_6609,N_6309,N_6539);
xor U6610 (N_6610,N_6321,N_6354);
xor U6611 (N_6611,N_6334,N_6442);
nor U6612 (N_6612,N_6395,N_6529);
xnor U6613 (N_6613,N_6344,N_6385);
or U6614 (N_6614,N_6358,N_6351);
nor U6615 (N_6615,N_6373,N_6443);
nor U6616 (N_6616,N_6537,N_6499);
nand U6617 (N_6617,N_6428,N_6595);
xor U6618 (N_6618,N_6462,N_6433);
and U6619 (N_6619,N_6304,N_6524);
or U6620 (N_6620,N_6417,N_6463);
nand U6621 (N_6621,N_6389,N_6363);
or U6622 (N_6622,N_6573,N_6425);
nor U6623 (N_6623,N_6515,N_6514);
and U6624 (N_6624,N_6592,N_6406);
or U6625 (N_6625,N_6584,N_6306);
and U6626 (N_6626,N_6598,N_6362);
or U6627 (N_6627,N_6545,N_6314);
xor U6628 (N_6628,N_6471,N_6340);
and U6629 (N_6629,N_6476,N_6331);
nand U6630 (N_6630,N_6536,N_6410);
nand U6631 (N_6631,N_6557,N_6313);
nand U6632 (N_6632,N_6318,N_6368);
nor U6633 (N_6633,N_6572,N_6550);
xnor U6634 (N_6634,N_6307,N_6597);
nor U6635 (N_6635,N_6458,N_6356);
xor U6636 (N_6636,N_6448,N_6342);
nand U6637 (N_6637,N_6452,N_6538);
xor U6638 (N_6638,N_6563,N_6386);
or U6639 (N_6639,N_6427,N_6420);
nor U6640 (N_6640,N_6470,N_6568);
or U6641 (N_6641,N_6405,N_6581);
or U6642 (N_6642,N_6345,N_6571);
nor U6643 (N_6643,N_6378,N_6349);
or U6644 (N_6644,N_6479,N_6311);
and U6645 (N_6645,N_6408,N_6370);
nor U6646 (N_6646,N_6361,N_6507);
nand U6647 (N_6647,N_6399,N_6352);
nand U6648 (N_6648,N_6468,N_6559);
xnor U6649 (N_6649,N_6560,N_6464);
and U6650 (N_6650,N_6517,N_6583);
and U6651 (N_6651,N_6453,N_6534);
or U6652 (N_6652,N_6511,N_6455);
nand U6653 (N_6653,N_6407,N_6400);
xor U6654 (N_6654,N_6409,N_6403);
nand U6655 (N_6655,N_6465,N_6301);
nor U6656 (N_6656,N_6308,N_6404);
xor U6657 (N_6657,N_6555,N_6552);
xnor U6658 (N_6658,N_6535,N_6580);
xor U6659 (N_6659,N_6429,N_6335);
and U6660 (N_6660,N_6381,N_6305);
xnor U6661 (N_6661,N_6501,N_6554);
and U6662 (N_6662,N_6549,N_6502);
xnor U6663 (N_6663,N_6543,N_6508);
xor U6664 (N_6664,N_6558,N_6325);
or U6665 (N_6665,N_6466,N_6522);
nand U6666 (N_6666,N_6577,N_6412);
xnor U6667 (N_6667,N_6493,N_6328);
nand U6668 (N_6668,N_6461,N_6451);
nor U6669 (N_6669,N_6477,N_6319);
xor U6670 (N_6670,N_6357,N_6388);
xor U6671 (N_6671,N_6491,N_6323);
and U6672 (N_6672,N_6431,N_6565);
nor U6673 (N_6673,N_6485,N_6413);
or U6674 (N_6674,N_6480,N_6329);
nor U6675 (N_6675,N_6570,N_6590);
xnor U6676 (N_6676,N_6435,N_6509);
nor U6677 (N_6677,N_6444,N_6588);
nand U6678 (N_6678,N_6398,N_6397);
nand U6679 (N_6679,N_6383,N_6422);
nor U6680 (N_6680,N_6366,N_6591);
or U6681 (N_6681,N_6582,N_6574);
and U6682 (N_6682,N_6364,N_6376);
xor U6683 (N_6683,N_6488,N_6542);
xnor U6684 (N_6684,N_6482,N_6439);
or U6685 (N_6685,N_6421,N_6379);
nand U6686 (N_6686,N_6490,N_6327);
nor U6687 (N_6687,N_6332,N_6569);
or U6688 (N_6688,N_6437,N_6372);
nor U6689 (N_6689,N_6396,N_6374);
and U6690 (N_6690,N_6415,N_6547);
nand U6691 (N_6691,N_6492,N_6546);
xnor U6692 (N_6692,N_6316,N_6481);
or U6693 (N_6693,N_6390,N_6530);
or U6694 (N_6694,N_6434,N_6467);
or U6695 (N_6695,N_6512,N_6523);
nor U6696 (N_6696,N_6337,N_6475);
nor U6697 (N_6697,N_6393,N_6326);
nor U6698 (N_6698,N_6520,N_6333);
or U6699 (N_6699,N_6387,N_6302);
xor U6700 (N_6700,N_6438,N_6496);
and U6701 (N_6701,N_6432,N_6472);
nand U6702 (N_6702,N_6317,N_6411);
or U6703 (N_6703,N_6564,N_6419);
or U6704 (N_6704,N_6353,N_6487);
nor U6705 (N_6705,N_6579,N_6449);
nor U6706 (N_6706,N_6575,N_6526);
nor U6707 (N_6707,N_6525,N_6365);
xor U6708 (N_6708,N_6516,N_6303);
xor U6709 (N_6709,N_6377,N_6359);
or U6710 (N_6710,N_6521,N_6556);
or U6711 (N_6711,N_6505,N_6540);
and U6712 (N_6712,N_6446,N_6324);
and U6713 (N_6713,N_6599,N_6566);
xor U6714 (N_6714,N_6382,N_6355);
nor U6715 (N_6715,N_6510,N_6506);
nand U6716 (N_6716,N_6402,N_6418);
and U6717 (N_6717,N_6445,N_6527);
or U6718 (N_6718,N_6469,N_6484);
xnor U6719 (N_6719,N_6500,N_6553);
nor U6720 (N_6720,N_6426,N_6459);
nor U6721 (N_6721,N_6585,N_6456);
nor U6722 (N_6722,N_6441,N_6341);
nand U6723 (N_6723,N_6518,N_6339);
nor U6724 (N_6724,N_6567,N_6336);
or U6725 (N_6725,N_6440,N_6541);
nor U6726 (N_6726,N_6300,N_6495);
xor U6727 (N_6727,N_6392,N_6561);
and U6728 (N_6728,N_6473,N_6322);
xor U6729 (N_6729,N_6519,N_6312);
and U6730 (N_6730,N_6531,N_6544);
xor U6731 (N_6731,N_6483,N_6414);
nand U6732 (N_6732,N_6338,N_6562);
nand U6733 (N_6733,N_6576,N_6587);
or U6734 (N_6734,N_6436,N_6586);
nor U6735 (N_6735,N_6310,N_6457);
nor U6736 (N_6736,N_6401,N_6367);
xor U6737 (N_6737,N_6360,N_6589);
nand U6738 (N_6738,N_6474,N_6343);
or U6739 (N_6739,N_6330,N_6528);
nor U6740 (N_6740,N_6486,N_6497);
nand U6741 (N_6741,N_6450,N_6369);
nand U6742 (N_6742,N_6596,N_6513);
nand U6743 (N_6743,N_6460,N_6532);
xor U6744 (N_6744,N_6350,N_6454);
nor U6745 (N_6745,N_6593,N_6447);
or U6746 (N_6746,N_6375,N_6503);
nor U6747 (N_6747,N_6424,N_6478);
and U6748 (N_6748,N_6391,N_6578);
xnor U6749 (N_6749,N_6320,N_6315);
or U6750 (N_6750,N_6360,N_6309);
nand U6751 (N_6751,N_6420,N_6344);
xnor U6752 (N_6752,N_6308,N_6486);
or U6753 (N_6753,N_6543,N_6378);
xnor U6754 (N_6754,N_6518,N_6595);
nand U6755 (N_6755,N_6494,N_6352);
nor U6756 (N_6756,N_6406,N_6501);
xor U6757 (N_6757,N_6406,N_6572);
nor U6758 (N_6758,N_6476,N_6379);
and U6759 (N_6759,N_6371,N_6349);
nand U6760 (N_6760,N_6562,N_6589);
nor U6761 (N_6761,N_6414,N_6539);
and U6762 (N_6762,N_6535,N_6437);
nor U6763 (N_6763,N_6339,N_6592);
and U6764 (N_6764,N_6487,N_6457);
and U6765 (N_6765,N_6349,N_6393);
xor U6766 (N_6766,N_6574,N_6573);
and U6767 (N_6767,N_6361,N_6594);
nor U6768 (N_6768,N_6511,N_6472);
xnor U6769 (N_6769,N_6427,N_6507);
nor U6770 (N_6770,N_6583,N_6417);
or U6771 (N_6771,N_6335,N_6354);
nor U6772 (N_6772,N_6465,N_6388);
or U6773 (N_6773,N_6577,N_6505);
or U6774 (N_6774,N_6447,N_6521);
or U6775 (N_6775,N_6477,N_6352);
and U6776 (N_6776,N_6373,N_6508);
or U6777 (N_6777,N_6381,N_6481);
or U6778 (N_6778,N_6541,N_6544);
nand U6779 (N_6779,N_6487,N_6503);
nand U6780 (N_6780,N_6591,N_6322);
and U6781 (N_6781,N_6424,N_6399);
and U6782 (N_6782,N_6400,N_6322);
nor U6783 (N_6783,N_6442,N_6357);
xnor U6784 (N_6784,N_6367,N_6477);
nor U6785 (N_6785,N_6334,N_6573);
xor U6786 (N_6786,N_6571,N_6353);
xnor U6787 (N_6787,N_6397,N_6371);
nand U6788 (N_6788,N_6497,N_6309);
xor U6789 (N_6789,N_6548,N_6590);
and U6790 (N_6790,N_6593,N_6333);
xor U6791 (N_6791,N_6518,N_6393);
nand U6792 (N_6792,N_6520,N_6306);
xnor U6793 (N_6793,N_6312,N_6388);
or U6794 (N_6794,N_6472,N_6583);
nor U6795 (N_6795,N_6434,N_6557);
nand U6796 (N_6796,N_6416,N_6543);
xor U6797 (N_6797,N_6450,N_6585);
nor U6798 (N_6798,N_6488,N_6565);
and U6799 (N_6799,N_6378,N_6344);
and U6800 (N_6800,N_6302,N_6322);
nand U6801 (N_6801,N_6347,N_6368);
or U6802 (N_6802,N_6556,N_6326);
or U6803 (N_6803,N_6430,N_6459);
and U6804 (N_6804,N_6351,N_6572);
nor U6805 (N_6805,N_6350,N_6349);
nor U6806 (N_6806,N_6403,N_6393);
xnor U6807 (N_6807,N_6536,N_6578);
nand U6808 (N_6808,N_6531,N_6397);
nor U6809 (N_6809,N_6411,N_6497);
nor U6810 (N_6810,N_6356,N_6381);
xor U6811 (N_6811,N_6304,N_6323);
nor U6812 (N_6812,N_6481,N_6594);
and U6813 (N_6813,N_6504,N_6484);
nand U6814 (N_6814,N_6509,N_6393);
or U6815 (N_6815,N_6420,N_6461);
and U6816 (N_6816,N_6516,N_6468);
nor U6817 (N_6817,N_6577,N_6543);
and U6818 (N_6818,N_6448,N_6556);
nand U6819 (N_6819,N_6305,N_6376);
xnor U6820 (N_6820,N_6576,N_6366);
or U6821 (N_6821,N_6429,N_6420);
or U6822 (N_6822,N_6569,N_6586);
and U6823 (N_6823,N_6397,N_6388);
and U6824 (N_6824,N_6477,N_6465);
or U6825 (N_6825,N_6490,N_6302);
nor U6826 (N_6826,N_6498,N_6503);
nor U6827 (N_6827,N_6566,N_6338);
xor U6828 (N_6828,N_6541,N_6416);
and U6829 (N_6829,N_6482,N_6545);
nand U6830 (N_6830,N_6539,N_6451);
and U6831 (N_6831,N_6302,N_6530);
nand U6832 (N_6832,N_6370,N_6366);
or U6833 (N_6833,N_6491,N_6585);
and U6834 (N_6834,N_6406,N_6413);
xnor U6835 (N_6835,N_6386,N_6305);
nand U6836 (N_6836,N_6596,N_6351);
and U6837 (N_6837,N_6575,N_6551);
nor U6838 (N_6838,N_6482,N_6489);
nand U6839 (N_6839,N_6387,N_6320);
xor U6840 (N_6840,N_6480,N_6554);
nand U6841 (N_6841,N_6391,N_6598);
or U6842 (N_6842,N_6505,N_6563);
xnor U6843 (N_6843,N_6513,N_6540);
and U6844 (N_6844,N_6442,N_6436);
and U6845 (N_6845,N_6313,N_6491);
and U6846 (N_6846,N_6541,N_6575);
xnor U6847 (N_6847,N_6409,N_6535);
or U6848 (N_6848,N_6529,N_6423);
xor U6849 (N_6849,N_6328,N_6340);
xnor U6850 (N_6850,N_6456,N_6319);
or U6851 (N_6851,N_6517,N_6358);
nor U6852 (N_6852,N_6568,N_6446);
or U6853 (N_6853,N_6424,N_6483);
nand U6854 (N_6854,N_6401,N_6586);
nand U6855 (N_6855,N_6558,N_6389);
nand U6856 (N_6856,N_6583,N_6304);
or U6857 (N_6857,N_6318,N_6547);
or U6858 (N_6858,N_6336,N_6489);
nor U6859 (N_6859,N_6504,N_6486);
xnor U6860 (N_6860,N_6463,N_6381);
nor U6861 (N_6861,N_6448,N_6492);
nor U6862 (N_6862,N_6557,N_6468);
and U6863 (N_6863,N_6594,N_6357);
and U6864 (N_6864,N_6536,N_6424);
xor U6865 (N_6865,N_6420,N_6300);
or U6866 (N_6866,N_6573,N_6527);
and U6867 (N_6867,N_6477,N_6441);
or U6868 (N_6868,N_6359,N_6590);
or U6869 (N_6869,N_6425,N_6417);
and U6870 (N_6870,N_6474,N_6553);
and U6871 (N_6871,N_6564,N_6453);
nor U6872 (N_6872,N_6428,N_6308);
and U6873 (N_6873,N_6312,N_6565);
nand U6874 (N_6874,N_6550,N_6546);
nand U6875 (N_6875,N_6412,N_6582);
nand U6876 (N_6876,N_6465,N_6398);
nand U6877 (N_6877,N_6510,N_6463);
nand U6878 (N_6878,N_6515,N_6535);
nor U6879 (N_6879,N_6481,N_6522);
nand U6880 (N_6880,N_6375,N_6451);
or U6881 (N_6881,N_6390,N_6538);
xnor U6882 (N_6882,N_6306,N_6511);
or U6883 (N_6883,N_6509,N_6382);
nor U6884 (N_6884,N_6401,N_6513);
xor U6885 (N_6885,N_6409,N_6484);
nand U6886 (N_6886,N_6490,N_6492);
or U6887 (N_6887,N_6350,N_6499);
and U6888 (N_6888,N_6418,N_6444);
xor U6889 (N_6889,N_6551,N_6531);
nor U6890 (N_6890,N_6550,N_6316);
nor U6891 (N_6891,N_6454,N_6592);
nor U6892 (N_6892,N_6308,N_6468);
xnor U6893 (N_6893,N_6508,N_6502);
nand U6894 (N_6894,N_6538,N_6419);
or U6895 (N_6895,N_6363,N_6583);
nand U6896 (N_6896,N_6326,N_6369);
nand U6897 (N_6897,N_6572,N_6519);
and U6898 (N_6898,N_6512,N_6444);
nor U6899 (N_6899,N_6357,N_6528);
nor U6900 (N_6900,N_6801,N_6678);
xor U6901 (N_6901,N_6860,N_6788);
nand U6902 (N_6902,N_6822,N_6893);
nand U6903 (N_6903,N_6891,N_6815);
nand U6904 (N_6904,N_6761,N_6866);
nor U6905 (N_6905,N_6722,N_6621);
nor U6906 (N_6906,N_6754,N_6870);
xnor U6907 (N_6907,N_6609,N_6718);
and U6908 (N_6908,N_6613,N_6742);
xnor U6909 (N_6909,N_6786,N_6881);
nor U6910 (N_6910,N_6819,N_6804);
or U6911 (N_6911,N_6665,N_6715);
nand U6912 (N_6912,N_6820,N_6651);
nand U6913 (N_6913,N_6646,N_6852);
or U6914 (N_6914,N_6814,N_6809);
nand U6915 (N_6915,N_6849,N_6762);
or U6916 (N_6916,N_6818,N_6636);
or U6917 (N_6917,N_6679,N_6812);
and U6918 (N_6918,N_6680,N_6791);
xor U6919 (N_6919,N_6682,N_6765);
xor U6920 (N_6920,N_6629,N_6645);
nand U6921 (N_6921,N_6630,N_6817);
nand U6922 (N_6922,N_6737,N_6760);
xor U6923 (N_6923,N_6769,N_6744);
nor U6924 (N_6924,N_6720,N_6698);
and U6925 (N_6925,N_6657,N_6787);
nor U6926 (N_6926,N_6869,N_6633);
and U6927 (N_6927,N_6702,N_6714);
xnor U6928 (N_6928,N_6644,N_6839);
nor U6929 (N_6929,N_6838,N_6634);
and U6930 (N_6930,N_6871,N_6894);
xnor U6931 (N_6931,N_6741,N_6846);
and U6932 (N_6932,N_6885,N_6851);
nor U6933 (N_6933,N_6616,N_6626);
nor U6934 (N_6934,N_6693,N_6705);
nand U6935 (N_6935,N_6627,N_6664);
nor U6936 (N_6936,N_6863,N_6631);
xnor U6937 (N_6937,N_6748,N_6637);
xnor U6938 (N_6938,N_6642,N_6623);
or U6939 (N_6939,N_6696,N_6811);
or U6940 (N_6940,N_6619,N_6607);
nand U6941 (N_6941,N_6602,N_6654);
and U6942 (N_6942,N_6643,N_6873);
xor U6943 (N_6943,N_6746,N_6600);
xnor U6944 (N_6944,N_6661,N_6777);
and U6945 (N_6945,N_6688,N_6671);
nand U6946 (N_6946,N_6875,N_6723);
xnor U6947 (N_6947,N_6675,N_6898);
nand U6948 (N_6948,N_6649,N_6874);
or U6949 (N_6949,N_6740,N_6750);
nand U6950 (N_6950,N_6897,N_6677);
xor U6951 (N_6951,N_6731,N_6794);
and U6952 (N_6952,N_6773,N_6694);
xnor U6953 (N_6953,N_6782,N_6758);
nand U6954 (N_6954,N_6639,N_6858);
or U6955 (N_6955,N_6796,N_6877);
xnor U6956 (N_6956,N_6895,N_6896);
nor U6957 (N_6957,N_6800,N_6721);
or U6958 (N_6958,N_6666,N_6681);
xnor U6959 (N_6959,N_6805,N_6756);
or U6960 (N_6960,N_6848,N_6717);
nand U6961 (N_6961,N_6727,N_6847);
nand U6962 (N_6962,N_6628,N_6691);
xnor U6963 (N_6963,N_6669,N_6662);
or U6964 (N_6964,N_6768,N_6807);
nand U6965 (N_6965,N_6729,N_6832);
and U6966 (N_6966,N_6776,N_6689);
and U6967 (N_6967,N_6763,N_6659);
nand U6968 (N_6968,N_6710,N_6620);
xor U6969 (N_6969,N_6861,N_6683);
nand U6970 (N_6970,N_6690,N_6615);
xnor U6971 (N_6971,N_6638,N_6658);
or U6972 (N_6972,N_6617,N_6855);
nand U6973 (N_6973,N_6808,N_6738);
nand U6974 (N_6974,N_6882,N_6719);
nor U6975 (N_6975,N_6784,N_6868);
xor U6976 (N_6976,N_6810,N_6663);
and U6977 (N_6977,N_6771,N_6752);
or U6978 (N_6978,N_6883,N_6793);
xnor U6979 (N_6979,N_6747,N_6701);
nor U6980 (N_6980,N_6608,N_6840);
or U6981 (N_6981,N_6716,N_6635);
nand U6982 (N_6982,N_6684,N_6803);
or U6983 (N_6983,N_6798,N_6655);
nand U6984 (N_6984,N_6745,N_6708);
nor U6985 (N_6985,N_6841,N_6743);
and U6986 (N_6986,N_6700,N_6753);
or U6987 (N_6987,N_6857,N_6844);
nand U6988 (N_6988,N_6706,N_6755);
or U6989 (N_6989,N_6884,N_6880);
and U6990 (N_6990,N_6618,N_6610);
nand U6991 (N_6991,N_6835,N_6892);
or U6992 (N_6992,N_6888,N_6843);
and U6993 (N_6993,N_6704,N_6890);
nor U6994 (N_6994,N_6640,N_6887);
nand U6995 (N_6995,N_6845,N_6699);
and U6996 (N_6996,N_6781,N_6648);
and U6997 (N_6997,N_6790,N_6695);
xnor U6998 (N_6998,N_6734,N_6886);
nand U6999 (N_6999,N_6842,N_6673);
and U7000 (N_7000,N_6672,N_6878);
or U7001 (N_7001,N_6826,N_6759);
nand U7002 (N_7002,N_6879,N_6725);
or U7003 (N_7003,N_6772,N_6732);
and U7004 (N_7004,N_6603,N_6606);
nor U7005 (N_7005,N_6806,N_6766);
xor U7006 (N_7006,N_6712,N_6624);
nand U7007 (N_7007,N_6831,N_6859);
nor U7008 (N_7008,N_6823,N_6876);
nand U7009 (N_7009,N_6780,N_6821);
or U7010 (N_7010,N_6865,N_6856);
and U7011 (N_7011,N_6816,N_6726);
and U7012 (N_7012,N_6676,N_6601);
nor U7013 (N_7013,N_6789,N_6674);
or U7014 (N_7014,N_6656,N_6853);
or U7015 (N_7015,N_6647,N_6774);
or U7016 (N_7016,N_6797,N_6829);
nor U7017 (N_7017,N_6828,N_6795);
nor U7018 (N_7018,N_6799,N_6632);
and U7019 (N_7019,N_6813,N_6783);
xor U7020 (N_7020,N_6739,N_6779);
nor U7021 (N_7021,N_6889,N_6770);
or U7022 (N_7022,N_6605,N_6736);
nor U7023 (N_7023,N_6730,N_6650);
nand U7024 (N_7024,N_6836,N_6713);
xor U7025 (N_7025,N_6854,N_6792);
xnor U7026 (N_7026,N_6830,N_6625);
and U7027 (N_7027,N_6707,N_6687);
and U7028 (N_7028,N_6709,N_6653);
nor U7029 (N_7029,N_6667,N_6837);
nand U7030 (N_7030,N_6641,N_6614);
nor U7031 (N_7031,N_6834,N_6867);
and U7032 (N_7032,N_6757,N_6785);
nand U7033 (N_7033,N_6827,N_6692);
and U7034 (N_7034,N_6724,N_6611);
and U7035 (N_7035,N_6749,N_6703);
or U7036 (N_7036,N_6711,N_6751);
nand U7037 (N_7037,N_6668,N_6697);
and U7038 (N_7038,N_6686,N_6862);
or U7039 (N_7039,N_6685,N_6652);
and U7040 (N_7040,N_6825,N_6833);
or U7041 (N_7041,N_6612,N_6824);
and U7042 (N_7042,N_6899,N_6733);
nor U7043 (N_7043,N_6778,N_6850);
nor U7044 (N_7044,N_6670,N_6802);
and U7045 (N_7045,N_6728,N_6735);
and U7046 (N_7046,N_6764,N_6604);
xor U7047 (N_7047,N_6872,N_6660);
nor U7048 (N_7048,N_6622,N_6864);
nor U7049 (N_7049,N_6767,N_6775);
nand U7050 (N_7050,N_6633,N_6619);
or U7051 (N_7051,N_6888,N_6720);
and U7052 (N_7052,N_6847,N_6859);
and U7053 (N_7053,N_6739,N_6644);
and U7054 (N_7054,N_6808,N_6649);
nand U7055 (N_7055,N_6623,N_6726);
xnor U7056 (N_7056,N_6714,N_6836);
xor U7057 (N_7057,N_6773,N_6678);
xor U7058 (N_7058,N_6854,N_6850);
xor U7059 (N_7059,N_6616,N_6610);
and U7060 (N_7060,N_6816,N_6783);
and U7061 (N_7061,N_6872,N_6713);
and U7062 (N_7062,N_6772,N_6703);
and U7063 (N_7063,N_6803,N_6637);
nor U7064 (N_7064,N_6674,N_6711);
and U7065 (N_7065,N_6886,N_6865);
nand U7066 (N_7066,N_6715,N_6820);
xor U7067 (N_7067,N_6776,N_6669);
or U7068 (N_7068,N_6791,N_6662);
and U7069 (N_7069,N_6712,N_6646);
or U7070 (N_7070,N_6875,N_6665);
or U7071 (N_7071,N_6753,N_6894);
xnor U7072 (N_7072,N_6734,N_6876);
and U7073 (N_7073,N_6876,N_6832);
and U7074 (N_7074,N_6761,N_6753);
or U7075 (N_7075,N_6883,N_6740);
nor U7076 (N_7076,N_6895,N_6795);
nor U7077 (N_7077,N_6801,N_6693);
nand U7078 (N_7078,N_6636,N_6616);
nand U7079 (N_7079,N_6700,N_6730);
nand U7080 (N_7080,N_6673,N_6827);
and U7081 (N_7081,N_6865,N_6698);
or U7082 (N_7082,N_6766,N_6835);
nand U7083 (N_7083,N_6615,N_6898);
and U7084 (N_7084,N_6819,N_6724);
nand U7085 (N_7085,N_6710,N_6742);
or U7086 (N_7086,N_6891,N_6647);
nor U7087 (N_7087,N_6698,N_6877);
and U7088 (N_7088,N_6816,N_6757);
and U7089 (N_7089,N_6615,N_6844);
nand U7090 (N_7090,N_6888,N_6858);
xnor U7091 (N_7091,N_6807,N_6701);
or U7092 (N_7092,N_6635,N_6659);
xor U7093 (N_7093,N_6714,N_6711);
and U7094 (N_7094,N_6856,N_6828);
or U7095 (N_7095,N_6612,N_6676);
nand U7096 (N_7096,N_6690,N_6867);
and U7097 (N_7097,N_6766,N_6868);
nand U7098 (N_7098,N_6864,N_6608);
nand U7099 (N_7099,N_6615,N_6715);
nand U7100 (N_7100,N_6685,N_6718);
and U7101 (N_7101,N_6838,N_6637);
or U7102 (N_7102,N_6863,N_6694);
nand U7103 (N_7103,N_6889,N_6799);
nor U7104 (N_7104,N_6639,N_6712);
or U7105 (N_7105,N_6641,N_6722);
nand U7106 (N_7106,N_6817,N_6656);
xnor U7107 (N_7107,N_6754,N_6621);
or U7108 (N_7108,N_6856,N_6780);
nand U7109 (N_7109,N_6882,N_6880);
xnor U7110 (N_7110,N_6792,N_6757);
nor U7111 (N_7111,N_6710,N_6607);
nand U7112 (N_7112,N_6713,N_6851);
nand U7113 (N_7113,N_6856,N_6617);
nor U7114 (N_7114,N_6701,N_6718);
xor U7115 (N_7115,N_6810,N_6762);
or U7116 (N_7116,N_6887,N_6760);
nand U7117 (N_7117,N_6713,N_6882);
nor U7118 (N_7118,N_6637,N_6740);
xor U7119 (N_7119,N_6679,N_6641);
nand U7120 (N_7120,N_6698,N_6611);
xor U7121 (N_7121,N_6606,N_6700);
nand U7122 (N_7122,N_6628,N_6654);
nor U7123 (N_7123,N_6805,N_6604);
or U7124 (N_7124,N_6652,N_6739);
or U7125 (N_7125,N_6776,N_6876);
nand U7126 (N_7126,N_6826,N_6868);
xor U7127 (N_7127,N_6708,N_6718);
nor U7128 (N_7128,N_6871,N_6723);
nor U7129 (N_7129,N_6699,N_6776);
xor U7130 (N_7130,N_6874,N_6636);
xnor U7131 (N_7131,N_6763,N_6857);
nand U7132 (N_7132,N_6624,N_6688);
nand U7133 (N_7133,N_6682,N_6749);
or U7134 (N_7134,N_6666,N_6607);
or U7135 (N_7135,N_6802,N_6692);
xor U7136 (N_7136,N_6806,N_6888);
xor U7137 (N_7137,N_6748,N_6761);
nand U7138 (N_7138,N_6671,N_6795);
or U7139 (N_7139,N_6624,N_6749);
nand U7140 (N_7140,N_6768,N_6650);
xnor U7141 (N_7141,N_6809,N_6889);
nand U7142 (N_7142,N_6665,N_6643);
and U7143 (N_7143,N_6891,N_6816);
xnor U7144 (N_7144,N_6818,N_6851);
and U7145 (N_7145,N_6758,N_6889);
nand U7146 (N_7146,N_6850,N_6652);
or U7147 (N_7147,N_6694,N_6734);
xnor U7148 (N_7148,N_6619,N_6758);
or U7149 (N_7149,N_6661,N_6623);
or U7150 (N_7150,N_6663,N_6622);
or U7151 (N_7151,N_6822,N_6873);
or U7152 (N_7152,N_6694,N_6759);
nor U7153 (N_7153,N_6607,N_6610);
xnor U7154 (N_7154,N_6872,N_6791);
and U7155 (N_7155,N_6808,N_6622);
xor U7156 (N_7156,N_6720,N_6736);
or U7157 (N_7157,N_6733,N_6632);
or U7158 (N_7158,N_6708,N_6801);
nor U7159 (N_7159,N_6625,N_6757);
xnor U7160 (N_7160,N_6679,N_6640);
nand U7161 (N_7161,N_6875,N_6882);
and U7162 (N_7162,N_6751,N_6621);
xor U7163 (N_7163,N_6633,N_6636);
and U7164 (N_7164,N_6771,N_6809);
nor U7165 (N_7165,N_6696,N_6800);
or U7166 (N_7166,N_6858,N_6665);
or U7167 (N_7167,N_6839,N_6742);
nand U7168 (N_7168,N_6631,N_6834);
xnor U7169 (N_7169,N_6769,N_6704);
or U7170 (N_7170,N_6631,N_6806);
or U7171 (N_7171,N_6729,N_6898);
xnor U7172 (N_7172,N_6721,N_6867);
and U7173 (N_7173,N_6662,N_6741);
or U7174 (N_7174,N_6704,N_6755);
nor U7175 (N_7175,N_6714,N_6838);
xnor U7176 (N_7176,N_6753,N_6843);
xnor U7177 (N_7177,N_6837,N_6676);
xor U7178 (N_7178,N_6722,N_6882);
nand U7179 (N_7179,N_6617,N_6621);
nor U7180 (N_7180,N_6603,N_6886);
and U7181 (N_7181,N_6723,N_6788);
nor U7182 (N_7182,N_6651,N_6725);
nand U7183 (N_7183,N_6822,N_6601);
and U7184 (N_7184,N_6625,N_6847);
and U7185 (N_7185,N_6718,N_6856);
or U7186 (N_7186,N_6660,N_6834);
and U7187 (N_7187,N_6712,N_6844);
nor U7188 (N_7188,N_6605,N_6841);
nor U7189 (N_7189,N_6856,N_6884);
and U7190 (N_7190,N_6687,N_6660);
or U7191 (N_7191,N_6774,N_6732);
xor U7192 (N_7192,N_6616,N_6685);
or U7193 (N_7193,N_6719,N_6645);
nor U7194 (N_7194,N_6894,N_6854);
nor U7195 (N_7195,N_6788,N_6636);
nor U7196 (N_7196,N_6606,N_6828);
xor U7197 (N_7197,N_6818,N_6692);
or U7198 (N_7198,N_6811,N_6880);
and U7199 (N_7199,N_6744,N_6723);
or U7200 (N_7200,N_6962,N_7048);
or U7201 (N_7201,N_6918,N_7196);
nand U7202 (N_7202,N_7109,N_7186);
nand U7203 (N_7203,N_7000,N_7027);
nor U7204 (N_7204,N_7056,N_6964);
and U7205 (N_7205,N_6936,N_7117);
xor U7206 (N_7206,N_7033,N_7185);
nor U7207 (N_7207,N_6900,N_7059);
nor U7208 (N_7208,N_7141,N_7014);
xnor U7209 (N_7209,N_6973,N_7124);
and U7210 (N_7210,N_6991,N_7040);
or U7211 (N_7211,N_6949,N_6954);
xnor U7212 (N_7212,N_7074,N_6980);
nor U7213 (N_7213,N_7022,N_7143);
nand U7214 (N_7214,N_6955,N_7049);
and U7215 (N_7215,N_6916,N_6914);
nor U7216 (N_7216,N_6913,N_6971);
or U7217 (N_7217,N_7197,N_6939);
nand U7218 (N_7218,N_6909,N_7144);
or U7219 (N_7219,N_6929,N_6968);
nand U7220 (N_7220,N_7047,N_7050);
nor U7221 (N_7221,N_7007,N_7035);
and U7222 (N_7222,N_6998,N_7176);
nor U7223 (N_7223,N_7188,N_7189);
xnor U7224 (N_7224,N_7094,N_7111);
or U7225 (N_7225,N_7116,N_6926);
xnor U7226 (N_7226,N_7023,N_7172);
xor U7227 (N_7227,N_7042,N_7164);
xor U7228 (N_7228,N_7129,N_7067);
nand U7229 (N_7229,N_7183,N_7063);
nand U7230 (N_7230,N_7003,N_6951);
or U7231 (N_7231,N_7179,N_6983);
nand U7232 (N_7232,N_7012,N_7066);
xnor U7233 (N_7233,N_6924,N_7153);
nand U7234 (N_7234,N_7140,N_6905);
or U7235 (N_7235,N_7064,N_7145);
nand U7236 (N_7236,N_7163,N_6935);
or U7237 (N_7237,N_7021,N_7118);
xnor U7238 (N_7238,N_6906,N_7070);
nor U7239 (N_7239,N_6985,N_7011);
nand U7240 (N_7240,N_7147,N_6903);
or U7241 (N_7241,N_7135,N_6981);
xnor U7242 (N_7242,N_6979,N_7092);
or U7243 (N_7243,N_7131,N_7065);
or U7244 (N_7244,N_7044,N_7103);
and U7245 (N_7245,N_7075,N_7113);
nor U7246 (N_7246,N_7087,N_7193);
or U7247 (N_7247,N_7194,N_7198);
nor U7248 (N_7248,N_7170,N_7130);
nor U7249 (N_7249,N_7161,N_7122);
nand U7250 (N_7250,N_7020,N_7032);
xor U7251 (N_7251,N_6992,N_7171);
xnor U7252 (N_7252,N_7138,N_7114);
nor U7253 (N_7253,N_6950,N_7098);
and U7254 (N_7254,N_6943,N_6970);
nor U7255 (N_7255,N_7015,N_7051);
and U7256 (N_7256,N_6944,N_7136);
or U7257 (N_7257,N_7085,N_6908);
xor U7258 (N_7258,N_7177,N_6948);
nor U7259 (N_7259,N_7181,N_7025);
nand U7260 (N_7260,N_7062,N_7110);
nor U7261 (N_7261,N_7091,N_7156);
or U7262 (N_7262,N_7013,N_6915);
or U7263 (N_7263,N_7008,N_6967);
and U7264 (N_7264,N_7061,N_7101);
nand U7265 (N_7265,N_7175,N_7083);
xnor U7266 (N_7266,N_7082,N_6957);
nor U7267 (N_7267,N_6987,N_7168);
or U7268 (N_7268,N_7010,N_7099);
or U7269 (N_7269,N_6988,N_7076);
nand U7270 (N_7270,N_7187,N_6947);
or U7271 (N_7271,N_7121,N_7126);
xor U7272 (N_7272,N_7072,N_7195);
and U7273 (N_7273,N_7055,N_7173);
and U7274 (N_7274,N_7115,N_6999);
nand U7275 (N_7275,N_6974,N_7134);
or U7276 (N_7276,N_7142,N_7026);
nor U7277 (N_7277,N_7146,N_7086);
nor U7278 (N_7278,N_6972,N_7096);
or U7279 (N_7279,N_7159,N_7155);
and U7280 (N_7280,N_6978,N_7192);
nor U7281 (N_7281,N_7037,N_7038);
nand U7282 (N_7282,N_7057,N_7154);
or U7283 (N_7283,N_6933,N_6963);
nor U7284 (N_7284,N_7018,N_7081);
nor U7285 (N_7285,N_7073,N_6965);
nand U7286 (N_7286,N_6958,N_7152);
nand U7287 (N_7287,N_7105,N_7184);
and U7288 (N_7288,N_7041,N_7001);
and U7289 (N_7289,N_7004,N_7100);
and U7290 (N_7290,N_6959,N_7123);
and U7291 (N_7291,N_7199,N_7137);
nand U7292 (N_7292,N_7052,N_7149);
nand U7293 (N_7293,N_7132,N_7165);
nand U7294 (N_7294,N_7178,N_7106);
and U7295 (N_7295,N_6925,N_6912);
and U7296 (N_7296,N_7191,N_7166);
and U7297 (N_7297,N_6960,N_6984);
nor U7298 (N_7298,N_7182,N_7016);
or U7299 (N_7299,N_6934,N_7039);
xor U7300 (N_7300,N_7120,N_6928);
and U7301 (N_7301,N_7167,N_6956);
xnor U7302 (N_7302,N_7029,N_7180);
nand U7303 (N_7303,N_7169,N_7005);
and U7304 (N_7304,N_6993,N_6907);
nand U7305 (N_7305,N_6953,N_7095);
or U7306 (N_7306,N_7160,N_7019);
nand U7307 (N_7307,N_6995,N_6942);
xor U7308 (N_7308,N_7006,N_6911);
nor U7309 (N_7309,N_7190,N_6952);
and U7310 (N_7310,N_6927,N_7088);
nand U7311 (N_7311,N_7079,N_7071);
and U7312 (N_7312,N_6904,N_6994);
and U7313 (N_7313,N_7157,N_6946);
or U7314 (N_7314,N_6937,N_7017);
nor U7315 (N_7315,N_6923,N_6922);
and U7316 (N_7316,N_7151,N_7058);
xnor U7317 (N_7317,N_6945,N_7009);
xor U7318 (N_7318,N_7119,N_7080);
xnor U7319 (N_7319,N_7139,N_7158);
xnor U7320 (N_7320,N_6901,N_6966);
and U7321 (N_7321,N_6989,N_7102);
xor U7322 (N_7322,N_7069,N_6996);
and U7323 (N_7323,N_7097,N_7174);
xor U7324 (N_7324,N_7108,N_6940);
nand U7325 (N_7325,N_6930,N_6921);
xnor U7326 (N_7326,N_7053,N_7034);
xnor U7327 (N_7327,N_6986,N_6917);
or U7328 (N_7328,N_6982,N_6902);
nand U7329 (N_7329,N_6977,N_7084);
and U7330 (N_7330,N_7148,N_7104);
xnor U7331 (N_7331,N_6997,N_7093);
nor U7332 (N_7332,N_6932,N_6920);
nand U7333 (N_7333,N_7045,N_7127);
nand U7334 (N_7334,N_7077,N_6975);
nand U7335 (N_7335,N_7150,N_6990);
nand U7336 (N_7336,N_7036,N_6910);
or U7337 (N_7337,N_7046,N_6938);
and U7338 (N_7338,N_6976,N_7024);
nand U7339 (N_7339,N_7031,N_7112);
nand U7340 (N_7340,N_7054,N_6919);
or U7341 (N_7341,N_7162,N_7002);
xor U7342 (N_7342,N_7043,N_7028);
xnor U7343 (N_7343,N_7068,N_6941);
nor U7344 (N_7344,N_6961,N_7133);
nand U7345 (N_7345,N_6931,N_7125);
or U7346 (N_7346,N_7107,N_6969);
and U7347 (N_7347,N_7089,N_7078);
and U7348 (N_7348,N_7090,N_7128);
xor U7349 (N_7349,N_7030,N_7060);
nand U7350 (N_7350,N_6910,N_7061);
xor U7351 (N_7351,N_7086,N_6947);
or U7352 (N_7352,N_6936,N_7112);
and U7353 (N_7353,N_7070,N_7155);
and U7354 (N_7354,N_7097,N_7175);
and U7355 (N_7355,N_7072,N_7004);
or U7356 (N_7356,N_7032,N_7071);
or U7357 (N_7357,N_7103,N_7150);
xor U7358 (N_7358,N_7196,N_7023);
or U7359 (N_7359,N_7106,N_7155);
and U7360 (N_7360,N_7006,N_6945);
or U7361 (N_7361,N_7150,N_7016);
nand U7362 (N_7362,N_7103,N_7002);
and U7363 (N_7363,N_7101,N_7174);
xor U7364 (N_7364,N_6999,N_7194);
or U7365 (N_7365,N_7113,N_7092);
xnor U7366 (N_7366,N_7186,N_7150);
nand U7367 (N_7367,N_6988,N_7187);
nand U7368 (N_7368,N_7065,N_6904);
and U7369 (N_7369,N_7063,N_7189);
or U7370 (N_7370,N_6973,N_7040);
and U7371 (N_7371,N_7074,N_7054);
xnor U7372 (N_7372,N_7079,N_7193);
nor U7373 (N_7373,N_7197,N_7100);
nand U7374 (N_7374,N_7199,N_7076);
or U7375 (N_7375,N_6929,N_7119);
nor U7376 (N_7376,N_7117,N_7168);
and U7377 (N_7377,N_6955,N_7166);
and U7378 (N_7378,N_7121,N_7175);
nor U7379 (N_7379,N_7066,N_7085);
xor U7380 (N_7380,N_7132,N_7074);
nor U7381 (N_7381,N_7077,N_7185);
and U7382 (N_7382,N_7035,N_7070);
or U7383 (N_7383,N_6980,N_7165);
nand U7384 (N_7384,N_7067,N_7046);
nand U7385 (N_7385,N_7052,N_7068);
or U7386 (N_7386,N_6912,N_7058);
nand U7387 (N_7387,N_6980,N_6923);
nand U7388 (N_7388,N_7127,N_6915);
xnor U7389 (N_7389,N_7106,N_6997);
xnor U7390 (N_7390,N_6926,N_6921);
nor U7391 (N_7391,N_7127,N_7156);
or U7392 (N_7392,N_7013,N_7090);
and U7393 (N_7393,N_7102,N_7044);
or U7394 (N_7394,N_6974,N_6989);
and U7395 (N_7395,N_7182,N_6943);
nand U7396 (N_7396,N_7047,N_7157);
xor U7397 (N_7397,N_6936,N_7028);
nand U7398 (N_7398,N_7065,N_7179);
and U7399 (N_7399,N_6924,N_6960);
and U7400 (N_7400,N_7110,N_7077);
nor U7401 (N_7401,N_7070,N_7099);
nor U7402 (N_7402,N_7074,N_7083);
or U7403 (N_7403,N_7057,N_7076);
xnor U7404 (N_7404,N_7095,N_7027);
and U7405 (N_7405,N_6905,N_6989);
nor U7406 (N_7406,N_6938,N_6998);
nor U7407 (N_7407,N_7009,N_7056);
xnor U7408 (N_7408,N_7029,N_6938);
and U7409 (N_7409,N_7182,N_6940);
nand U7410 (N_7410,N_7145,N_7116);
nand U7411 (N_7411,N_7111,N_6920);
nor U7412 (N_7412,N_6959,N_6972);
nand U7413 (N_7413,N_7083,N_7159);
or U7414 (N_7414,N_6934,N_7164);
or U7415 (N_7415,N_6981,N_7034);
nor U7416 (N_7416,N_6934,N_6939);
nand U7417 (N_7417,N_7114,N_6914);
and U7418 (N_7418,N_7174,N_6907);
or U7419 (N_7419,N_7187,N_6985);
nor U7420 (N_7420,N_7130,N_7153);
or U7421 (N_7421,N_6953,N_7159);
nor U7422 (N_7422,N_6934,N_7025);
nand U7423 (N_7423,N_7196,N_7184);
or U7424 (N_7424,N_6924,N_7092);
nor U7425 (N_7425,N_7054,N_6901);
nor U7426 (N_7426,N_6930,N_7115);
xnor U7427 (N_7427,N_6952,N_7123);
nor U7428 (N_7428,N_6985,N_7049);
or U7429 (N_7429,N_7017,N_6924);
or U7430 (N_7430,N_7176,N_6973);
nand U7431 (N_7431,N_7177,N_7009);
xor U7432 (N_7432,N_7083,N_7095);
xnor U7433 (N_7433,N_6971,N_7001);
xnor U7434 (N_7434,N_6973,N_7091);
nand U7435 (N_7435,N_6979,N_7099);
or U7436 (N_7436,N_6923,N_7025);
nor U7437 (N_7437,N_7046,N_7129);
nor U7438 (N_7438,N_6973,N_7000);
xnor U7439 (N_7439,N_6948,N_7032);
or U7440 (N_7440,N_7187,N_6960);
nand U7441 (N_7441,N_7196,N_6950);
nand U7442 (N_7442,N_6903,N_7183);
nand U7443 (N_7443,N_6964,N_7024);
nor U7444 (N_7444,N_7009,N_6957);
and U7445 (N_7445,N_7017,N_7057);
or U7446 (N_7446,N_7195,N_7158);
and U7447 (N_7447,N_7038,N_7122);
nand U7448 (N_7448,N_7077,N_6949);
or U7449 (N_7449,N_7193,N_6951);
nand U7450 (N_7450,N_6918,N_7127);
nor U7451 (N_7451,N_7094,N_7188);
and U7452 (N_7452,N_7109,N_6983);
nor U7453 (N_7453,N_7157,N_6954);
nor U7454 (N_7454,N_6985,N_7084);
or U7455 (N_7455,N_7155,N_6918);
or U7456 (N_7456,N_7097,N_7125);
and U7457 (N_7457,N_7054,N_7199);
nand U7458 (N_7458,N_6949,N_7079);
xnor U7459 (N_7459,N_7029,N_7005);
and U7460 (N_7460,N_7074,N_7124);
nor U7461 (N_7461,N_6976,N_7067);
and U7462 (N_7462,N_6975,N_6950);
or U7463 (N_7463,N_7073,N_7079);
nand U7464 (N_7464,N_6912,N_7000);
or U7465 (N_7465,N_7050,N_7087);
or U7466 (N_7466,N_6935,N_7170);
xnor U7467 (N_7467,N_7132,N_6909);
nor U7468 (N_7468,N_7139,N_6917);
nor U7469 (N_7469,N_7023,N_7099);
nand U7470 (N_7470,N_6944,N_6943);
and U7471 (N_7471,N_7018,N_6911);
or U7472 (N_7472,N_7100,N_7122);
xnor U7473 (N_7473,N_7174,N_7145);
and U7474 (N_7474,N_7149,N_6942);
or U7475 (N_7475,N_7172,N_6959);
nand U7476 (N_7476,N_6931,N_7131);
nor U7477 (N_7477,N_6944,N_7040);
nor U7478 (N_7478,N_7184,N_6954);
xor U7479 (N_7479,N_6985,N_6956);
or U7480 (N_7480,N_7021,N_7101);
nor U7481 (N_7481,N_7191,N_6981);
and U7482 (N_7482,N_7044,N_6989);
xor U7483 (N_7483,N_7176,N_6939);
nor U7484 (N_7484,N_7054,N_6994);
nor U7485 (N_7485,N_7131,N_7032);
nand U7486 (N_7486,N_6987,N_6931);
and U7487 (N_7487,N_7093,N_6922);
nand U7488 (N_7488,N_6917,N_6914);
and U7489 (N_7489,N_7088,N_6980);
xor U7490 (N_7490,N_7133,N_7107);
nand U7491 (N_7491,N_7141,N_7005);
or U7492 (N_7492,N_6954,N_7183);
xor U7493 (N_7493,N_7005,N_7108);
xnor U7494 (N_7494,N_7090,N_7059);
nor U7495 (N_7495,N_6925,N_7042);
nor U7496 (N_7496,N_7173,N_7099);
and U7497 (N_7497,N_6902,N_7123);
and U7498 (N_7498,N_6925,N_7170);
and U7499 (N_7499,N_7141,N_7137);
xnor U7500 (N_7500,N_7478,N_7465);
nand U7501 (N_7501,N_7460,N_7380);
xor U7502 (N_7502,N_7336,N_7368);
xnor U7503 (N_7503,N_7260,N_7303);
nor U7504 (N_7504,N_7337,N_7376);
nor U7505 (N_7505,N_7426,N_7239);
xor U7506 (N_7506,N_7348,N_7206);
and U7507 (N_7507,N_7231,N_7497);
nor U7508 (N_7508,N_7405,N_7471);
and U7509 (N_7509,N_7383,N_7322);
nand U7510 (N_7510,N_7352,N_7272);
nand U7511 (N_7511,N_7452,N_7349);
nand U7512 (N_7512,N_7274,N_7398);
or U7513 (N_7513,N_7312,N_7411);
and U7514 (N_7514,N_7433,N_7448);
or U7515 (N_7515,N_7404,N_7384);
or U7516 (N_7516,N_7232,N_7418);
nor U7517 (N_7517,N_7373,N_7245);
xor U7518 (N_7518,N_7249,N_7314);
nor U7519 (N_7519,N_7470,N_7489);
nor U7520 (N_7520,N_7356,N_7269);
and U7521 (N_7521,N_7412,N_7354);
xnor U7522 (N_7522,N_7391,N_7325);
or U7523 (N_7523,N_7227,N_7487);
or U7524 (N_7524,N_7221,N_7277);
or U7525 (N_7525,N_7342,N_7392);
and U7526 (N_7526,N_7488,N_7270);
xor U7527 (N_7527,N_7493,N_7358);
or U7528 (N_7528,N_7390,N_7324);
nand U7529 (N_7529,N_7297,N_7319);
nand U7530 (N_7530,N_7375,N_7455);
nor U7531 (N_7531,N_7468,N_7399);
nor U7532 (N_7532,N_7236,N_7402);
and U7533 (N_7533,N_7369,N_7432);
xor U7534 (N_7534,N_7450,N_7428);
xnor U7535 (N_7535,N_7326,N_7273);
xnor U7536 (N_7536,N_7279,N_7423);
or U7537 (N_7537,N_7265,N_7284);
nand U7538 (N_7538,N_7422,N_7440);
nand U7539 (N_7539,N_7256,N_7299);
nand U7540 (N_7540,N_7327,N_7400);
and U7541 (N_7541,N_7222,N_7242);
and U7542 (N_7542,N_7357,N_7479);
or U7543 (N_7543,N_7481,N_7235);
nor U7544 (N_7544,N_7301,N_7309);
or U7545 (N_7545,N_7438,N_7371);
nand U7546 (N_7546,N_7499,N_7469);
xnor U7547 (N_7547,N_7416,N_7291);
nor U7548 (N_7548,N_7425,N_7292);
and U7549 (N_7549,N_7230,N_7459);
or U7550 (N_7550,N_7344,N_7238);
or U7551 (N_7551,N_7341,N_7490);
xnor U7552 (N_7552,N_7364,N_7208);
nand U7553 (N_7553,N_7494,N_7262);
and U7554 (N_7554,N_7317,N_7485);
or U7555 (N_7555,N_7372,N_7366);
and U7556 (N_7556,N_7210,N_7486);
nor U7557 (N_7557,N_7293,N_7436);
nor U7558 (N_7558,N_7307,N_7286);
xor U7559 (N_7559,N_7281,N_7271);
or U7560 (N_7560,N_7473,N_7255);
or U7561 (N_7561,N_7339,N_7464);
or U7562 (N_7562,N_7431,N_7382);
nor U7563 (N_7563,N_7280,N_7439);
xor U7564 (N_7564,N_7374,N_7367);
xor U7565 (N_7565,N_7267,N_7288);
and U7566 (N_7566,N_7406,N_7211);
or U7567 (N_7567,N_7244,N_7483);
nand U7568 (N_7568,N_7330,N_7201);
or U7569 (N_7569,N_7226,N_7296);
xnor U7570 (N_7570,N_7237,N_7442);
xor U7571 (N_7571,N_7443,N_7410);
nand U7572 (N_7572,N_7491,N_7306);
and U7573 (N_7573,N_7467,N_7229);
xor U7574 (N_7574,N_7300,N_7219);
and U7575 (N_7575,N_7395,N_7430);
nor U7576 (N_7576,N_7320,N_7456);
or U7577 (N_7577,N_7214,N_7234);
or U7578 (N_7578,N_7477,N_7261);
nand U7579 (N_7579,N_7401,N_7449);
and U7580 (N_7580,N_7247,N_7216);
xor U7581 (N_7581,N_7379,N_7453);
or U7582 (N_7582,N_7290,N_7409);
xnor U7583 (N_7583,N_7205,N_7318);
or U7584 (N_7584,N_7263,N_7340);
and U7585 (N_7585,N_7305,N_7496);
xor U7586 (N_7586,N_7435,N_7387);
xnor U7587 (N_7587,N_7484,N_7254);
nor U7588 (N_7588,N_7268,N_7233);
and U7589 (N_7589,N_7276,N_7347);
and U7590 (N_7590,N_7225,N_7454);
nor U7591 (N_7591,N_7350,N_7355);
nor U7592 (N_7592,N_7359,N_7437);
nand U7593 (N_7593,N_7209,N_7346);
or U7594 (N_7594,N_7360,N_7389);
nor U7595 (N_7595,N_7492,N_7302);
nor U7596 (N_7596,N_7212,N_7444);
or U7597 (N_7597,N_7240,N_7458);
xor U7598 (N_7598,N_7451,N_7363);
xor U7599 (N_7599,N_7228,N_7408);
xnor U7600 (N_7600,N_7415,N_7396);
or U7601 (N_7601,N_7203,N_7353);
nor U7602 (N_7602,N_7257,N_7298);
and U7603 (N_7603,N_7315,N_7200);
xor U7604 (N_7604,N_7393,N_7407);
and U7605 (N_7605,N_7202,N_7386);
nand U7606 (N_7606,N_7217,N_7220);
or U7607 (N_7607,N_7328,N_7335);
xor U7608 (N_7608,N_7289,N_7207);
xnor U7609 (N_7609,N_7381,N_7213);
nand U7610 (N_7610,N_7287,N_7251);
xor U7611 (N_7611,N_7463,N_7308);
nand U7612 (N_7612,N_7414,N_7365);
or U7613 (N_7613,N_7204,N_7295);
xnor U7614 (N_7614,N_7329,N_7447);
and U7615 (N_7615,N_7403,N_7385);
or U7616 (N_7616,N_7394,N_7278);
nand U7617 (N_7617,N_7441,N_7446);
nor U7618 (N_7618,N_7304,N_7313);
nor U7619 (N_7619,N_7321,N_7218);
and U7620 (N_7620,N_7370,N_7316);
or U7621 (N_7621,N_7351,N_7243);
nand U7622 (N_7622,N_7397,N_7323);
and U7623 (N_7623,N_7480,N_7417);
nor U7624 (N_7624,N_7338,N_7246);
and U7625 (N_7625,N_7362,N_7275);
nand U7626 (N_7626,N_7445,N_7332);
or U7627 (N_7627,N_7476,N_7223);
xor U7628 (N_7628,N_7427,N_7361);
nor U7629 (N_7629,N_7429,N_7462);
nor U7630 (N_7630,N_7252,N_7377);
nor U7631 (N_7631,N_7264,N_7331);
and U7632 (N_7632,N_7434,N_7248);
nand U7633 (N_7633,N_7224,N_7241);
nand U7634 (N_7634,N_7424,N_7311);
nor U7635 (N_7635,N_7259,N_7250);
or U7636 (N_7636,N_7475,N_7420);
xor U7637 (N_7637,N_7215,N_7498);
nor U7638 (N_7638,N_7258,N_7310);
xnor U7639 (N_7639,N_7461,N_7388);
and U7640 (N_7640,N_7334,N_7253);
and U7641 (N_7641,N_7285,N_7266);
nand U7642 (N_7642,N_7474,N_7419);
or U7643 (N_7643,N_7333,N_7413);
or U7644 (N_7644,N_7378,N_7472);
nand U7645 (N_7645,N_7294,N_7482);
nor U7646 (N_7646,N_7345,N_7282);
nor U7647 (N_7647,N_7421,N_7466);
or U7648 (N_7648,N_7457,N_7495);
or U7649 (N_7649,N_7343,N_7283);
or U7650 (N_7650,N_7477,N_7254);
or U7651 (N_7651,N_7346,N_7464);
nand U7652 (N_7652,N_7247,N_7461);
xnor U7653 (N_7653,N_7242,N_7273);
xor U7654 (N_7654,N_7464,N_7328);
xnor U7655 (N_7655,N_7239,N_7230);
and U7656 (N_7656,N_7469,N_7353);
xor U7657 (N_7657,N_7259,N_7405);
xnor U7658 (N_7658,N_7338,N_7255);
and U7659 (N_7659,N_7421,N_7402);
and U7660 (N_7660,N_7298,N_7234);
xnor U7661 (N_7661,N_7391,N_7358);
nor U7662 (N_7662,N_7256,N_7231);
nand U7663 (N_7663,N_7250,N_7294);
nor U7664 (N_7664,N_7441,N_7400);
and U7665 (N_7665,N_7414,N_7324);
nand U7666 (N_7666,N_7316,N_7281);
and U7667 (N_7667,N_7495,N_7267);
xor U7668 (N_7668,N_7323,N_7227);
and U7669 (N_7669,N_7318,N_7455);
and U7670 (N_7670,N_7425,N_7247);
nand U7671 (N_7671,N_7372,N_7386);
nand U7672 (N_7672,N_7236,N_7345);
nor U7673 (N_7673,N_7461,N_7234);
nand U7674 (N_7674,N_7209,N_7311);
xor U7675 (N_7675,N_7401,N_7417);
nor U7676 (N_7676,N_7208,N_7313);
nand U7677 (N_7677,N_7467,N_7357);
and U7678 (N_7678,N_7292,N_7374);
xor U7679 (N_7679,N_7422,N_7362);
nor U7680 (N_7680,N_7242,N_7327);
nor U7681 (N_7681,N_7392,N_7245);
nor U7682 (N_7682,N_7335,N_7272);
nand U7683 (N_7683,N_7344,N_7355);
or U7684 (N_7684,N_7468,N_7260);
and U7685 (N_7685,N_7468,N_7252);
nand U7686 (N_7686,N_7237,N_7386);
and U7687 (N_7687,N_7473,N_7283);
or U7688 (N_7688,N_7326,N_7344);
and U7689 (N_7689,N_7304,N_7210);
and U7690 (N_7690,N_7331,N_7412);
xor U7691 (N_7691,N_7410,N_7438);
nand U7692 (N_7692,N_7382,N_7292);
or U7693 (N_7693,N_7454,N_7258);
nor U7694 (N_7694,N_7434,N_7224);
or U7695 (N_7695,N_7318,N_7350);
nand U7696 (N_7696,N_7243,N_7450);
and U7697 (N_7697,N_7353,N_7391);
nor U7698 (N_7698,N_7336,N_7247);
or U7699 (N_7699,N_7486,N_7329);
nor U7700 (N_7700,N_7256,N_7353);
nand U7701 (N_7701,N_7385,N_7460);
or U7702 (N_7702,N_7353,N_7386);
or U7703 (N_7703,N_7471,N_7319);
or U7704 (N_7704,N_7305,N_7360);
or U7705 (N_7705,N_7384,N_7480);
nand U7706 (N_7706,N_7428,N_7246);
nor U7707 (N_7707,N_7455,N_7294);
xor U7708 (N_7708,N_7381,N_7228);
nand U7709 (N_7709,N_7213,N_7321);
xor U7710 (N_7710,N_7384,N_7348);
and U7711 (N_7711,N_7417,N_7264);
or U7712 (N_7712,N_7453,N_7272);
and U7713 (N_7713,N_7411,N_7443);
nor U7714 (N_7714,N_7400,N_7226);
xor U7715 (N_7715,N_7491,N_7224);
nand U7716 (N_7716,N_7413,N_7415);
nand U7717 (N_7717,N_7355,N_7441);
nand U7718 (N_7718,N_7399,N_7378);
nand U7719 (N_7719,N_7498,N_7257);
nand U7720 (N_7720,N_7326,N_7346);
nand U7721 (N_7721,N_7454,N_7213);
nand U7722 (N_7722,N_7341,N_7226);
or U7723 (N_7723,N_7342,N_7459);
or U7724 (N_7724,N_7440,N_7490);
nand U7725 (N_7725,N_7383,N_7283);
xor U7726 (N_7726,N_7287,N_7329);
and U7727 (N_7727,N_7471,N_7341);
and U7728 (N_7728,N_7398,N_7303);
and U7729 (N_7729,N_7463,N_7357);
and U7730 (N_7730,N_7326,N_7457);
nor U7731 (N_7731,N_7280,N_7335);
or U7732 (N_7732,N_7461,N_7365);
or U7733 (N_7733,N_7431,N_7310);
and U7734 (N_7734,N_7342,N_7240);
and U7735 (N_7735,N_7483,N_7208);
nor U7736 (N_7736,N_7420,N_7302);
nand U7737 (N_7737,N_7345,N_7284);
nand U7738 (N_7738,N_7229,N_7384);
and U7739 (N_7739,N_7474,N_7471);
or U7740 (N_7740,N_7452,N_7344);
and U7741 (N_7741,N_7356,N_7464);
xnor U7742 (N_7742,N_7465,N_7453);
and U7743 (N_7743,N_7459,N_7431);
and U7744 (N_7744,N_7437,N_7232);
or U7745 (N_7745,N_7286,N_7481);
nor U7746 (N_7746,N_7472,N_7316);
or U7747 (N_7747,N_7226,N_7217);
nand U7748 (N_7748,N_7325,N_7373);
nor U7749 (N_7749,N_7435,N_7412);
nand U7750 (N_7750,N_7357,N_7266);
and U7751 (N_7751,N_7427,N_7367);
and U7752 (N_7752,N_7337,N_7427);
or U7753 (N_7753,N_7306,N_7278);
nor U7754 (N_7754,N_7480,N_7303);
nor U7755 (N_7755,N_7281,N_7368);
and U7756 (N_7756,N_7282,N_7467);
or U7757 (N_7757,N_7386,N_7407);
or U7758 (N_7758,N_7321,N_7230);
xnor U7759 (N_7759,N_7397,N_7398);
and U7760 (N_7760,N_7253,N_7263);
xnor U7761 (N_7761,N_7442,N_7308);
xnor U7762 (N_7762,N_7387,N_7491);
or U7763 (N_7763,N_7464,N_7347);
nand U7764 (N_7764,N_7471,N_7455);
nor U7765 (N_7765,N_7403,N_7451);
or U7766 (N_7766,N_7262,N_7398);
or U7767 (N_7767,N_7343,N_7342);
nand U7768 (N_7768,N_7271,N_7453);
xnor U7769 (N_7769,N_7310,N_7355);
or U7770 (N_7770,N_7392,N_7280);
xnor U7771 (N_7771,N_7409,N_7388);
nand U7772 (N_7772,N_7312,N_7231);
and U7773 (N_7773,N_7492,N_7375);
nand U7774 (N_7774,N_7364,N_7201);
xnor U7775 (N_7775,N_7462,N_7276);
and U7776 (N_7776,N_7314,N_7469);
and U7777 (N_7777,N_7406,N_7226);
nand U7778 (N_7778,N_7231,N_7420);
nor U7779 (N_7779,N_7420,N_7222);
or U7780 (N_7780,N_7361,N_7291);
and U7781 (N_7781,N_7427,N_7275);
nor U7782 (N_7782,N_7288,N_7381);
xnor U7783 (N_7783,N_7431,N_7395);
nor U7784 (N_7784,N_7462,N_7407);
nand U7785 (N_7785,N_7337,N_7290);
or U7786 (N_7786,N_7449,N_7337);
nand U7787 (N_7787,N_7385,N_7317);
or U7788 (N_7788,N_7426,N_7460);
nor U7789 (N_7789,N_7303,N_7352);
nor U7790 (N_7790,N_7240,N_7413);
xnor U7791 (N_7791,N_7494,N_7218);
nand U7792 (N_7792,N_7266,N_7389);
or U7793 (N_7793,N_7291,N_7227);
or U7794 (N_7794,N_7350,N_7429);
nand U7795 (N_7795,N_7455,N_7396);
or U7796 (N_7796,N_7245,N_7360);
nand U7797 (N_7797,N_7309,N_7457);
xnor U7798 (N_7798,N_7286,N_7220);
xnor U7799 (N_7799,N_7468,N_7296);
and U7800 (N_7800,N_7681,N_7669);
xor U7801 (N_7801,N_7513,N_7764);
nand U7802 (N_7802,N_7683,N_7742);
or U7803 (N_7803,N_7697,N_7791);
xor U7804 (N_7804,N_7627,N_7675);
xnor U7805 (N_7805,N_7540,N_7708);
and U7806 (N_7806,N_7636,N_7704);
or U7807 (N_7807,N_7759,N_7528);
nor U7808 (N_7808,N_7637,N_7797);
xor U7809 (N_7809,N_7617,N_7628);
nor U7810 (N_7810,N_7502,N_7721);
and U7811 (N_7811,N_7756,N_7747);
and U7812 (N_7812,N_7700,N_7726);
or U7813 (N_7813,N_7761,N_7622);
nor U7814 (N_7814,N_7547,N_7733);
nand U7815 (N_7815,N_7505,N_7750);
or U7816 (N_7816,N_7736,N_7525);
xnor U7817 (N_7817,N_7664,N_7551);
nor U7818 (N_7818,N_7580,N_7757);
or U7819 (N_7819,N_7650,N_7793);
or U7820 (N_7820,N_7530,N_7666);
and U7821 (N_7821,N_7686,N_7788);
nand U7822 (N_7822,N_7725,N_7663);
and U7823 (N_7823,N_7615,N_7500);
nor U7824 (N_7824,N_7511,N_7651);
and U7825 (N_7825,N_7705,N_7732);
or U7826 (N_7826,N_7526,N_7604);
nor U7827 (N_7827,N_7515,N_7631);
xor U7828 (N_7828,N_7577,N_7644);
or U7829 (N_7829,N_7659,N_7509);
and U7830 (N_7830,N_7657,N_7755);
nand U7831 (N_7831,N_7533,N_7593);
and U7832 (N_7832,N_7519,N_7536);
or U7833 (N_7833,N_7749,N_7779);
nand U7834 (N_7834,N_7696,N_7595);
nor U7835 (N_7835,N_7699,N_7694);
or U7836 (N_7836,N_7522,N_7562);
and U7837 (N_7837,N_7751,N_7799);
xnor U7838 (N_7838,N_7527,N_7770);
nand U7839 (N_7839,N_7620,N_7692);
nand U7840 (N_7840,N_7569,N_7711);
xnor U7841 (N_7841,N_7744,N_7717);
and U7842 (N_7842,N_7701,N_7618);
or U7843 (N_7843,N_7714,N_7662);
nor U7844 (N_7844,N_7762,N_7576);
and U7845 (N_7845,N_7611,N_7677);
xnor U7846 (N_7846,N_7671,N_7518);
xnor U7847 (N_7847,N_7695,N_7643);
nand U7848 (N_7848,N_7575,N_7646);
nand U7849 (N_7849,N_7592,N_7703);
xnor U7850 (N_7850,N_7767,N_7790);
and U7851 (N_7851,N_7534,N_7786);
xnor U7852 (N_7852,N_7605,N_7738);
or U7853 (N_7853,N_7652,N_7782);
or U7854 (N_7854,N_7794,N_7648);
nor U7855 (N_7855,N_7710,N_7709);
and U7856 (N_7856,N_7514,N_7579);
nor U7857 (N_7857,N_7586,N_7630);
xnor U7858 (N_7858,N_7680,N_7792);
nand U7859 (N_7859,N_7563,N_7546);
and U7860 (N_7860,N_7568,N_7501);
xnor U7861 (N_7861,N_7587,N_7521);
and U7862 (N_7862,N_7538,N_7582);
nand U7863 (N_7863,N_7512,N_7523);
nand U7864 (N_7864,N_7689,N_7589);
xnor U7865 (N_7865,N_7691,N_7578);
or U7866 (N_7866,N_7544,N_7787);
or U7867 (N_7867,N_7581,N_7775);
xor U7868 (N_7868,N_7517,N_7571);
xor U7869 (N_7869,N_7690,N_7789);
nand U7870 (N_7870,N_7784,N_7549);
or U7871 (N_7871,N_7539,N_7625);
nor U7872 (N_7872,N_7723,N_7613);
nand U7873 (N_7873,N_7655,N_7573);
nand U7874 (N_7874,N_7504,N_7785);
and U7875 (N_7875,N_7753,N_7554);
and U7876 (N_7876,N_7591,N_7745);
nor U7877 (N_7877,N_7621,N_7614);
nor U7878 (N_7878,N_7629,N_7719);
xor U7879 (N_7879,N_7735,N_7559);
nand U7880 (N_7880,N_7772,N_7552);
nor U7881 (N_7881,N_7550,N_7640);
nand U7882 (N_7882,N_7653,N_7673);
or U7883 (N_7883,N_7558,N_7682);
nor U7884 (N_7884,N_7545,N_7771);
and U7885 (N_7885,N_7722,N_7707);
and U7886 (N_7886,N_7769,N_7510);
nand U7887 (N_7887,N_7555,N_7678);
nor U7888 (N_7888,N_7556,N_7503);
nand U7889 (N_7889,N_7602,N_7565);
nand U7890 (N_7890,N_7642,N_7760);
nor U7891 (N_7891,N_7773,N_7780);
nand U7892 (N_7892,N_7574,N_7674);
or U7893 (N_7893,N_7766,N_7619);
or U7894 (N_7894,N_7609,N_7668);
or U7895 (N_7895,N_7715,N_7672);
nor U7896 (N_7896,N_7743,N_7740);
xor U7897 (N_7897,N_7601,N_7507);
nor U7898 (N_7898,N_7720,N_7516);
xor U7899 (N_7899,N_7553,N_7597);
xor U7900 (N_7900,N_7566,N_7713);
xnor U7901 (N_7901,N_7665,N_7783);
and U7902 (N_7902,N_7638,N_7684);
nor U7903 (N_7903,N_7739,N_7693);
or U7904 (N_7904,N_7603,N_7583);
xor U7905 (N_7905,N_7647,N_7541);
nor U7906 (N_7906,N_7535,N_7660);
and U7907 (N_7907,N_7746,N_7520);
xnor U7908 (N_7908,N_7765,N_7676);
and U7909 (N_7909,N_7670,N_7531);
or U7910 (N_7910,N_7798,N_7658);
nand U7911 (N_7911,N_7537,N_7634);
nor U7912 (N_7912,N_7560,N_7641);
and U7913 (N_7913,N_7612,N_7570);
or U7914 (N_7914,N_7716,N_7564);
xor U7915 (N_7915,N_7698,N_7633);
and U7916 (N_7916,N_7758,N_7584);
nor U7917 (N_7917,N_7754,N_7763);
nand U7918 (N_7918,N_7508,N_7632);
xnor U7919 (N_7919,N_7532,N_7688);
and U7920 (N_7920,N_7781,N_7585);
nor U7921 (N_7921,N_7623,N_7654);
xnor U7922 (N_7922,N_7731,N_7561);
nand U7923 (N_7923,N_7626,N_7778);
nor U7924 (N_7924,N_7795,N_7685);
or U7925 (N_7925,N_7667,N_7661);
and U7926 (N_7926,N_7702,N_7567);
nand U7927 (N_7927,N_7712,N_7728);
nor U7928 (N_7928,N_7542,N_7706);
nand U7929 (N_7929,N_7776,N_7748);
xnor U7930 (N_7930,N_7752,N_7606);
xor U7931 (N_7931,N_7529,N_7741);
and U7932 (N_7932,N_7506,N_7645);
xnor U7933 (N_7933,N_7656,N_7572);
and U7934 (N_7934,N_7639,N_7590);
nand U7935 (N_7935,N_7616,N_7594);
nor U7936 (N_7936,N_7524,N_7796);
and U7937 (N_7937,N_7727,N_7635);
and U7938 (N_7938,N_7598,N_7724);
xnor U7939 (N_7939,N_7718,N_7588);
xor U7940 (N_7940,N_7624,N_7687);
nor U7941 (N_7941,N_7543,N_7768);
nor U7942 (N_7942,N_7548,N_7610);
xor U7943 (N_7943,N_7729,N_7774);
or U7944 (N_7944,N_7599,N_7596);
or U7945 (N_7945,N_7557,N_7730);
nor U7946 (N_7946,N_7607,N_7649);
or U7947 (N_7947,N_7679,N_7734);
and U7948 (N_7948,N_7608,N_7777);
xnor U7949 (N_7949,N_7737,N_7600);
and U7950 (N_7950,N_7516,N_7575);
nor U7951 (N_7951,N_7770,N_7632);
xor U7952 (N_7952,N_7613,N_7538);
or U7953 (N_7953,N_7685,N_7738);
nand U7954 (N_7954,N_7620,N_7587);
or U7955 (N_7955,N_7627,N_7585);
xor U7956 (N_7956,N_7787,N_7792);
xnor U7957 (N_7957,N_7584,N_7676);
or U7958 (N_7958,N_7782,N_7555);
xnor U7959 (N_7959,N_7637,N_7522);
or U7960 (N_7960,N_7630,N_7675);
nor U7961 (N_7961,N_7615,N_7646);
and U7962 (N_7962,N_7776,N_7525);
nand U7963 (N_7963,N_7590,N_7557);
nand U7964 (N_7964,N_7599,N_7610);
and U7965 (N_7965,N_7646,N_7644);
xnor U7966 (N_7966,N_7557,N_7541);
or U7967 (N_7967,N_7576,N_7732);
or U7968 (N_7968,N_7568,N_7508);
nor U7969 (N_7969,N_7598,N_7528);
and U7970 (N_7970,N_7634,N_7716);
or U7971 (N_7971,N_7585,N_7666);
nor U7972 (N_7972,N_7695,N_7601);
nor U7973 (N_7973,N_7566,N_7687);
and U7974 (N_7974,N_7606,N_7608);
or U7975 (N_7975,N_7725,N_7690);
nor U7976 (N_7976,N_7792,N_7775);
and U7977 (N_7977,N_7649,N_7537);
nand U7978 (N_7978,N_7516,N_7602);
nand U7979 (N_7979,N_7676,N_7731);
nor U7980 (N_7980,N_7502,N_7628);
or U7981 (N_7981,N_7566,N_7759);
xor U7982 (N_7982,N_7561,N_7683);
or U7983 (N_7983,N_7697,N_7529);
nor U7984 (N_7984,N_7579,N_7518);
nor U7985 (N_7985,N_7686,N_7786);
or U7986 (N_7986,N_7740,N_7637);
xor U7987 (N_7987,N_7765,N_7674);
xnor U7988 (N_7988,N_7640,N_7642);
or U7989 (N_7989,N_7552,N_7660);
nor U7990 (N_7990,N_7671,N_7545);
xor U7991 (N_7991,N_7631,N_7786);
and U7992 (N_7992,N_7646,N_7596);
and U7993 (N_7993,N_7699,N_7781);
or U7994 (N_7994,N_7531,N_7745);
or U7995 (N_7995,N_7719,N_7750);
nand U7996 (N_7996,N_7604,N_7733);
xor U7997 (N_7997,N_7776,N_7569);
or U7998 (N_7998,N_7537,N_7695);
nor U7999 (N_7999,N_7576,N_7759);
xnor U8000 (N_8000,N_7535,N_7772);
or U8001 (N_8001,N_7758,N_7717);
or U8002 (N_8002,N_7678,N_7521);
or U8003 (N_8003,N_7775,N_7557);
nand U8004 (N_8004,N_7663,N_7695);
xnor U8005 (N_8005,N_7791,N_7575);
or U8006 (N_8006,N_7520,N_7601);
and U8007 (N_8007,N_7675,N_7744);
nand U8008 (N_8008,N_7741,N_7587);
and U8009 (N_8009,N_7678,N_7784);
nand U8010 (N_8010,N_7559,N_7517);
nand U8011 (N_8011,N_7629,N_7576);
nand U8012 (N_8012,N_7562,N_7605);
or U8013 (N_8013,N_7627,N_7731);
xor U8014 (N_8014,N_7534,N_7606);
nand U8015 (N_8015,N_7743,N_7654);
xnor U8016 (N_8016,N_7534,N_7608);
xnor U8017 (N_8017,N_7626,N_7550);
and U8018 (N_8018,N_7608,N_7744);
nand U8019 (N_8019,N_7640,N_7721);
or U8020 (N_8020,N_7580,N_7522);
and U8021 (N_8021,N_7515,N_7637);
nor U8022 (N_8022,N_7792,N_7659);
nor U8023 (N_8023,N_7766,N_7719);
or U8024 (N_8024,N_7507,N_7566);
nand U8025 (N_8025,N_7579,N_7749);
xnor U8026 (N_8026,N_7674,N_7516);
nand U8027 (N_8027,N_7752,N_7713);
nand U8028 (N_8028,N_7714,N_7756);
nor U8029 (N_8029,N_7634,N_7554);
nor U8030 (N_8030,N_7572,N_7631);
and U8031 (N_8031,N_7736,N_7738);
and U8032 (N_8032,N_7532,N_7671);
nand U8033 (N_8033,N_7625,N_7637);
or U8034 (N_8034,N_7796,N_7741);
and U8035 (N_8035,N_7790,N_7769);
xnor U8036 (N_8036,N_7673,N_7644);
nor U8037 (N_8037,N_7648,N_7567);
nand U8038 (N_8038,N_7590,N_7696);
xnor U8039 (N_8039,N_7696,N_7752);
and U8040 (N_8040,N_7677,N_7533);
or U8041 (N_8041,N_7614,N_7623);
or U8042 (N_8042,N_7754,N_7641);
nor U8043 (N_8043,N_7728,N_7549);
xnor U8044 (N_8044,N_7655,N_7657);
nand U8045 (N_8045,N_7534,N_7552);
nand U8046 (N_8046,N_7589,N_7790);
and U8047 (N_8047,N_7614,N_7685);
nand U8048 (N_8048,N_7537,N_7619);
or U8049 (N_8049,N_7623,N_7767);
nand U8050 (N_8050,N_7583,N_7670);
nor U8051 (N_8051,N_7691,N_7777);
and U8052 (N_8052,N_7553,N_7564);
or U8053 (N_8053,N_7677,N_7768);
nand U8054 (N_8054,N_7766,N_7635);
and U8055 (N_8055,N_7721,N_7651);
xor U8056 (N_8056,N_7537,N_7755);
or U8057 (N_8057,N_7591,N_7664);
nand U8058 (N_8058,N_7739,N_7687);
or U8059 (N_8059,N_7527,N_7535);
xnor U8060 (N_8060,N_7583,N_7732);
nor U8061 (N_8061,N_7508,N_7729);
nor U8062 (N_8062,N_7708,N_7617);
and U8063 (N_8063,N_7697,N_7724);
nor U8064 (N_8064,N_7757,N_7602);
and U8065 (N_8065,N_7769,N_7627);
nor U8066 (N_8066,N_7649,N_7687);
or U8067 (N_8067,N_7646,N_7551);
nor U8068 (N_8068,N_7573,N_7671);
nor U8069 (N_8069,N_7791,N_7618);
xor U8070 (N_8070,N_7677,N_7729);
nand U8071 (N_8071,N_7631,N_7605);
nor U8072 (N_8072,N_7588,N_7692);
and U8073 (N_8073,N_7763,N_7741);
nand U8074 (N_8074,N_7759,N_7639);
xnor U8075 (N_8075,N_7523,N_7631);
nand U8076 (N_8076,N_7757,N_7735);
nor U8077 (N_8077,N_7685,N_7545);
nor U8078 (N_8078,N_7775,N_7543);
or U8079 (N_8079,N_7561,N_7583);
nand U8080 (N_8080,N_7586,N_7704);
nand U8081 (N_8081,N_7594,N_7734);
or U8082 (N_8082,N_7778,N_7755);
and U8083 (N_8083,N_7777,N_7542);
nand U8084 (N_8084,N_7687,N_7510);
and U8085 (N_8085,N_7793,N_7584);
or U8086 (N_8086,N_7531,N_7638);
and U8087 (N_8087,N_7506,N_7759);
xnor U8088 (N_8088,N_7732,N_7508);
nand U8089 (N_8089,N_7541,N_7590);
or U8090 (N_8090,N_7689,N_7734);
nand U8091 (N_8091,N_7630,N_7745);
nor U8092 (N_8092,N_7549,N_7570);
xnor U8093 (N_8093,N_7535,N_7723);
nor U8094 (N_8094,N_7677,N_7624);
nand U8095 (N_8095,N_7542,N_7601);
xnor U8096 (N_8096,N_7505,N_7717);
nand U8097 (N_8097,N_7714,N_7631);
xnor U8098 (N_8098,N_7728,N_7627);
nand U8099 (N_8099,N_7558,N_7753);
and U8100 (N_8100,N_7817,N_8003);
and U8101 (N_8101,N_8018,N_8041);
nor U8102 (N_8102,N_7911,N_7931);
and U8103 (N_8103,N_7903,N_7842);
nand U8104 (N_8104,N_7997,N_8068);
or U8105 (N_8105,N_7833,N_8030);
and U8106 (N_8106,N_7802,N_7875);
or U8107 (N_8107,N_7916,N_8097);
or U8108 (N_8108,N_7999,N_7941);
nor U8109 (N_8109,N_8020,N_7990);
nand U8110 (N_8110,N_7900,N_8066);
nand U8111 (N_8111,N_7850,N_7813);
or U8112 (N_8112,N_7882,N_7947);
nand U8113 (N_8113,N_7945,N_8059);
and U8114 (N_8114,N_7840,N_7811);
xnor U8115 (N_8115,N_7878,N_7991);
xnor U8116 (N_8116,N_7958,N_7907);
xnor U8117 (N_8117,N_7898,N_7905);
nor U8118 (N_8118,N_7950,N_7843);
nand U8119 (N_8119,N_7922,N_8058);
nor U8120 (N_8120,N_7979,N_8096);
and U8121 (N_8121,N_7956,N_7890);
or U8122 (N_8122,N_8025,N_7927);
nand U8123 (N_8123,N_7888,N_7928);
or U8124 (N_8124,N_7880,N_8094);
or U8125 (N_8125,N_7835,N_7913);
and U8126 (N_8126,N_7870,N_7884);
xnor U8127 (N_8127,N_7822,N_7868);
or U8128 (N_8128,N_7883,N_7845);
or U8129 (N_8129,N_7964,N_8010);
or U8130 (N_8130,N_7871,N_8019);
or U8131 (N_8131,N_7946,N_7937);
or U8132 (N_8132,N_7820,N_8065);
nor U8133 (N_8133,N_8044,N_7984);
and U8134 (N_8134,N_8090,N_8039);
or U8135 (N_8135,N_7978,N_7961);
xor U8136 (N_8136,N_8022,N_7825);
nor U8137 (N_8137,N_7861,N_7877);
nand U8138 (N_8138,N_7851,N_7926);
xor U8139 (N_8139,N_7887,N_7803);
nor U8140 (N_8140,N_7943,N_8040);
nand U8141 (N_8141,N_7954,N_7998);
and U8142 (N_8142,N_7976,N_7806);
or U8143 (N_8143,N_8038,N_7992);
and U8144 (N_8144,N_7853,N_8055);
xor U8145 (N_8145,N_8075,N_7908);
xnor U8146 (N_8146,N_8083,N_7929);
xnor U8147 (N_8147,N_7989,N_7818);
nor U8148 (N_8148,N_8057,N_8052);
or U8149 (N_8149,N_7988,N_7859);
nor U8150 (N_8150,N_7860,N_7801);
nand U8151 (N_8151,N_7986,N_8054);
nor U8152 (N_8152,N_7968,N_7856);
nor U8153 (N_8153,N_7971,N_7969);
nand U8154 (N_8154,N_7891,N_8079);
xor U8155 (N_8155,N_8067,N_7899);
or U8156 (N_8156,N_7932,N_8036);
and U8157 (N_8157,N_7930,N_7854);
xor U8158 (N_8158,N_7821,N_7841);
xor U8159 (N_8159,N_7959,N_7920);
or U8160 (N_8160,N_7844,N_7893);
or U8161 (N_8161,N_8032,N_7938);
nor U8162 (N_8162,N_7919,N_7885);
or U8163 (N_8163,N_8043,N_8017);
nor U8164 (N_8164,N_8015,N_8001);
and U8165 (N_8165,N_7995,N_7879);
or U8166 (N_8166,N_8069,N_7852);
nor U8167 (N_8167,N_7894,N_8006);
or U8168 (N_8168,N_7948,N_7977);
xnor U8169 (N_8169,N_7804,N_8063);
nand U8170 (N_8170,N_8081,N_7914);
nor U8171 (N_8171,N_8086,N_7872);
xnor U8172 (N_8172,N_8080,N_7963);
xor U8173 (N_8173,N_8095,N_7962);
xnor U8174 (N_8174,N_7909,N_7970);
xnor U8175 (N_8175,N_7829,N_8046);
or U8176 (N_8176,N_7924,N_8061);
xor U8177 (N_8177,N_7966,N_8007);
and U8178 (N_8178,N_7994,N_8026);
xnor U8179 (N_8179,N_7892,N_8076);
and U8180 (N_8180,N_7967,N_8028);
xnor U8181 (N_8181,N_8029,N_7925);
xnor U8182 (N_8182,N_8023,N_7855);
nand U8183 (N_8183,N_7944,N_8048);
nor U8184 (N_8184,N_8073,N_7873);
xnor U8185 (N_8185,N_8070,N_8060);
nand U8186 (N_8186,N_7936,N_8089);
nand U8187 (N_8187,N_7831,N_7912);
xnor U8188 (N_8188,N_8035,N_8031);
nor U8189 (N_8189,N_7996,N_8027);
xor U8190 (N_8190,N_7917,N_7939);
nand U8191 (N_8191,N_8011,N_7808);
nor U8192 (N_8192,N_7933,N_7823);
xnor U8193 (N_8193,N_7866,N_7858);
and U8194 (N_8194,N_7923,N_8005);
nand U8195 (N_8195,N_8078,N_7857);
nor U8196 (N_8196,N_7874,N_8084);
or U8197 (N_8197,N_7983,N_7934);
xnor U8198 (N_8198,N_7921,N_8049);
or U8199 (N_8199,N_8004,N_8037);
nand U8200 (N_8200,N_8008,N_7869);
nor U8201 (N_8201,N_7824,N_7864);
and U8202 (N_8202,N_8053,N_7815);
nor U8203 (N_8203,N_8056,N_7863);
nand U8204 (N_8204,N_8085,N_7904);
or U8205 (N_8205,N_7942,N_8093);
and U8206 (N_8206,N_7838,N_7940);
nor U8207 (N_8207,N_7980,N_7993);
nand U8208 (N_8208,N_8077,N_7816);
nand U8209 (N_8209,N_7965,N_7830);
nand U8210 (N_8210,N_8000,N_8099);
and U8211 (N_8211,N_7827,N_8012);
and U8212 (N_8212,N_8045,N_7881);
or U8213 (N_8213,N_7867,N_8047);
or U8214 (N_8214,N_7832,N_8062);
xnor U8215 (N_8215,N_8050,N_8092);
nor U8216 (N_8216,N_8082,N_8021);
xnor U8217 (N_8217,N_7951,N_7819);
nand U8218 (N_8218,N_7975,N_7836);
or U8219 (N_8219,N_8087,N_7849);
and U8220 (N_8220,N_7876,N_7805);
xor U8221 (N_8221,N_7837,N_7897);
nor U8222 (N_8222,N_8088,N_8098);
nor U8223 (N_8223,N_8009,N_7865);
nor U8224 (N_8224,N_7826,N_7910);
nand U8225 (N_8225,N_7952,N_7960);
and U8226 (N_8226,N_8071,N_7834);
nor U8227 (N_8227,N_8013,N_7906);
nand U8228 (N_8228,N_7800,N_8002);
and U8229 (N_8229,N_8064,N_7902);
xor U8230 (N_8230,N_7955,N_7982);
xnor U8231 (N_8231,N_7828,N_8014);
and U8232 (N_8232,N_7896,N_7889);
nand U8233 (N_8233,N_7949,N_7809);
nand U8234 (N_8234,N_7953,N_7972);
nor U8235 (N_8235,N_8042,N_7812);
or U8236 (N_8236,N_7814,N_7973);
nand U8237 (N_8237,N_7957,N_7839);
or U8238 (N_8238,N_7810,N_7915);
and U8239 (N_8239,N_7974,N_8024);
and U8240 (N_8240,N_7981,N_7918);
nand U8241 (N_8241,N_7807,N_8072);
or U8242 (N_8242,N_7847,N_7846);
xnor U8243 (N_8243,N_8016,N_8091);
nor U8244 (N_8244,N_7901,N_7935);
and U8245 (N_8245,N_7886,N_8033);
or U8246 (N_8246,N_7985,N_7987);
or U8247 (N_8247,N_8034,N_7848);
nand U8248 (N_8248,N_8074,N_7862);
and U8249 (N_8249,N_8051,N_7895);
or U8250 (N_8250,N_7827,N_8056);
or U8251 (N_8251,N_8030,N_8098);
xor U8252 (N_8252,N_7881,N_7825);
and U8253 (N_8253,N_7931,N_7899);
nor U8254 (N_8254,N_7812,N_8016);
nor U8255 (N_8255,N_7875,N_8053);
or U8256 (N_8256,N_7958,N_7802);
and U8257 (N_8257,N_8048,N_7885);
nand U8258 (N_8258,N_8031,N_8042);
and U8259 (N_8259,N_7921,N_7802);
and U8260 (N_8260,N_7904,N_7977);
or U8261 (N_8261,N_7841,N_8076);
and U8262 (N_8262,N_8016,N_8033);
nor U8263 (N_8263,N_7945,N_8031);
xor U8264 (N_8264,N_7945,N_8024);
and U8265 (N_8265,N_8067,N_7959);
nor U8266 (N_8266,N_8044,N_8082);
or U8267 (N_8267,N_8071,N_8046);
nor U8268 (N_8268,N_8013,N_7998);
or U8269 (N_8269,N_7904,N_7867);
nand U8270 (N_8270,N_7807,N_7929);
nor U8271 (N_8271,N_7959,N_7879);
nand U8272 (N_8272,N_7965,N_7977);
nand U8273 (N_8273,N_7866,N_7892);
nor U8274 (N_8274,N_8050,N_7815);
xnor U8275 (N_8275,N_8047,N_7945);
nand U8276 (N_8276,N_7969,N_7893);
nor U8277 (N_8277,N_7867,N_7990);
nand U8278 (N_8278,N_8071,N_8068);
nor U8279 (N_8279,N_8039,N_8021);
or U8280 (N_8280,N_8002,N_7826);
nor U8281 (N_8281,N_8066,N_7835);
nor U8282 (N_8282,N_8087,N_7963);
nand U8283 (N_8283,N_8036,N_7807);
nor U8284 (N_8284,N_7923,N_7843);
xor U8285 (N_8285,N_7982,N_8061);
xor U8286 (N_8286,N_7950,N_8037);
nor U8287 (N_8287,N_8057,N_8070);
and U8288 (N_8288,N_8007,N_7814);
nor U8289 (N_8289,N_7947,N_7838);
and U8290 (N_8290,N_7893,N_7803);
and U8291 (N_8291,N_8023,N_8082);
xnor U8292 (N_8292,N_8051,N_7839);
and U8293 (N_8293,N_8038,N_7898);
xnor U8294 (N_8294,N_7930,N_7899);
and U8295 (N_8295,N_8014,N_7960);
nand U8296 (N_8296,N_7806,N_7955);
nand U8297 (N_8297,N_8089,N_7848);
or U8298 (N_8298,N_7946,N_7917);
xor U8299 (N_8299,N_8086,N_8038);
nand U8300 (N_8300,N_7873,N_7925);
and U8301 (N_8301,N_7911,N_7897);
nor U8302 (N_8302,N_7825,N_8017);
nand U8303 (N_8303,N_7888,N_7914);
nor U8304 (N_8304,N_7989,N_8088);
xor U8305 (N_8305,N_7937,N_7984);
xor U8306 (N_8306,N_8064,N_8022);
nand U8307 (N_8307,N_8000,N_7815);
nor U8308 (N_8308,N_8080,N_8007);
nor U8309 (N_8309,N_7933,N_8038);
and U8310 (N_8310,N_8043,N_8039);
and U8311 (N_8311,N_7951,N_7890);
xor U8312 (N_8312,N_7873,N_8078);
xor U8313 (N_8313,N_7998,N_8028);
or U8314 (N_8314,N_7916,N_7866);
xnor U8315 (N_8315,N_7949,N_7935);
or U8316 (N_8316,N_8066,N_8010);
or U8317 (N_8317,N_8006,N_7911);
or U8318 (N_8318,N_7912,N_8097);
or U8319 (N_8319,N_7910,N_8092);
or U8320 (N_8320,N_7841,N_7859);
and U8321 (N_8321,N_7840,N_7860);
nor U8322 (N_8322,N_8093,N_7919);
nor U8323 (N_8323,N_7865,N_7988);
nor U8324 (N_8324,N_7870,N_8048);
nand U8325 (N_8325,N_7891,N_7911);
xor U8326 (N_8326,N_7850,N_8007);
xnor U8327 (N_8327,N_8053,N_7913);
nor U8328 (N_8328,N_7911,N_7859);
or U8329 (N_8329,N_8058,N_7856);
xnor U8330 (N_8330,N_8012,N_7895);
xnor U8331 (N_8331,N_8072,N_8051);
and U8332 (N_8332,N_7946,N_8014);
nand U8333 (N_8333,N_7871,N_7860);
xor U8334 (N_8334,N_7992,N_8076);
xnor U8335 (N_8335,N_8049,N_7949);
and U8336 (N_8336,N_7820,N_8008);
xor U8337 (N_8337,N_7952,N_8052);
xor U8338 (N_8338,N_7983,N_8006);
or U8339 (N_8339,N_8065,N_8093);
nor U8340 (N_8340,N_8003,N_8085);
and U8341 (N_8341,N_7974,N_8019);
xnor U8342 (N_8342,N_7932,N_7931);
or U8343 (N_8343,N_7874,N_7984);
nor U8344 (N_8344,N_8033,N_7819);
nand U8345 (N_8345,N_7811,N_7981);
and U8346 (N_8346,N_7807,N_7985);
or U8347 (N_8347,N_8098,N_8026);
nor U8348 (N_8348,N_7891,N_8067);
nor U8349 (N_8349,N_8049,N_8009);
and U8350 (N_8350,N_8035,N_7854);
xnor U8351 (N_8351,N_7828,N_7822);
or U8352 (N_8352,N_7929,N_7907);
or U8353 (N_8353,N_7955,N_8087);
nor U8354 (N_8354,N_7862,N_7814);
xnor U8355 (N_8355,N_7807,N_8043);
nor U8356 (N_8356,N_7957,N_8001);
nand U8357 (N_8357,N_7869,N_7906);
nor U8358 (N_8358,N_7951,N_7900);
nor U8359 (N_8359,N_7919,N_8051);
and U8360 (N_8360,N_7946,N_7965);
or U8361 (N_8361,N_7940,N_7980);
or U8362 (N_8362,N_7897,N_8045);
or U8363 (N_8363,N_8027,N_8037);
nand U8364 (N_8364,N_8008,N_8034);
nor U8365 (N_8365,N_7802,N_8078);
nor U8366 (N_8366,N_8005,N_7909);
nor U8367 (N_8367,N_7856,N_7883);
nand U8368 (N_8368,N_7865,N_7869);
nor U8369 (N_8369,N_7807,N_7960);
or U8370 (N_8370,N_8000,N_7887);
or U8371 (N_8371,N_8009,N_7922);
nor U8372 (N_8372,N_7983,N_7810);
nand U8373 (N_8373,N_7948,N_7857);
xnor U8374 (N_8374,N_8035,N_8028);
or U8375 (N_8375,N_7881,N_8001);
nor U8376 (N_8376,N_8034,N_7949);
or U8377 (N_8377,N_8072,N_8023);
or U8378 (N_8378,N_7895,N_7916);
nand U8379 (N_8379,N_7860,N_7883);
and U8380 (N_8380,N_8082,N_8058);
and U8381 (N_8381,N_8013,N_7893);
xnor U8382 (N_8382,N_7921,N_7824);
xor U8383 (N_8383,N_7985,N_7821);
and U8384 (N_8384,N_7896,N_8011);
nand U8385 (N_8385,N_7967,N_7802);
or U8386 (N_8386,N_7946,N_8033);
nor U8387 (N_8387,N_8083,N_8042);
and U8388 (N_8388,N_7910,N_7977);
nand U8389 (N_8389,N_8098,N_7854);
or U8390 (N_8390,N_8046,N_7860);
nor U8391 (N_8391,N_8036,N_7937);
or U8392 (N_8392,N_7867,N_7821);
xor U8393 (N_8393,N_7984,N_7864);
and U8394 (N_8394,N_8073,N_7866);
and U8395 (N_8395,N_7919,N_7950);
nand U8396 (N_8396,N_8071,N_7885);
or U8397 (N_8397,N_8064,N_7809);
or U8398 (N_8398,N_7948,N_7863);
xor U8399 (N_8399,N_7977,N_7830);
or U8400 (N_8400,N_8295,N_8108);
xor U8401 (N_8401,N_8172,N_8340);
nand U8402 (N_8402,N_8345,N_8151);
nor U8403 (N_8403,N_8220,N_8190);
nand U8404 (N_8404,N_8229,N_8334);
and U8405 (N_8405,N_8223,N_8319);
nand U8406 (N_8406,N_8141,N_8337);
and U8407 (N_8407,N_8324,N_8250);
xor U8408 (N_8408,N_8361,N_8393);
xnor U8409 (N_8409,N_8242,N_8308);
and U8410 (N_8410,N_8124,N_8283);
and U8411 (N_8411,N_8188,N_8367);
and U8412 (N_8412,N_8146,N_8145);
and U8413 (N_8413,N_8318,N_8132);
nand U8414 (N_8414,N_8373,N_8320);
nor U8415 (N_8415,N_8336,N_8221);
xnor U8416 (N_8416,N_8139,N_8355);
nor U8417 (N_8417,N_8398,N_8384);
nor U8418 (N_8418,N_8115,N_8249);
nand U8419 (N_8419,N_8225,N_8125);
nand U8420 (N_8420,N_8271,N_8187);
xor U8421 (N_8421,N_8363,N_8206);
xor U8422 (N_8422,N_8230,N_8321);
nor U8423 (N_8423,N_8289,N_8153);
or U8424 (N_8424,N_8222,N_8325);
or U8425 (N_8425,N_8200,N_8241);
and U8426 (N_8426,N_8245,N_8121);
nor U8427 (N_8427,N_8300,N_8240);
nor U8428 (N_8428,N_8226,N_8148);
xor U8429 (N_8429,N_8281,N_8284);
and U8430 (N_8430,N_8117,N_8196);
or U8431 (N_8431,N_8353,N_8191);
nor U8432 (N_8432,N_8282,N_8227);
nand U8433 (N_8433,N_8143,N_8297);
nor U8434 (N_8434,N_8235,N_8365);
or U8435 (N_8435,N_8199,N_8239);
or U8436 (N_8436,N_8286,N_8105);
nor U8437 (N_8437,N_8306,N_8322);
and U8438 (N_8438,N_8182,N_8338);
nor U8439 (N_8439,N_8211,N_8328);
nor U8440 (N_8440,N_8260,N_8381);
or U8441 (N_8441,N_8195,N_8386);
xor U8442 (N_8442,N_8238,N_8327);
xor U8443 (N_8443,N_8377,N_8233);
xor U8444 (N_8444,N_8309,N_8287);
nand U8445 (N_8445,N_8290,N_8272);
nor U8446 (N_8446,N_8179,N_8301);
xor U8447 (N_8447,N_8378,N_8127);
xnor U8448 (N_8448,N_8362,N_8294);
nor U8449 (N_8449,N_8307,N_8269);
and U8450 (N_8450,N_8326,N_8280);
xor U8451 (N_8451,N_8347,N_8257);
nor U8452 (N_8452,N_8263,N_8285);
nor U8453 (N_8453,N_8293,N_8142);
nor U8454 (N_8454,N_8270,N_8312);
or U8455 (N_8455,N_8255,N_8185);
xnor U8456 (N_8456,N_8159,N_8331);
nand U8457 (N_8457,N_8277,N_8110);
and U8458 (N_8458,N_8382,N_8204);
nor U8459 (N_8459,N_8104,N_8112);
xnor U8460 (N_8460,N_8228,N_8134);
xor U8461 (N_8461,N_8164,N_8126);
nor U8462 (N_8462,N_8296,N_8354);
nand U8463 (N_8463,N_8133,N_8246);
and U8464 (N_8464,N_8383,N_8210);
nor U8465 (N_8465,N_8243,N_8155);
xnor U8466 (N_8466,N_8219,N_8166);
or U8467 (N_8467,N_8106,N_8311);
or U8468 (N_8468,N_8154,N_8313);
xor U8469 (N_8469,N_8275,N_8380);
and U8470 (N_8470,N_8276,N_8303);
or U8471 (N_8471,N_8109,N_8256);
and U8472 (N_8472,N_8129,N_8399);
and U8473 (N_8473,N_8176,N_8169);
nand U8474 (N_8474,N_8209,N_8278);
nor U8475 (N_8475,N_8379,N_8356);
nand U8476 (N_8476,N_8335,N_8150);
and U8477 (N_8477,N_8314,N_8247);
or U8478 (N_8478,N_8122,N_8123);
or U8479 (N_8479,N_8259,N_8258);
nor U8480 (N_8480,N_8273,N_8248);
and U8481 (N_8481,N_8349,N_8302);
xnor U8482 (N_8482,N_8348,N_8184);
nor U8483 (N_8483,N_8234,N_8304);
nand U8484 (N_8484,N_8152,N_8376);
and U8485 (N_8485,N_8174,N_8118);
xor U8486 (N_8486,N_8180,N_8217);
nor U8487 (N_8487,N_8279,N_8396);
nand U8488 (N_8488,N_8344,N_8252);
or U8489 (N_8489,N_8103,N_8391);
and U8490 (N_8490,N_8385,N_8343);
nand U8491 (N_8491,N_8147,N_8102);
xor U8492 (N_8492,N_8114,N_8157);
xnor U8493 (N_8493,N_8310,N_8203);
xnor U8494 (N_8494,N_8161,N_8137);
nor U8495 (N_8495,N_8168,N_8130);
and U8496 (N_8496,N_8298,N_8333);
or U8497 (N_8497,N_8330,N_8205);
nand U8498 (N_8498,N_8237,N_8254);
nor U8499 (N_8499,N_8352,N_8372);
or U8500 (N_8500,N_8107,N_8170);
or U8501 (N_8501,N_8357,N_8236);
and U8502 (N_8502,N_8389,N_8315);
or U8503 (N_8503,N_8197,N_8135);
or U8504 (N_8504,N_8186,N_8216);
xor U8505 (N_8505,N_8138,N_8156);
and U8506 (N_8506,N_8368,N_8369);
nor U8507 (N_8507,N_8232,N_8251);
nand U8508 (N_8508,N_8264,N_8339);
nand U8509 (N_8509,N_8371,N_8394);
nor U8510 (N_8510,N_8111,N_8201);
xor U8511 (N_8511,N_8291,N_8202);
nor U8512 (N_8512,N_8208,N_8167);
nand U8513 (N_8513,N_8288,N_8136);
nor U8514 (N_8514,N_8267,N_8342);
nand U8515 (N_8515,N_8265,N_8224);
xor U8516 (N_8516,N_8128,N_8218);
nand U8517 (N_8517,N_8194,N_8198);
xor U8518 (N_8518,N_8171,N_8329);
nor U8519 (N_8519,N_8351,N_8317);
nand U8520 (N_8520,N_8158,N_8163);
nor U8521 (N_8521,N_8100,N_8116);
and U8522 (N_8522,N_8212,N_8370);
xor U8523 (N_8523,N_8305,N_8192);
nor U8524 (N_8524,N_8215,N_8323);
nor U8525 (N_8525,N_8341,N_8316);
or U8526 (N_8526,N_8261,N_8165);
xnor U8527 (N_8527,N_8193,N_8231);
nand U8528 (N_8528,N_8144,N_8395);
nor U8529 (N_8529,N_8213,N_8177);
nand U8530 (N_8530,N_8160,N_8183);
or U8531 (N_8531,N_8181,N_8292);
xor U8532 (N_8532,N_8113,N_8360);
nand U8533 (N_8533,N_8101,N_8173);
nand U8534 (N_8534,N_8175,N_8268);
xor U8535 (N_8535,N_8162,N_8274);
nand U8536 (N_8536,N_8140,N_8374);
and U8537 (N_8537,N_8359,N_8189);
and U8538 (N_8538,N_8375,N_8214);
or U8539 (N_8539,N_8366,N_8178);
xnor U8540 (N_8540,N_8253,N_8299);
nand U8541 (N_8541,N_8266,N_8149);
nand U8542 (N_8542,N_8262,N_8390);
and U8543 (N_8543,N_8364,N_8350);
and U8544 (N_8544,N_8387,N_8388);
nor U8545 (N_8545,N_8392,N_8119);
and U8546 (N_8546,N_8397,N_8358);
nor U8547 (N_8547,N_8332,N_8244);
nor U8548 (N_8548,N_8346,N_8131);
nor U8549 (N_8549,N_8120,N_8207);
nand U8550 (N_8550,N_8305,N_8105);
and U8551 (N_8551,N_8130,N_8243);
or U8552 (N_8552,N_8248,N_8120);
nor U8553 (N_8553,N_8330,N_8396);
nand U8554 (N_8554,N_8264,N_8319);
and U8555 (N_8555,N_8188,N_8197);
and U8556 (N_8556,N_8159,N_8310);
and U8557 (N_8557,N_8290,N_8265);
or U8558 (N_8558,N_8332,N_8152);
or U8559 (N_8559,N_8186,N_8142);
or U8560 (N_8560,N_8363,N_8399);
or U8561 (N_8561,N_8207,N_8341);
xnor U8562 (N_8562,N_8340,N_8349);
nand U8563 (N_8563,N_8312,N_8368);
or U8564 (N_8564,N_8220,N_8312);
xor U8565 (N_8565,N_8336,N_8359);
nand U8566 (N_8566,N_8280,N_8150);
and U8567 (N_8567,N_8213,N_8378);
xnor U8568 (N_8568,N_8362,N_8131);
xor U8569 (N_8569,N_8158,N_8190);
nor U8570 (N_8570,N_8316,N_8333);
nor U8571 (N_8571,N_8112,N_8391);
or U8572 (N_8572,N_8324,N_8317);
and U8573 (N_8573,N_8135,N_8170);
xor U8574 (N_8574,N_8274,N_8147);
and U8575 (N_8575,N_8376,N_8340);
or U8576 (N_8576,N_8298,N_8294);
and U8577 (N_8577,N_8287,N_8299);
nand U8578 (N_8578,N_8232,N_8342);
and U8579 (N_8579,N_8195,N_8300);
and U8580 (N_8580,N_8174,N_8200);
nor U8581 (N_8581,N_8159,N_8369);
and U8582 (N_8582,N_8277,N_8280);
or U8583 (N_8583,N_8221,N_8392);
nand U8584 (N_8584,N_8331,N_8253);
nand U8585 (N_8585,N_8300,N_8216);
xnor U8586 (N_8586,N_8314,N_8213);
or U8587 (N_8587,N_8143,N_8147);
or U8588 (N_8588,N_8227,N_8372);
nand U8589 (N_8589,N_8153,N_8254);
or U8590 (N_8590,N_8336,N_8144);
xor U8591 (N_8591,N_8131,N_8200);
nor U8592 (N_8592,N_8146,N_8216);
xor U8593 (N_8593,N_8371,N_8316);
or U8594 (N_8594,N_8339,N_8308);
nand U8595 (N_8595,N_8365,N_8159);
xor U8596 (N_8596,N_8239,N_8123);
nand U8597 (N_8597,N_8268,N_8205);
or U8598 (N_8598,N_8180,N_8362);
nor U8599 (N_8599,N_8166,N_8308);
xnor U8600 (N_8600,N_8341,N_8122);
nand U8601 (N_8601,N_8213,N_8319);
nor U8602 (N_8602,N_8211,N_8224);
nor U8603 (N_8603,N_8127,N_8281);
nand U8604 (N_8604,N_8368,N_8362);
and U8605 (N_8605,N_8375,N_8177);
nand U8606 (N_8606,N_8342,N_8345);
xnor U8607 (N_8607,N_8163,N_8160);
nand U8608 (N_8608,N_8393,N_8261);
or U8609 (N_8609,N_8156,N_8394);
xor U8610 (N_8610,N_8100,N_8320);
xor U8611 (N_8611,N_8353,N_8358);
xor U8612 (N_8612,N_8363,N_8303);
xor U8613 (N_8613,N_8290,N_8387);
and U8614 (N_8614,N_8259,N_8151);
and U8615 (N_8615,N_8395,N_8193);
nor U8616 (N_8616,N_8252,N_8186);
xnor U8617 (N_8617,N_8235,N_8102);
xnor U8618 (N_8618,N_8384,N_8301);
nor U8619 (N_8619,N_8133,N_8354);
nand U8620 (N_8620,N_8374,N_8185);
xnor U8621 (N_8621,N_8383,N_8332);
xor U8622 (N_8622,N_8204,N_8269);
xor U8623 (N_8623,N_8184,N_8216);
and U8624 (N_8624,N_8296,N_8234);
nand U8625 (N_8625,N_8320,N_8283);
nor U8626 (N_8626,N_8357,N_8346);
xnor U8627 (N_8627,N_8369,N_8280);
and U8628 (N_8628,N_8135,N_8285);
nor U8629 (N_8629,N_8233,N_8247);
and U8630 (N_8630,N_8386,N_8128);
xnor U8631 (N_8631,N_8136,N_8308);
or U8632 (N_8632,N_8361,N_8387);
nor U8633 (N_8633,N_8377,N_8285);
xnor U8634 (N_8634,N_8357,N_8349);
xnor U8635 (N_8635,N_8204,N_8149);
and U8636 (N_8636,N_8180,N_8246);
and U8637 (N_8637,N_8208,N_8385);
nor U8638 (N_8638,N_8335,N_8259);
and U8639 (N_8639,N_8232,N_8278);
nor U8640 (N_8640,N_8388,N_8199);
xnor U8641 (N_8641,N_8122,N_8353);
nand U8642 (N_8642,N_8244,N_8241);
xnor U8643 (N_8643,N_8124,N_8361);
or U8644 (N_8644,N_8342,N_8374);
nor U8645 (N_8645,N_8109,N_8232);
nand U8646 (N_8646,N_8233,N_8361);
and U8647 (N_8647,N_8150,N_8360);
and U8648 (N_8648,N_8157,N_8322);
xor U8649 (N_8649,N_8126,N_8117);
or U8650 (N_8650,N_8309,N_8197);
nor U8651 (N_8651,N_8240,N_8235);
nor U8652 (N_8652,N_8191,N_8365);
nand U8653 (N_8653,N_8283,N_8211);
nand U8654 (N_8654,N_8153,N_8108);
and U8655 (N_8655,N_8103,N_8329);
or U8656 (N_8656,N_8273,N_8287);
nand U8657 (N_8657,N_8162,N_8115);
nor U8658 (N_8658,N_8195,N_8209);
or U8659 (N_8659,N_8161,N_8228);
xnor U8660 (N_8660,N_8379,N_8253);
and U8661 (N_8661,N_8126,N_8220);
nand U8662 (N_8662,N_8119,N_8248);
xnor U8663 (N_8663,N_8126,N_8210);
nor U8664 (N_8664,N_8245,N_8156);
or U8665 (N_8665,N_8318,N_8155);
or U8666 (N_8666,N_8103,N_8250);
nand U8667 (N_8667,N_8204,N_8265);
xnor U8668 (N_8668,N_8188,N_8175);
and U8669 (N_8669,N_8388,N_8167);
or U8670 (N_8670,N_8137,N_8178);
nand U8671 (N_8671,N_8313,N_8153);
or U8672 (N_8672,N_8219,N_8376);
nor U8673 (N_8673,N_8166,N_8267);
nand U8674 (N_8674,N_8360,N_8218);
and U8675 (N_8675,N_8128,N_8357);
nand U8676 (N_8676,N_8381,N_8101);
xnor U8677 (N_8677,N_8354,N_8100);
nor U8678 (N_8678,N_8151,N_8261);
nor U8679 (N_8679,N_8130,N_8248);
nand U8680 (N_8680,N_8318,N_8275);
nor U8681 (N_8681,N_8127,N_8341);
nor U8682 (N_8682,N_8233,N_8264);
and U8683 (N_8683,N_8136,N_8330);
xnor U8684 (N_8684,N_8297,N_8236);
or U8685 (N_8685,N_8109,N_8273);
nand U8686 (N_8686,N_8295,N_8134);
and U8687 (N_8687,N_8367,N_8133);
nor U8688 (N_8688,N_8217,N_8335);
or U8689 (N_8689,N_8175,N_8223);
nand U8690 (N_8690,N_8170,N_8238);
or U8691 (N_8691,N_8244,N_8136);
nor U8692 (N_8692,N_8199,N_8288);
or U8693 (N_8693,N_8317,N_8300);
or U8694 (N_8694,N_8365,N_8381);
or U8695 (N_8695,N_8230,N_8323);
and U8696 (N_8696,N_8115,N_8294);
nor U8697 (N_8697,N_8176,N_8218);
or U8698 (N_8698,N_8279,N_8101);
xor U8699 (N_8699,N_8376,N_8196);
nor U8700 (N_8700,N_8637,N_8664);
nand U8701 (N_8701,N_8523,N_8446);
and U8702 (N_8702,N_8692,N_8688);
and U8703 (N_8703,N_8682,N_8576);
nand U8704 (N_8704,N_8425,N_8528);
xor U8705 (N_8705,N_8615,N_8668);
xnor U8706 (N_8706,N_8421,N_8478);
nand U8707 (N_8707,N_8582,N_8594);
nand U8708 (N_8708,N_8550,N_8456);
xnor U8709 (N_8709,N_8424,N_8479);
xnor U8710 (N_8710,N_8548,N_8647);
or U8711 (N_8711,N_8572,N_8465);
or U8712 (N_8712,N_8649,N_8434);
nor U8713 (N_8713,N_8689,N_8524);
nor U8714 (N_8714,N_8498,N_8571);
or U8715 (N_8715,N_8448,N_8566);
or U8716 (N_8716,N_8665,N_8461);
nor U8717 (N_8717,N_8584,N_8451);
nor U8718 (N_8718,N_8629,N_8504);
nor U8719 (N_8719,N_8678,N_8640);
nor U8720 (N_8720,N_8501,N_8502);
or U8721 (N_8721,N_8454,N_8654);
nor U8722 (N_8722,N_8488,N_8507);
xor U8723 (N_8723,N_8441,N_8493);
nor U8724 (N_8724,N_8432,N_8557);
and U8725 (N_8725,N_8542,N_8540);
nor U8726 (N_8726,N_8453,N_8631);
nand U8727 (N_8727,N_8458,N_8574);
nand U8728 (N_8728,N_8402,N_8617);
xor U8729 (N_8729,N_8603,N_8477);
nand U8730 (N_8730,N_8568,N_8527);
nor U8731 (N_8731,N_8419,N_8552);
xnor U8732 (N_8732,N_8470,N_8623);
nand U8733 (N_8733,N_8522,N_8506);
xnor U8734 (N_8734,N_8619,N_8618);
and U8735 (N_8735,N_8436,N_8601);
nor U8736 (N_8736,N_8567,N_8683);
nor U8737 (N_8737,N_8691,N_8579);
and U8738 (N_8738,N_8455,N_8481);
or U8739 (N_8739,N_8559,N_8680);
nor U8740 (N_8740,N_8410,N_8467);
or U8741 (N_8741,N_8518,N_8437);
nor U8742 (N_8742,N_8652,N_8537);
and U8743 (N_8743,N_8643,N_8471);
xor U8744 (N_8744,N_8480,N_8677);
or U8745 (N_8745,N_8473,N_8575);
nor U8746 (N_8746,N_8696,N_8604);
or U8747 (N_8747,N_8610,N_8562);
nand U8748 (N_8748,N_8641,N_8476);
or U8749 (N_8749,N_8698,N_8492);
nor U8750 (N_8750,N_8433,N_8500);
and U8751 (N_8751,N_8491,N_8588);
and U8752 (N_8752,N_8521,N_8627);
or U8753 (N_8753,N_8685,N_8538);
and U8754 (N_8754,N_8636,N_8444);
nor U8755 (N_8755,N_8416,N_8485);
and U8756 (N_8756,N_8406,N_8529);
or U8757 (N_8757,N_8472,N_8580);
nor U8758 (N_8758,N_8534,N_8427);
and U8759 (N_8759,N_8560,N_8541);
nand U8760 (N_8760,N_8670,N_8577);
or U8761 (N_8761,N_8407,N_8551);
nand U8762 (N_8762,N_8586,N_8620);
and U8763 (N_8763,N_8558,N_8658);
nand U8764 (N_8764,N_8675,N_8663);
nor U8765 (N_8765,N_8442,N_8445);
and U8766 (N_8766,N_8602,N_8495);
xor U8767 (N_8767,N_8468,N_8638);
or U8768 (N_8768,N_8430,N_8535);
or U8769 (N_8769,N_8564,N_8694);
nand U8770 (N_8770,N_8447,N_8418);
nand U8771 (N_8771,N_8599,N_8639);
nand U8772 (N_8772,N_8517,N_8474);
nand U8773 (N_8773,N_8565,N_8549);
nand U8774 (N_8774,N_8686,N_8463);
nand U8775 (N_8775,N_8672,N_8484);
nor U8776 (N_8776,N_8578,N_8435);
and U8777 (N_8777,N_8657,N_8412);
nand U8778 (N_8778,N_8606,N_8699);
nor U8779 (N_8779,N_8648,N_8674);
and U8780 (N_8780,N_8431,N_8590);
xor U8781 (N_8781,N_8429,N_8642);
nor U8782 (N_8782,N_8547,N_8646);
nand U8783 (N_8783,N_8645,N_8612);
xor U8784 (N_8784,N_8400,N_8449);
or U8785 (N_8785,N_8581,N_8591);
xor U8786 (N_8786,N_8666,N_8519);
nor U8787 (N_8787,N_8555,N_8589);
xnor U8788 (N_8788,N_8530,N_8622);
or U8789 (N_8789,N_8462,N_8693);
xnor U8790 (N_8790,N_8650,N_8592);
or U8791 (N_8791,N_8625,N_8630);
xnor U8792 (N_8792,N_8597,N_8439);
and U8793 (N_8793,N_8553,N_8409);
xor U8794 (N_8794,N_8420,N_8614);
nor U8795 (N_8795,N_8525,N_8687);
nand U8796 (N_8796,N_8408,N_8405);
xnor U8797 (N_8797,N_8546,N_8673);
and U8798 (N_8798,N_8659,N_8561);
xnor U8799 (N_8799,N_8596,N_8452);
and U8800 (N_8800,N_8697,N_8684);
nor U8801 (N_8801,N_8450,N_8422);
xor U8802 (N_8802,N_8644,N_8624);
and U8803 (N_8803,N_8482,N_8514);
nor U8804 (N_8804,N_8516,N_8632);
or U8805 (N_8805,N_8403,N_8600);
nor U8806 (N_8806,N_8554,N_8633);
and U8807 (N_8807,N_8608,N_8413);
nor U8808 (N_8808,N_8613,N_8544);
xnor U8809 (N_8809,N_8426,N_8545);
nand U8810 (N_8810,N_8539,N_8499);
nand U8811 (N_8811,N_8526,N_8585);
nor U8812 (N_8812,N_8671,N_8628);
nand U8813 (N_8813,N_8616,N_8404);
xor U8814 (N_8814,N_8593,N_8512);
and U8815 (N_8815,N_8605,N_8563);
or U8816 (N_8816,N_8509,N_8469);
and U8817 (N_8817,N_8475,N_8513);
xor U8818 (N_8818,N_8459,N_8595);
and U8819 (N_8819,N_8634,N_8532);
and U8820 (N_8820,N_8440,N_8508);
xnor U8821 (N_8821,N_8653,N_8609);
nor U8822 (N_8822,N_8423,N_8415);
nand U8823 (N_8823,N_8669,N_8569);
nor U8824 (N_8824,N_8655,N_8443);
nand U8825 (N_8825,N_8661,N_8583);
xor U8826 (N_8826,N_8543,N_8679);
or U8827 (N_8827,N_8607,N_8662);
xnor U8828 (N_8828,N_8556,N_8681);
xor U8829 (N_8829,N_8536,N_8487);
nand U8830 (N_8830,N_8401,N_8428);
and U8831 (N_8831,N_8486,N_8466);
or U8832 (N_8832,N_8667,N_8457);
and U8833 (N_8833,N_8510,N_8483);
nand U8834 (N_8834,N_8460,N_8515);
nor U8835 (N_8835,N_8690,N_8651);
nor U8836 (N_8836,N_8490,N_8533);
xnor U8837 (N_8837,N_8531,N_8635);
nor U8838 (N_8838,N_8676,N_8570);
xor U8839 (N_8839,N_8494,N_8464);
and U8840 (N_8840,N_8621,N_8626);
nand U8841 (N_8841,N_8496,N_8497);
and U8842 (N_8842,N_8511,N_8656);
nor U8843 (N_8843,N_8411,N_8417);
nand U8844 (N_8844,N_8660,N_8695);
or U8845 (N_8845,N_8611,N_8573);
nor U8846 (N_8846,N_8414,N_8587);
and U8847 (N_8847,N_8489,N_8598);
nor U8848 (N_8848,N_8503,N_8505);
nor U8849 (N_8849,N_8438,N_8520);
xor U8850 (N_8850,N_8463,N_8650);
nor U8851 (N_8851,N_8478,N_8467);
or U8852 (N_8852,N_8470,N_8459);
nor U8853 (N_8853,N_8584,N_8676);
nor U8854 (N_8854,N_8544,N_8511);
xor U8855 (N_8855,N_8498,N_8584);
xor U8856 (N_8856,N_8457,N_8605);
xnor U8857 (N_8857,N_8623,N_8697);
and U8858 (N_8858,N_8515,N_8679);
or U8859 (N_8859,N_8431,N_8419);
nor U8860 (N_8860,N_8638,N_8596);
or U8861 (N_8861,N_8651,N_8685);
and U8862 (N_8862,N_8679,N_8500);
and U8863 (N_8863,N_8583,N_8406);
nand U8864 (N_8864,N_8547,N_8449);
nand U8865 (N_8865,N_8651,N_8580);
nor U8866 (N_8866,N_8542,N_8584);
nor U8867 (N_8867,N_8506,N_8553);
or U8868 (N_8868,N_8631,N_8515);
xnor U8869 (N_8869,N_8679,N_8598);
or U8870 (N_8870,N_8698,N_8519);
or U8871 (N_8871,N_8458,N_8410);
nor U8872 (N_8872,N_8671,N_8596);
nand U8873 (N_8873,N_8549,N_8546);
or U8874 (N_8874,N_8570,N_8551);
and U8875 (N_8875,N_8557,N_8506);
nor U8876 (N_8876,N_8460,N_8656);
and U8877 (N_8877,N_8586,N_8461);
nor U8878 (N_8878,N_8631,N_8537);
nand U8879 (N_8879,N_8460,N_8474);
and U8880 (N_8880,N_8504,N_8498);
nand U8881 (N_8881,N_8472,N_8426);
and U8882 (N_8882,N_8563,N_8547);
xnor U8883 (N_8883,N_8672,N_8450);
or U8884 (N_8884,N_8433,N_8464);
and U8885 (N_8885,N_8468,N_8619);
nand U8886 (N_8886,N_8515,N_8491);
or U8887 (N_8887,N_8682,N_8445);
and U8888 (N_8888,N_8485,N_8528);
nor U8889 (N_8889,N_8666,N_8400);
nor U8890 (N_8890,N_8572,N_8558);
xor U8891 (N_8891,N_8413,N_8618);
nand U8892 (N_8892,N_8481,N_8650);
nand U8893 (N_8893,N_8598,N_8686);
or U8894 (N_8894,N_8650,N_8670);
or U8895 (N_8895,N_8426,N_8543);
xor U8896 (N_8896,N_8537,N_8552);
nand U8897 (N_8897,N_8577,N_8658);
xnor U8898 (N_8898,N_8663,N_8487);
or U8899 (N_8899,N_8601,N_8405);
and U8900 (N_8900,N_8499,N_8689);
xor U8901 (N_8901,N_8536,N_8516);
xnor U8902 (N_8902,N_8621,N_8506);
nand U8903 (N_8903,N_8460,N_8429);
or U8904 (N_8904,N_8477,N_8544);
or U8905 (N_8905,N_8546,N_8525);
and U8906 (N_8906,N_8469,N_8660);
nand U8907 (N_8907,N_8576,N_8501);
or U8908 (N_8908,N_8423,N_8632);
and U8909 (N_8909,N_8685,N_8588);
xor U8910 (N_8910,N_8676,N_8681);
nor U8911 (N_8911,N_8577,N_8464);
xor U8912 (N_8912,N_8477,N_8532);
or U8913 (N_8913,N_8589,N_8539);
and U8914 (N_8914,N_8420,N_8433);
nand U8915 (N_8915,N_8685,N_8600);
xor U8916 (N_8916,N_8537,N_8461);
or U8917 (N_8917,N_8691,N_8690);
xor U8918 (N_8918,N_8643,N_8416);
nor U8919 (N_8919,N_8408,N_8699);
or U8920 (N_8920,N_8487,N_8569);
and U8921 (N_8921,N_8443,N_8615);
or U8922 (N_8922,N_8471,N_8688);
or U8923 (N_8923,N_8673,N_8465);
nand U8924 (N_8924,N_8657,N_8474);
and U8925 (N_8925,N_8436,N_8524);
xor U8926 (N_8926,N_8630,N_8519);
and U8927 (N_8927,N_8563,N_8509);
or U8928 (N_8928,N_8570,N_8577);
and U8929 (N_8929,N_8424,N_8557);
nand U8930 (N_8930,N_8691,N_8536);
or U8931 (N_8931,N_8502,N_8592);
or U8932 (N_8932,N_8670,N_8436);
xor U8933 (N_8933,N_8610,N_8516);
nor U8934 (N_8934,N_8542,N_8627);
and U8935 (N_8935,N_8590,N_8460);
nand U8936 (N_8936,N_8692,N_8433);
nor U8937 (N_8937,N_8409,N_8434);
nor U8938 (N_8938,N_8680,N_8417);
nor U8939 (N_8939,N_8603,N_8557);
nor U8940 (N_8940,N_8671,N_8423);
nand U8941 (N_8941,N_8585,N_8441);
nor U8942 (N_8942,N_8610,N_8611);
and U8943 (N_8943,N_8460,N_8588);
or U8944 (N_8944,N_8630,N_8440);
or U8945 (N_8945,N_8452,N_8639);
xnor U8946 (N_8946,N_8669,N_8527);
and U8947 (N_8947,N_8521,N_8460);
nor U8948 (N_8948,N_8668,N_8618);
xor U8949 (N_8949,N_8450,N_8671);
nand U8950 (N_8950,N_8602,N_8528);
xnor U8951 (N_8951,N_8418,N_8693);
or U8952 (N_8952,N_8441,N_8610);
nand U8953 (N_8953,N_8566,N_8642);
nand U8954 (N_8954,N_8632,N_8545);
nand U8955 (N_8955,N_8696,N_8595);
xnor U8956 (N_8956,N_8437,N_8487);
nand U8957 (N_8957,N_8671,N_8422);
and U8958 (N_8958,N_8415,N_8699);
or U8959 (N_8959,N_8433,N_8416);
nor U8960 (N_8960,N_8555,N_8538);
xnor U8961 (N_8961,N_8584,N_8579);
and U8962 (N_8962,N_8541,N_8486);
nor U8963 (N_8963,N_8420,N_8489);
nand U8964 (N_8964,N_8652,N_8481);
xor U8965 (N_8965,N_8561,N_8644);
or U8966 (N_8966,N_8631,N_8561);
and U8967 (N_8967,N_8492,N_8517);
xnor U8968 (N_8968,N_8498,N_8597);
and U8969 (N_8969,N_8517,N_8608);
or U8970 (N_8970,N_8545,N_8654);
or U8971 (N_8971,N_8601,N_8486);
and U8972 (N_8972,N_8541,N_8543);
xor U8973 (N_8973,N_8570,N_8483);
or U8974 (N_8974,N_8562,N_8403);
nor U8975 (N_8975,N_8538,N_8627);
and U8976 (N_8976,N_8675,N_8574);
nand U8977 (N_8977,N_8562,N_8515);
xor U8978 (N_8978,N_8425,N_8587);
nor U8979 (N_8979,N_8484,N_8523);
nor U8980 (N_8980,N_8483,N_8646);
and U8981 (N_8981,N_8531,N_8521);
or U8982 (N_8982,N_8699,N_8573);
and U8983 (N_8983,N_8661,N_8595);
and U8984 (N_8984,N_8678,N_8459);
and U8985 (N_8985,N_8690,N_8502);
or U8986 (N_8986,N_8558,N_8483);
and U8987 (N_8987,N_8409,N_8432);
nand U8988 (N_8988,N_8426,N_8580);
nor U8989 (N_8989,N_8687,N_8512);
xor U8990 (N_8990,N_8445,N_8627);
xor U8991 (N_8991,N_8577,N_8514);
xor U8992 (N_8992,N_8502,N_8484);
and U8993 (N_8993,N_8638,N_8476);
nor U8994 (N_8994,N_8477,N_8671);
nand U8995 (N_8995,N_8591,N_8418);
and U8996 (N_8996,N_8486,N_8567);
xor U8997 (N_8997,N_8621,N_8667);
and U8998 (N_8998,N_8629,N_8610);
nor U8999 (N_8999,N_8412,N_8568);
xnor U9000 (N_9000,N_8801,N_8755);
nand U9001 (N_9001,N_8826,N_8944);
nand U9002 (N_9002,N_8713,N_8783);
or U9003 (N_9003,N_8867,N_8973);
nand U9004 (N_9004,N_8721,N_8759);
nor U9005 (N_9005,N_8769,N_8991);
or U9006 (N_9006,N_8756,N_8817);
or U9007 (N_9007,N_8785,N_8833);
nor U9008 (N_9008,N_8834,N_8799);
and U9009 (N_9009,N_8966,N_8981);
and U9010 (N_9010,N_8749,N_8999);
nand U9011 (N_9011,N_8997,N_8731);
nand U9012 (N_9012,N_8923,N_8924);
nand U9013 (N_9013,N_8816,N_8881);
or U9014 (N_9014,N_8972,N_8908);
or U9015 (N_9015,N_8717,N_8959);
nand U9016 (N_9016,N_8800,N_8917);
or U9017 (N_9017,N_8748,N_8998);
and U9018 (N_9018,N_8821,N_8968);
and U9019 (N_9019,N_8847,N_8722);
xnor U9020 (N_9020,N_8876,N_8763);
and U9021 (N_9021,N_8711,N_8761);
and U9022 (N_9022,N_8980,N_8901);
xor U9023 (N_9023,N_8793,N_8762);
or U9024 (N_9024,N_8789,N_8878);
xor U9025 (N_9025,N_8928,N_8956);
nand U9026 (N_9026,N_8927,N_8774);
and U9027 (N_9027,N_8825,N_8712);
nand U9028 (N_9028,N_8898,N_8879);
nor U9029 (N_9029,N_8828,N_8845);
xor U9030 (N_9030,N_8839,N_8736);
and U9031 (N_9031,N_8855,N_8720);
nand U9032 (N_9032,N_8709,N_8880);
and U9033 (N_9033,N_8975,N_8773);
or U9034 (N_9034,N_8710,N_8910);
or U9035 (N_9035,N_8779,N_8951);
xor U9036 (N_9036,N_8838,N_8822);
nand U9037 (N_9037,N_8921,N_8814);
and U9038 (N_9038,N_8806,N_8895);
and U9039 (N_9039,N_8813,N_8940);
and U9040 (N_9040,N_8703,N_8704);
or U9041 (N_9041,N_8714,N_8708);
xnor U9042 (N_9042,N_8893,N_8729);
and U9043 (N_9043,N_8996,N_8915);
xnor U9044 (N_9044,N_8824,N_8848);
nand U9045 (N_9045,N_8738,N_8913);
xnor U9046 (N_9046,N_8970,N_8957);
nor U9047 (N_9047,N_8994,N_8877);
xnor U9048 (N_9048,N_8982,N_8752);
and U9049 (N_9049,N_8767,N_8757);
xor U9050 (N_9050,N_8850,N_8760);
nand U9051 (N_9051,N_8844,N_8835);
and U9052 (N_9052,N_8790,N_8952);
and U9053 (N_9053,N_8766,N_8819);
or U9054 (N_9054,N_8730,N_8791);
xor U9055 (N_9055,N_8931,N_8930);
or U9056 (N_9056,N_8914,N_8939);
xnor U9057 (N_9057,N_8772,N_8937);
xnor U9058 (N_9058,N_8700,N_8754);
nor U9059 (N_9059,N_8943,N_8912);
xor U9060 (N_9060,N_8853,N_8870);
xor U9061 (N_9061,N_8858,N_8836);
or U9062 (N_9062,N_8929,N_8865);
and U9063 (N_9063,N_8885,N_8967);
or U9064 (N_9064,N_8889,N_8891);
nor U9065 (N_9065,N_8784,N_8960);
xor U9066 (N_9066,N_8792,N_8753);
nand U9067 (N_9067,N_8932,N_8907);
nor U9068 (N_9068,N_8995,N_8740);
and U9069 (N_9069,N_8770,N_8707);
xor U9070 (N_9070,N_8742,N_8781);
nor U9071 (N_9071,N_8987,N_8827);
nand U9072 (N_9072,N_8808,N_8734);
and U9073 (N_9073,N_8984,N_8771);
and U9074 (N_9074,N_8977,N_8979);
nor U9075 (N_9075,N_8829,N_8747);
and U9076 (N_9076,N_8971,N_8884);
and U9077 (N_9077,N_8856,N_8925);
nor U9078 (N_9078,N_8948,N_8727);
nor U9079 (N_9079,N_8989,N_8776);
xnor U9080 (N_9080,N_8872,N_8715);
nand U9081 (N_9081,N_8724,N_8735);
or U9082 (N_9082,N_8905,N_8983);
nor U9083 (N_9083,N_8904,N_8843);
and U9084 (N_9084,N_8739,N_8963);
nand U9085 (N_9085,N_8886,N_8765);
nor U9086 (N_9086,N_8725,N_8933);
or U9087 (N_9087,N_8892,N_8955);
xor U9088 (N_9088,N_8811,N_8902);
or U9089 (N_9089,N_8744,N_8807);
xor U9090 (N_9090,N_8859,N_8887);
nor U9091 (N_9091,N_8920,N_8961);
or U9092 (N_9092,N_8860,N_8949);
nor U9093 (N_9093,N_8954,N_8976);
or U9094 (N_9094,N_8906,N_8726);
and U9095 (N_9095,N_8716,N_8849);
nand U9096 (N_9096,N_8818,N_8863);
nand U9097 (N_9097,N_8798,N_8974);
nor U9098 (N_9098,N_8823,N_8841);
or U9099 (N_9099,N_8986,N_8953);
nor U9100 (N_9100,N_8926,N_8861);
and U9101 (N_9101,N_8992,N_8840);
nor U9102 (N_9102,N_8851,N_8705);
or U9103 (N_9103,N_8810,N_8899);
and U9104 (N_9104,N_8882,N_8751);
or U9105 (N_9105,N_8750,N_8922);
nor U9106 (N_9106,N_8888,N_8719);
nand U9107 (N_9107,N_8775,N_8702);
and U9108 (N_9108,N_8780,N_8862);
or U9109 (N_9109,N_8778,N_8869);
or U9110 (N_9110,N_8797,N_8978);
nor U9111 (N_9111,N_8936,N_8786);
and U9112 (N_9112,N_8890,N_8965);
nand U9113 (N_9113,N_8874,N_8815);
nand U9114 (N_9114,N_8962,N_8897);
nand U9115 (N_9115,N_8846,N_8894);
nand U9116 (N_9116,N_8728,N_8741);
and U9117 (N_9117,N_8758,N_8875);
or U9118 (N_9118,N_8871,N_8988);
or U9119 (N_9119,N_8732,N_8900);
nand U9120 (N_9120,N_8903,N_8916);
and U9121 (N_9121,N_8883,N_8934);
xor U9122 (N_9122,N_8868,N_8802);
xor U9123 (N_9123,N_8854,N_8935);
and U9124 (N_9124,N_8909,N_8942);
xnor U9125 (N_9125,N_8803,N_8896);
xnor U9126 (N_9126,N_8852,N_8985);
xor U9127 (N_9127,N_8873,N_8969);
or U9128 (N_9128,N_8794,N_8788);
nand U9129 (N_9129,N_8911,N_8919);
nand U9130 (N_9130,N_8820,N_8764);
and U9131 (N_9131,N_8743,N_8706);
and U9132 (N_9132,N_8964,N_8857);
and U9133 (N_9133,N_8864,N_8918);
xnor U9134 (N_9134,N_8795,N_8768);
nor U9135 (N_9135,N_8830,N_8805);
and U9136 (N_9136,N_8777,N_8812);
xnor U9137 (N_9137,N_8746,N_8745);
nor U9138 (N_9138,N_8804,N_8993);
xnor U9139 (N_9139,N_8958,N_8723);
and U9140 (N_9140,N_8831,N_8796);
and U9141 (N_9141,N_8990,N_8832);
or U9142 (N_9142,N_8945,N_8787);
nor U9143 (N_9143,N_8950,N_8733);
nand U9144 (N_9144,N_8809,N_8941);
and U9145 (N_9145,N_8837,N_8947);
nor U9146 (N_9146,N_8782,N_8938);
nor U9147 (N_9147,N_8946,N_8718);
or U9148 (N_9148,N_8701,N_8866);
and U9149 (N_9149,N_8737,N_8842);
and U9150 (N_9150,N_8781,N_8851);
nor U9151 (N_9151,N_8734,N_8790);
and U9152 (N_9152,N_8926,N_8822);
or U9153 (N_9153,N_8784,N_8982);
and U9154 (N_9154,N_8974,N_8713);
and U9155 (N_9155,N_8895,N_8918);
or U9156 (N_9156,N_8701,N_8916);
or U9157 (N_9157,N_8796,N_8958);
nand U9158 (N_9158,N_8705,N_8948);
nor U9159 (N_9159,N_8920,N_8747);
or U9160 (N_9160,N_8715,N_8844);
nand U9161 (N_9161,N_8868,N_8904);
nor U9162 (N_9162,N_8830,N_8943);
xor U9163 (N_9163,N_8882,N_8707);
nor U9164 (N_9164,N_8775,N_8903);
nor U9165 (N_9165,N_8969,N_8906);
nand U9166 (N_9166,N_8996,N_8958);
xor U9167 (N_9167,N_8795,N_8746);
and U9168 (N_9168,N_8883,N_8956);
nor U9169 (N_9169,N_8918,N_8932);
or U9170 (N_9170,N_8721,N_8971);
or U9171 (N_9171,N_8774,N_8713);
nor U9172 (N_9172,N_8997,N_8925);
xnor U9173 (N_9173,N_8771,N_8842);
and U9174 (N_9174,N_8917,N_8930);
or U9175 (N_9175,N_8857,N_8977);
xor U9176 (N_9176,N_8725,N_8864);
and U9177 (N_9177,N_8921,N_8965);
and U9178 (N_9178,N_8766,N_8908);
or U9179 (N_9179,N_8755,N_8915);
xor U9180 (N_9180,N_8957,N_8850);
and U9181 (N_9181,N_8788,N_8810);
xor U9182 (N_9182,N_8990,N_8821);
xor U9183 (N_9183,N_8932,N_8977);
and U9184 (N_9184,N_8960,N_8771);
and U9185 (N_9185,N_8743,N_8962);
nor U9186 (N_9186,N_8865,N_8831);
xor U9187 (N_9187,N_8713,N_8902);
and U9188 (N_9188,N_8949,N_8880);
xor U9189 (N_9189,N_8999,N_8758);
nor U9190 (N_9190,N_8913,N_8707);
and U9191 (N_9191,N_8779,N_8923);
and U9192 (N_9192,N_8944,N_8960);
nand U9193 (N_9193,N_8900,N_8830);
or U9194 (N_9194,N_8773,N_8753);
or U9195 (N_9195,N_8934,N_8900);
and U9196 (N_9196,N_8719,N_8797);
or U9197 (N_9197,N_8841,N_8886);
or U9198 (N_9198,N_8851,N_8850);
nor U9199 (N_9199,N_8860,N_8794);
xnor U9200 (N_9200,N_8846,N_8863);
nor U9201 (N_9201,N_8956,N_8762);
xor U9202 (N_9202,N_8942,N_8711);
or U9203 (N_9203,N_8762,N_8873);
and U9204 (N_9204,N_8999,N_8943);
nand U9205 (N_9205,N_8967,N_8897);
or U9206 (N_9206,N_8739,N_8988);
and U9207 (N_9207,N_8745,N_8973);
and U9208 (N_9208,N_8962,N_8724);
or U9209 (N_9209,N_8905,N_8935);
nand U9210 (N_9210,N_8875,N_8841);
or U9211 (N_9211,N_8946,N_8959);
nor U9212 (N_9212,N_8728,N_8822);
or U9213 (N_9213,N_8965,N_8728);
and U9214 (N_9214,N_8820,N_8921);
nor U9215 (N_9215,N_8789,N_8723);
nor U9216 (N_9216,N_8829,N_8808);
xor U9217 (N_9217,N_8753,N_8876);
xor U9218 (N_9218,N_8828,N_8818);
nor U9219 (N_9219,N_8831,N_8972);
xor U9220 (N_9220,N_8789,N_8826);
xnor U9221 (N_9221,N_8972,N_8912);
nand U9222 (N_9222,N_8853,N_8840);
xnor U9223 (N_9223,N_8803,N_8793);
xnor U9224 (N_9224,N_8750,N_8855);
and U9225 (N_9225,N_8816,N_8815);
and U9226 (N_9226,N_8816,N_8755);
nor U9227 (N_9227,N_8941,N_8709);
and U9228 (N_9228,N_8744,N_8960);
and U9229 (N_9229,N_8783,N_8700);
xnor U9230 (N_9230,N_8757,N_8761);
xnor U9231 (N_9231,N_8852,N_8868);
or U9232 (N_9232,N_8766,N_8818);
nand U9233 (N_9233,N_8783,N_8735);
nand U9234 (N_9234,N_8714,N_8773);
nor U9235 (N_9235,N_8993,N_8778);
xor U9236 (N_9236,N_8984,N_8877);
and U9237 (N_9237,N_8832,N_8739);
nand U9238 (N_9238,N_8822,N_8813);
or U9239 (N_9239,N_8880,N_8929);
and U9240 (N_9240,N_8819,N_8812);
nand U9241 (N_9241,N_8770,N_8782);
or U9242 (N_9242,N_8815,N_8854);
nand U9243 (N_9243,N_8829,N_8955);
and U9244 (N_9244,N_8755,N_8962);
nor U9245 (N_9245,N_8778,N_8949);
nor U9246 (N_9246,N_8961,N_8818);
nand U9247 (N_9247,N_8921,N_8705);
and U9248 (N_9248,N_8943,N_8705);
nand U9249 (N_9249,N_8945,N_8814);
or U9250 (N_9250,N_8726,N_8905);
nand U9251 (N_9251,N_8835,N_8941);
nor U9252 (N_9252,N_8843,N_8956);
nand U9253 (N_9253,N_8947,N_8714);
and U9254 (N_9254,N_8827,N_8884);
xor U9255 (N_9255,N_8710,N_8954);
xor U9256 (N_9256,N_8903,N_8870);
and U9257 (N_9257,N_8716,N_8893);
or U9258 (N_9258,N_8812,N_8853);
nand U9259 (N_9259,N_8770,N_8843);
nand U9260 (N_9260,N_8725,N_8794);
nor U9261 (N_9261,N_8759,N_8787);
nor U9262 (N_9262,N_8731,N_8882);
or U9263 (N_9263,N_8872,N_8780);
and U9264 (N_9264,N_8968,N_8708);
nand U9265 (N_9265,N_8755,N_8860);
xor U9266 (N_9266,N_8798,N_8961);
nor U9267 (N_9267,N_8909,N_8718);
nor U9268 (N_9268,N_8825,N_8844);
xnor U9269 (N_9269,N_8764,N_8923);
xor U9270 (N_9270,N_8857,N_8861);
nand U9271 (N_9271,N_8948,N_8778);
nor U9272 (N_9272,N_8859,N_8949);
or U9273 (N_9273,N_8705,N_8732);
or U9274 (N_9274,N_8869,N_8918);
xnor U9275 (N_9275,N_8727,N_8754);
or U9276 (N_9276,N_8978,N_8901);
nand U9277 (N_9277,N_8931,N_8759);
nand U9278 (N_9278,N_8749,N_8704);
nor U9279 (N_9279,N_8778,N_8712);
nor U9280 (N_9280,N_8984,N_8802);
or U9281 (N_9281,N_8765,N_8846);
and U9282 (N_9282,N_8925,N_8834);
and U9283 (N_9283,N_8844,N_8819);
or U9284 (N_9284,N_8850,N_8971);
nand U9285 (N_9285,N_8977,N_8749);
or U9286 (N_9286,N_8816,N_8925);
or U9287 (N_9287,N_8897,N_8830);
or U9288 (N_9288,N_8889,N_8997);
xnor U9289 (N_9289,N_8746,N_8847);
or U9290 (N_9290,N_8744,N_8813);
and U9291 (N_9291,N_8951,N_8956);
nand U9292 (N_9292,N_8845,N_8837);
xnor U9293 (N_9293,N_8780,N_8940);
and U9294 (N_9294,N_8915,N_8939);
or U9295 (N_9295,N_8862,N_8934);
nand U9296 (N_9296,N_8735,N_8763);
nor U9297 (N_9297,N_8809,N_8706);
xor U9298 (N_9298,N_8896,N_8931);
or U9299 (N_9299,N_8837,N_8720);
nor U9300 (N_9300,N_9294,N_9217);
xnor U9301 (N_9301,N_9163,N_9154);
and U9302 (N_9302,N_9110,N_9033);
xor U9303 (N_9303,N_9038,N_9075);
or U9304 (N_9304,N_9046,N_9172);
nand U9305 (N_9305,N_9288,N_9167);
xor U9306 (N_9306,N_9067,N_9203);
nand U9307 (N_9307,N_9042,N_9199);
or U9308 (N_9308,N_9099,N_9037);
and U9309 (N_9309,N_9202,N_9159);
nand U9310 (N_9310,N_9255,N_9149);
nor U9311 (N_9311,N_9086,N_9185);
and U9312 (N_9312,N_9162,N_9239);
nor U9313 (N_9313,N_9122,N_9085);
and U9314 (N_9314,N_9137,N_9136);
nor U9315 (N_9315,N_9277,N_9032);
xor U9316 (N_9316,N_9257,N_9230);
xnor U9317 (N_9317,N_9215,N_9201);
nand U9318 (N_9318,N_9283,N_9270);
and U9319 (N_9319,N_9226,N_9282);
nor U9320 (N_9320,N_9152,N_9015);
xor U9321 (N_9321,N_9285,N_9281);
or U9322 (N_9322,N_9054,N_9145);
nand U9323 (N_9323,N_9036,N_9275);
nor U9324 (N_9324,N_9263,N_9092);
nand U9325 (N_9325,N_9237,N_9018);
nand U9326 (N_9326,N_9213,N_9229);
or U9327 (N_9327,N_9168,N_9048);
xor U9328 (N_9328,N_9000,N_9095);
xor U9329 (N_9329,N_9200,N_9039);
nor U9330 (N_9330,N_9093,N_9076);
or U9331 (N_9331,N_9197,N_9274);
or U9332 (N_9332,N_9296,N_9125);
nor U9333 (N_9333,N_9141,N_9166);
xnor U9334 (N_9334,N_9248,N_9132);
or U9335 (N_9335,N_9266,N_9205);
nor U9336 (N_9336,N_9254,N_9004);
and U9337 (N_9337,N_9026,N_9105);
and U9338 (N_9338,N_9279,N_9135);
nor U9339 (N_9339,N_9102,N_9051);
nand U9340 (N_9340,N_9251,N_9225);
and U9341 (N_9341,N_9078,N_9264);
nand U9342 (N_9342,N_9118,N_9231);
and U9343 (N_9343,N_9252,N_9035);
xor U9344 (N_9344,N_9169,N_9227);
or U9345 (N_9345,N_9209,N_9176);
and U9346 (N_9346,N_9216,N_9009);
and U9347 (N_9347,N_9190,N_9265);
and U9348 (N_9348,N_9074,N_9187);
nor U9349 (N_9349,N_9043,N_9045);
nand U9350 (N_9350,N_9170,N_9047);
nand U9351 (N_9351,N_9193,N_9220);
and U9352 (N_9352,N_9267,N_9134);
nand U9353 (N_9353,N_9029,N_9082);
xor U9354 (N_9354,N_9147,N_9208);
nor U9355 (N_9355,N_9072,N_9040);
or U9356 (N_9356,N_9014,N_9222);
and U9357 (N_9357,N_9057,N_9269);
nand U9358 (N_9358,N_9174,N_9061);
nand U9359 (N_9359,N_9240,N_9272);
nor U9360 (N_9360,N_9052,N_9089);
and U9361 (N_9361,N_9184,N_9115);
or U9362 (N_9362,N_9025,N_9242);
and U9363 (N_9363,N_9073,N_9234);
nor U9364 (N_9364,N_9148,N_9022);
nor U9365 (N_9365,N_9010,N_9210);
nand U9366 (N_9366,N_9214,N_9001);
or U9367 (N_9367,N_9293,N_9101);
nor U9368 (N_9368,N_9084,N_9117);
and U9369 (N_9369,N_9171,N_9273);
xor U9370 (N_9370,N_9256,N_9188);
nor U9371 (N_9371,N_9005,N_9276);
nand U9372 (N_9372,N_9204,N_9080);
nor U9373 (N_9373,N_9056,N_9280);
xor U9374 (N_9374,N_9183,N_9060);
nor U9375 (N_9375,N_9070,N_9112);
nand U9376 (N_9376,N_9278,N_9238);
nand U9377 (N_9377,N_9108,N_9262);
nand U9378 (N_9378,N_9245,N_9103);
xnor U9379 (N_9379,N_9151,N_9104);
or U9380 (N_9380,N_9059,N_9156);
nor U9381 (N_9381,N_9268,N_9109);
or U9382 (N_9382,N_9153,N_9123);
nor U9383 (N_9383,N_9027,N_9236);
xor U9384 (N_9384,N_9195,N_9250);
and U9385 (N_9385,N_9116,N_9003);
or U9386 (N_9386,N_9142,N_9131);
nor U9387 (N_9387,N_9299,N_9058);
and U9388 (N_9388,N_9194,N_9140);
or U9389 (N_9389,N_9207,N_9191);
and U9390 (N_9390,N_9287,N_9212);
xnor U9391 (N_9391,N_9249,N_9106);
nand U9392 (N_9392,N_9120,N_9077);
or U9393 (N_9393,N_9081,N_9121);
nor U9394 (N_9394,N_9062,N_9177);
nand U9395 (N_9395,N_9011,N_9138);
or U9396 (N_9396,N_9161,N_9111);
nor U9397 (N_9397,N_9087,N_9007);
nor U9398 (N_9398,N_9083,N_9126);
xnor U9399 (N_9399,N_9139,N_9173);
and U9400 (N_9400,N_9016,N_9066);
and U9401 (N_9401,N_9253,N_9259);
nand U9402 (N_9402,N_9098,N_9164);
nor U9403 (N_9403,N_9198,N_9019);
or U9404 (N_9404,N_9258,N_9063);
xor U9405 (N_9405,N_9157,N_9144);
and U9406 (N_9406,N_9069,N_9097);
nor U9407 (N_9407,N_9224,N_9064);
xor U9408 (N_9408,N_9289,N_9295);
or U9409 (N_9409,N_9002,N_9178);
nor U9410 (N_9410,N_9179,N_9182);
xor U9411 (N_9411,N_9020,N_9119);
and U9412 (N_9412,N_9206,N_9053);
and U9413 (N_9413,N_9133,N_9124);
xor U9414 (N_9414,N_9013,N_9271);
or U9415 (N_9415,N_9290,N_9291);
nand U9416 (N_9416,N_9247,N_9050);
nand U9417 (N_9417,N_9079,N_9286);
xnor U9418 (N_9418,N_9127,N_9243);
nor U9419 (N_9419,N_9186,N_9219);
xor U9420 (N_9420,N_9006,N_9071);
nor U9421 (N_9421,N_9260,N_9146);
xnor U9422 (N_9422,N_9088,N_9114);
and U9423 (N_9423,N_9246,N_9100);
and U9424 (N_9424,N_9158,N_9041);
xnor U9425 (N_9425,N_9223,N_9091);
nor U9426 (N_9426,N_9030,N_9155);
xnor U9427 (N_9427,N_9192,N_9021);
xnor U9428 (N_9428,N_9297,N_9284);
nor U9429 (N_9429,N_9189,N_9024);
nor U9430 (N_9430,N_9008,N_9044);
and U9431 (N_9431,N_9128,N_9107);
nor U9432 (N_9432,N_9096,N_9143);
or U9433 (N_9433,N_9160,N_9065);
nor U9434 (N_9434,N_9221,N_9232);
nand U9435 (N_9435,N_9094,N_9023);
nor U9436 (N_9436,N_9175,N_9068);
nand U9437 (N_9437,N_9012,N_9235);
nand U9438 (N_9438,N_9049,N_9031);
nor U9439 (N_9439,N_9113,N_9090);
nor U9440 (N_9440,N_9211,N_9028);
xor U9441 (N_9441,N_9233,N_9129);
xnor U9442 (N_9442,N_9261,N_9180);
xnor U9443 (N_9443,N_9150,N_9292);
xnor U9444 (N_9444,N_9055,N_9228);
nand U9445 (N_9445,N_9218,N_9034);
nand U9446 (N_9446,N_9017,N_9130);
or U9447 (N_9447,N_9165,N_9244);
nand U9448 (N_9448,N_9298,N_9181);
and U9449 (N_9449,N_9241,N_9196);
nand U9450 (N_9450,N_9202,N_9115);
and U9451 (N_9451,N_9192,N_9024);
nand U9452 (N_9452,N_9234,N_9014);
nand U9453 (N_9453,N_9089,N_9050);
and U9454 (N_9454,N_9186,N_9093);
xor U9455 (N_9455,N_9167,N_9231);
nor U9456 (N_9456,N_9174,N_9203);
and U9457 (N_9457,N_9206,N_9151);
and U9458 (N_9458,N_9120,N_9243);
xor U9459 (N_9459,N_9055,N_9034);
or U9460 (N_9460,N_9261,N_9032);
nor U9461 (N_9461,N_9277,N_9186);
xor U9462 (N_9462,N_9248,N_9285);
and U9463 (N_9463,N_9027,N_9222);
and U9464 (N_9464,N_9152,N_9029);
nor U9465 (N_9465,N_9122,N_9143);
nor U9466 (N_9466,N_9026,N_9123);
and U9467 (N_9467,N_9224,N_9267);
and U9468 (N_9468,N_9030,N_9217);
or U9469 (N_9469,N_9191,N_9087);
and U9470 (N_9470,N_9161,N_9285);
and U9471 (N_9471,N_9255,N_9223);
and U9472 (N_9472,N_9091,N_9088);
or U9473 (N_9473,N_9234,N_9089);
nor U9474 (N_9474,N_9275,N_9243);
nor U9475 (N_9475,N_9153,N_9030);
and U9476 (N_9476,N_9220,N_9200);
nand U9477 (N_9477,N_9025,N_9043);
xnor U9478 (N_9478,N_9028,N_9164);
nor U9479 (N_9479,N_9126,N_9166);
xnor U9480 (N_9480,N_9234,N_9038);
and U9481 (N_9481,N_9001,N_9027);
and U9482 (N_9482,N_9087,N_9136);
nor U9483 (N_9483,N_9187,N_9121);
or U9484 (N_9484,N_9004,N_9002);
nor U9485 (N_9485,N_9080,N_9183);
or U9486 (N_9486,N_9047,N_9262);
and U9487 (N_9487,N_9283,N_9121);
xnor U9488 (N_9488,N_9279,N_9066);
and U9489 (N_9489,N_9140,N_9117);
nand U9490 (N_9490,N_9072,N_9202);
xor U9491 (N_9491,N_9125,N_9092);
nor U9492 (N_9492,N_9227,N_9253);
nand U9493 (N_9493,N_9185,N_9275);
and U9494 (N_9494,N_9190,N_9169);
or U9495 (N_9495,N_9196,N_9244);
nor U9496 (N_9496,N_9245,N_9184);
and U9497 (N_9497,N_9235,N_9069);
nand U9498 (N_9498,N_9029,N_9031);
or U9499 (N_9499,N_9273,N_9162);
nand U9500 (N_9500,N_9269,N_9001);
or U9501 (N_9501,N_9156,N_9092);
nand U9502 (N_9502,N_9212,N_9184);
or U9503 (N_9503,N_9107,N_9113);
and U9504 (N_9504,N_9172,N_9189);
and U9505 (N_9505,N_9194,N_9059);
or U9506 (N_9506,N_9091,N_9200);
xor U9507 (N_9507,N_9025,N_9079);
nand U9508 (N_9508,N_9287,N_9279);
or U9509 (N_9509,N_9277,N_9219);
or U9510 (N_9510,N_9132,N_9247);
nor U9511 (N_9511,N_9289,N_9197);
nand U9512 (N_9512,N_9141,N_9267);
nor U9513 (N_9513,N_9063,N_9227);
and U9514 (N_9514,N_9213,N_9237);
and U9515 (N_9515,N_9077,N_9082);
and U9516 (N_9516,N_9100,N_9193);
or U9517 (N_9517,N_9041,N_9234);
or U9518 (N_9518,N_9110,N_9082);
or U9519 (N_9519,N_9024,N_9221);
nand U9520 (N_9520,N_9020,N_9286);
nand U9521 (N_9521,N_9206,N_9294);
xor U9522 (N_9522,N_9065,N_9063);
xnor U9523 (N_9523,N_9161,N_9073);
nand U9524 (N_9524,N_9125,N_9286);
nor U9525 (N_9525,N_9008,N_9094);
or U9526 (N_9526,N_9208,N_9045);
xor U9527 (N_9527,N_9130,N_9299);
or U9528 (N_9528,N_9214,N_9150);
or U9529 (N_9529,N_9150,N_9299);
nor U9530 (N_9530,N_9197,N_9278);
or U9531 (N_9531,N_9178,N_9240);
or U9532 (N_9532,N_9261,N_9270);
or U9533 (N_9533,N_9271,N_9240);
xor U9534 (N_9534,N_9016,N_9279);
nor U9535 (N_9535,N_9032,N_9109);
xor U9536 (N_9536,N_9064,N_9112);
nor U9537 (N_9537,N_9023,N_9271);
xnor U9538 (N_9538,N_9094,N_9257);
nor U9539 (N_9539,N_9105,N_9265);
nor U9540 (N_9540,N_9116,N_9290);
nand U9541 (N_9541,N_9125,N_9021);
nand U9542 (N_9542,N_9290,N_9101);
and U9543 (N_9543,N_9295,N_9028);
xnor U9544 (N_9544,N_9202,N_9158);
or U9545 (N_9545,N_9091,N_9023);
nand U9546 (N_9546,N_9098,N_9248);
nand U9547 (N_9547,N_9179,N_9253);
xor U9548 (N_9548,N_9066,N_9175);
nand U9549 (N_9549,N_9277,N_9207);
and U9550 (N_9550,N_9135,N_9266);
nor U9551 (N_9551,N_9117,N_9214);
and U9552 (N_9552,N_9155,N_9119);
xnor U9553 (N_9553,N_9195,N_9013);
and U9554 (N_9554,N_9245,N_9015);
or U9555 (N_9555,N_9105,N_9078);
xnor U9556 (N_9556,N_9030,N_9052);
and U9557 (N_9557,N_9259,N_9080);
and U9558 (N_9558,N_9098,N_9113);
or U9559 (N_9559,N_9075,N_9227);
nor U9560 (N_9560,N_9056,N_9024);
nor U9561 (N_9561,N_9275,N_9058);
or U9562 (N_9562,N_9100,N_9223);
nand U9563 (N_9563,N_9172,N_9073);
and U9564 (N_9564,N_9274,N_9222);
and U9565 (N_9565,N_9193,N_9098);
and U9566 (N_9566,N_9089,N_9280);
and U9567 (N_9567,N_9271,N_9136);
nand U9568 (N_9568,N_9292,N_9031);
nand U9569 (N_9569,N_9113,N_9128);
nor U9570 (N_9570,N_9027,N_9102);
nand U9571 (N_9571,N_9152,N_9018);
nand U9572 (N_9572,N_9184,N_9131);
xnor U9573 (N_9573,N_9091,N_9258);
and U9574 (N_9574,N_9184,N_9022);
and U9575 (N_9575,N_9003,N_9257);
nand U9576 (N_9576,N_9290,N_9006);
or U9577 (N_9577,N_9041,N_9214);
nand U9578 (N_9578,N_9262,N_9066);
and U9579 (N_9579,N_9143,N_9167);
and U9580 (N_9580,N_9180,N_9249);
xnor U9581 (N_9581,N_9116,N_9210);
or U9582 (N_9582,N_9086,N_9000);
xnor U9583 (N_9583,N_9262,N_9266);
xor U9584 (N_9584,N_9086,N_9178);
nand U9585 (N_9585,N_9030,N_9163);
or U9586 (N_9586,N_9216,N_9276);
and U9587 (N_9587,N_9048,N_9109);
xor U9588 (N_9588,N_9005,N_9213);
or U9589 (N_9589,N_9150,N_9144);
xor U9590 (N_9590,N_9032,N_9252);
nor U9591 (N_9591,N_9239,N_9191);
xor U9592 (N_9592,N_9240,N_9126);
nor U9593 (N_9593,N_9057,N_9145);
nor U9594 (N_9594,N_9143,N_9273);
xor U9595 (N_9595,N_9261,N_9265);
nor U9596 (N_9596,N_9192,N_9017);
or U9597 (N_9597,N_9107,N_9117);
nor U9598 (N_9598,N_9295,N_9041);
xnor U9599 (N_9599,N_9254,N_9152);
or U9600 (N_9600,N_9598,N_9327);
and U9601 (N_9601,N_9574,N_9521);
nand U9602 (N_9602,N_9566,N_9539);
or U9603 (N_9603,N_9340,N_9302);
xnor U9604 (N_9604,N_9424,N_9338);
and U9605 (N_9605,N_9357,N_9353);
or U9606 (N_9606,N_9569,N_9456);
or U9607 (N_9607,N_9570,N_9467);
or U9608 (N_9608,N_9563,N_9323);
xor U9609 (N_9609,N_9442,N_9422);
nand U9610 (N_9610,N_9313,N_9520);
nor U9611 (N_9611,N_9492,N_9334);
xor U9612 (N_9612,N_9412,N_9317);
xor U9613 (N_9613,N_9502,N_9330);
nand U9614 (N_9614,N_9537,N_9371);
and U9615 (N_9615,N_9562,N_9505);
nor U9616 (N_9616,N_9497,N_9361);
and U9617 (N_9617,N_9420,N_9465);
and U9618 (N_9618,N_9552,N_9413);
nand U9619 (N_9619,N_9544,N_9447);
xor U9620 (N_9620,N_9540,N_9386);
or U9621 (N_9621,N_9364,N_9575);
xnor U9622 (N_9622,N_9564,N_9449);
or U9623 (N_9623,N_9488,N_9428);
nand U9624 (N_9624,N_9446,N_9518);
or U9625 (N_9625,N_9304,N_9486);
nor U9626 (N_9626,N_9565,N_9365);
nor U9627 (N_9627,N_9337,N_9469);
xnor U9628 (N_9628,N_9410,N_9438);
and U9629 (N_9629,N_9587,N_9345);
xor U9630 (N_9630,N_9470,N_9431);
and U9631 (N_9631,N_9579,N_9557);
and U9632 (N_9632,N_9362,N_9400);
xor U9633 (N_9633,N_9390,N_9310);
xnor U9634 (N_9634,N_9483,N_9545);
nand U9635 (N_9635,N_9482,N_9439);
nand U9636 (N_9636,N_9528,N_9315);
or U9637 (N_9637,N_9454,N_9550);
or U9638 (N_9638,N_9331,N_9382);
or U9639 (N_9639,N_9335,N_9504);
nor U9640 (N_9640,N_9395,N_9584);
or U9641 (N_9641,N_9393,N_9548);
or U9642 (N_9642,N_9402,N_9450);
or U9643 (N_9643,N_9534,N_9326);
xnor U9644 (N_9644,N_9491,N_9307);
nor U9645 (N_9645,N_9549,N_9471);
or U9646 (N_9646,N_9383,N_9527);
and U9647 (N_9647,N_9476,N_9509);
or U9648 (N_9648,N_9592,N_9322);
xnor U9649 (N_9649,N_9347,N_9519);
nor U9650 (N_9650,N_9358,N_9464);
xnor U9651 (N_9651,N_9314,N_9378);
and U9652 (N_9652,N_9484,N_9372);
or U9653 (N_9653,N_9342,N_9455);
nand U9654 (N_9654,N_9384,N_9501);
nand U9655 (N_9655,N_9517,N_9498);
nand U9656 (N_9656,N_9558,N_9434);
and U9657 (N_9657,N_9418,N_9503);
xor U9658 (N_9658,N_9419,N_9524);
and U9659 (N_9659,N_9523,N_9405);
nand U9660 (N_9660,N_9485,N_9453);
nand U9661 (N_9661,N_9487,N_9448);
or U9662 (N_9662,N_9332,N_9568);
or U9663 (N_9663,N_9514,N_9481);
nand U9664 (N_9664,N_9445,N_9573);
nor U9665 (N_9665,N_9468,N_9451);
and U9666 (N_9666,N_9588,N_9379);
or U9667 (N_9667,N_9586,N_9407);
xnor U9668 (N_9668,N_9321,N_9525);
and U9669 (N_9669,N_9462,N_9328);
nor U9670 (N_9670,N_9560,N_9533);
or U9671 (N_9671,N_9333,N_9336);
or U9672 (N_9672,N_9473,N_9499);
and U9673 (N_9673,N_9436,N_9392);
nand U9674 (N_9674,N_9325,N_9368);
xnor U9675 (N_9675,N_9356,N_9561);
xnor U9676 (N_9676,N_9542,N_9512);
nand U9677 (N_9677,N_9318,N_9309);
nor U9678 (N_9678,N_9572,N_9427);
xnor U9679 (N_9679,N_9414,N_9496);
and U9680 (N_9680,N_9515,N_9359);
nor U9681 (N_9681,N_9507,N_9411);
or U9682 (N_9682,N_9529,N_9308);
xnor U9683 (N_9683,N_9443,N_9316);
xnor U9684 (N_9684,N_9437,N_9597);
and U9685 (N_9685,N_9329,N_9432);
nand U9686 (N_9686,N_9554,N_9425);
and U9687 (N_9687,N_9590,N_9460);
or U9688 (N_9688,N_9478,N_9417);
and U9689 (N_9689,N_9435,N_9547);
and U9690 (N_9690,N_9377,N_9343);
or U9691 (N_9691,N_9466,N_9580);
or U9692 (N_9692,N_9522,N_9532);
nand U9693 (N_9693,N_9538,N_9511);
or U9694 (N_9694,N_9508,N_9408);
or U9695 (N_9695,N_9369,N_9354);
xor U9696 (N_9696,N_9489,N_9394);
nor U9697 (N_9697,N_9409,N_9416);
nor U9698 (N_9698,N_9404,N_9595);
xor U9699 (N_9699,N_9474,N_9480);
and U9700 (N_9700,N_9578,N_9433);
and U9701 (N_9701,N_9324,N_9301);
or U9702 (N_9702,N_9388,N_9594);
xor U9703 (N_9703,N_9583,N_9306);
and U9704 (N_9704,N_9319,N_9513);
or U9705 (N_9705,N_9571,N_9459);
and U9706 (N_9706,N_9444,N_9530);
and U9707 (N_9707,N_9472,N_9366);
and U9708 (N_9708,N_9387,N_9596);
nand U9709 (N_9709,N_9350,N_9463);
nand U9710 (N_9710,N_9389,N_9370);
nand U9711 (N_9711,N_9376,N_9576);
xnor U9712 (N_9712,N_9536,N_9348);
or U9713 (N_9713,N_9399,N_9320);
or U9714 (N_9714,N_9458,N_9300);
or U9715 (N_9715,N_9589,N_9500);
nand U9716 (N_9716,N_9440,N_9352);
and U9717 (N_9717,N_9506,N_9423);
and U9718 (N_9718,N_9396,N_9475);
nand U9719 (N_9719,N_9426,N_9526);
nand U9720 (N_9720,N_9591,N_9349);
nor U9721 (N_9721,N_9546,N_9510);
xnor U9722 (N_9722,N_9441,N_9593);
or U9723 (N_9723,N_9585,N_9375);
xor U9724 (N_9724,N_9599,N_9495);
nor U9725 (N_9725,N_9351,N_9567);
nor U9726 (N_9726,N_9461,N_9477);
xnor U9727 (N_9727,N_9311,N_9344);
and U9728 (N_9728,N_9555,N_9494);
nand U9729 (N_9729,N_9421,N_9493);
and U9730 (N_9730,N_9551,N_9535);
and U9731 (N_9731,N_9553,N_9490);
nand U9732 (N_9732,N_9341,N_9360);
xor U9733 (N_9733,N_9380,N_9429);
or U9734 (N_9734,N_9543,N_9457);
nand U9735 (N_9735,N_9312,N_9391);
nand U9736 (N_9736,N_9403,N_9381);
nand U9737 (N_9737,N_9581,N_9346);
and U9738 (N_9738,N_9374,N_9582);
xnor U9739 (N_9739,N_9556,N_9397);
nand U9740 (N_9740,N_9577,N_9541);
nor U9741 (N_9741,N_9479,N_9339);
nand U9742 (N_9742,N_9398,N_9367);
and U9743 (N_9743,N_9559,N_9355);
and U9744 (N_9744,N_9531,N_9430);
nand U9745 (N_9745,N_9385,N_9363);
nand U9746 (N_9746,N_9452,N_9415);
or U9747 (N_9747,N_9516,N_9406);
nand U9748 (N_9748,N_9401,N_9373);
or U9749 (N_9749,N_9305,N_9303);
or U9750 (N_9750,N_9304,N_9595);
and U9751 (N_9751,N_9436,N_9529);
nand U9752 (N_9752,N_9375,N_9557);
and U9753 (N_9753,N_9364,N_9555);
and U9754 (N_9754,N_9551,N_9562);
or U9755 (N_9755,N_9373,N_9415);
and U9756 (N_9756,N_9556,N_9386);
nand U9757 (N_9757,N_9313,N_9374);
xor U9758 (N_9758,N_9593,N_9374);
nor U9759 (N_9759,N_9421,N_9416);
or U9760 (N_9760,N_9529,N_9325);
and U9761 (N_9761,N_9472,N_9478);
xor U9762 (N_9762,N_9419,N_9370);
and U9763 (N_9763,N_9340,N_9336);
or U9764 (N_9764,N_9489,N_9548);
nor U9765 (N_9765,N_9570,N_9495);
nor U9766 (N_9766,N_9405,N_9319);
and U9767 (N_9767,N_9539,N_9561);
and U9768 (N_9768,N_9351,N_9375);
and U9769 (N_9769,N_9494,N_9437);
nand U9770 (N_9770,N_9358,N_9552);
and U9771 (N_9771,N_9301,N_9317);
and U9772 (N_9772,N_9442,N_9551);
and U9773 (N_9773,N_9584,N_9597);
nand U9774 (N_9774,N_9472,N_9374);
nor U9775 (N_9775,N_9333,N_9576);
nand U9776 (N_9776,N_9379,N_9360);
nor U9777 (N_9777,N_9380,N_9557);
and U9778 (N_9778,N_9364,N_9303);
nor U9779 (N_9779,N_9477,N_9409);
nand U9780 (N_9780,N_9597,N_9388);
or U9781 (N_9781,N_9459,N_9390);
nand U9782 (N_9782,N_9545,N_9411);
and U9783 (N_9783,N_9339,N_9516);
xnor U9784 (N_9784,N_9411,N_9587);
nand U9785 (N_9785,N_9310,N_9344);
or U9786 (N_9786,N_9568,N_9548);
xnor U9787 (N_9787,N_9535,N_9465);
nand U9788 (N_9788,N_9395,N_9524);
xor U9789 (N_9789,N_9546,N_9580);
and U9790 (N_9790,N_9357,N_9559);
and U9791 (N_9791,N_9396,N_9484);
or U9792 (N_9792,N_9488,N_9585);
nor U9793 (N_9793,N_9318,N_9432);
nor U9794 (N_9794,N_9329,N_9468);
or U9795 (N_9795,N_9597,N_9461);
nor U9796 (N_9796,N_9424,N_9392);
and U9797 (N_9797,N_9472,N_9340);
and U9798 (N_9798,N_9471,N_9570);
nor U9799 (N_9799,N_9405,N_9430);
nand U9800 (N_9800,N_9598,N_9502);
xor U9801 (N_9801,N_9426,N_9534);
nand U9802 (N_9802,N_9310,N_9548);
xnor U9803 (N_9803,N_9455,N_9461);
or U9804 (N_9804,N_9539,N_9410);
xor U9805 (N_9805,N_9591,N_9353);
or U9806 (N_9806,N_9522,N_9484);
and U9807 (N_9807,N_9434,N_9510);
and U9808 (N_9808,N_9520,N_9557);
xor U9809 (N_9809,N_9304,N_9577);
and U9810 (N_9810,N_9554,N_9367);
nand U9811 (N_9811,N_9508,N_9329);
or U9812 (N_9812,N_9598,N_9330);
nand U9813 (N_9813,N_9529,N_9460);
nand U9814 (N_9814,N_9369,N_9379);
nor U9815 (N_9815,N_9590,N_9323);
and U9816 (N_9816,N_9466,N_9596);
nand U9817 (N_9817,N_9417,N_9379);
nand U9818 (N_9818,N_9393,N_9322);
xnor U9819 (N_9819,N_9344,N_9536);
and U9820 (N_9820,N_9465,N_9392);
nor U9821 (N_9821,N_9356,N_9501);
nor U9822 (N_9822,N_9592,N_9423);
or U9823 (N_9823,N_9362,N_9564);
or U9824 (N_9824,N_9409,N_9410);
nand U9825 (N_9825,N_9555,N_9362);
nor U9826 (N_9826,N_9571,N_9584);
xnor U9827 (N_9827,N_9399,N_9502);
or U9828 (N_9828,N_9564,N_9532);
nand U9829 (N_9829,N_9599,N_9379);
or U9830 (N_9830,N_9529,N_9540);
nor U9831 (N_9831,N_9391,N_9528);
and U9832 (N_9832,N_9451,N_9324);
nand U9833 (N_9833,N_9543,N_9569);
and U9834 (N_9834,N_9590,N_9336);
xnor U9835 (N_9835,N_9479,N_9593);
nor U9836 (N_9836,N_9452,N_9405);
nand U9837 (N_9837,N_9482,N_9474);
or U9838 (N_9838,N_9392,N_9596);
nand U9839 (N_9839,N_9368,N_9324);
nand U9840 (N_9840,N_9386,N_9516);
nor U9841 (N_9841,N_9509,N_9313);
and U9842 (N_9842,N_9306,N_9327);
and U9843 (N_9843,N_9329,N_9433);
or U9844 (N_9844,N_9470,N_9521);
or U9845 (N_9845,N_9357,N_9528);
or U9846 (N_9846,N_9577,N_9391);
or U9847 (N_9847,N_9482,N_9333);
and U9848 (N_9848,N_9581,N_9558);
xnor U9849 (N_9849,N_9400,N_9329);
xor U9850 (N_9850,N_9302,N_9514);
or U9851 (N_9851,N_9305,N_9474);
xor U9852 (N_9852,N_9572,N_9548);
xnor U9853 (N_9853,N_9491,N_9479);
or U9854 (N_9854,N_9380,N_9457);
xnor U9855 (N_9855,N_9426,N_9550);
and U9856 (N_9856,N_9365,N_9302);
nand U9857 (N_9857,N_9323,N_9426);
nor U9858 (N_9858,N_9589,N_9300);
xor U9859 (N_9859,N_9507,N_9550);
nand U9860 (N_9860,N_9430,N_9424);
or U9861 (N_9861,N_9370,N_9560);
and U9862 (N_9862,N_9477,N_9595);
xnor U9863 (N_9863,N_9368,N_9308);
xnor U9864 (N_9864,N_9551,N_9582);
nor U9865 (N_9865,N_9563,N_9531);
and U9866 (N_9866,N_9383,N_9479);
xor U9867 (N_9867,N_9408,N_9512);
nor U9868 (N_9868,N_9420,N_9445);
or U9869 (N_9869,N_9497,N_9533);
and U9870 (N_9870,N_9401,N_9526);
or U9871 (N_9871,N_9595,N_9337);
and U9872 (N_9872,N_9451,N_9507);
xnor U9873 (N_9873,N_9478,N_9411);
nor U9874 (N_9874,N_9365,N_9358);
nand U9875 (N_9875,N_9597,N_9520);
nand U9876 (N_9876,N_9547,N_9510);
nor U9877 (N_9877,N_9464,N_9415);
and U9878 (N_9878,N_9503,N_9395);
xor U9879 (N_9879,N_9556,N_9365);
and U9880 (N_9880,N_9494,N_9582);
nand U9881 (N_9881,N_9372,N_9304);
and U9882 (N_9882,N_9346,N_9302);
and U9883 (N_9883,N_9433,N_9454);
and U9884 (N_9884,N_9319,N_9420);
or U9885 (N_9885,N_9438,N_9368);
xor U9886 (N_9886,N_9380,N_9482);
or U9887 (N_9887,N_9361,N_9420);
nand U9888 (N_9888,N_9469,N_9305);
nor U9889 (N_9889,N_9591,N_9590);
or U9890 (N_9890,N_9542,N_9395);
xor U9891 (N_9891,N_9319,N_9587);
or U9892 (N_9892,N_9456,N_9440);
and U9893 (N_9893,N_9485,N_9329);
nand U9894 (N_9894,N_9343,N_9322);
xor U9895 (N_9895,N_9498,N_9387);
nand U9896 (N_9896,N_9474,N_9331);
or U9897 (N_9897,N_9527,N_9499);
nand U9898 (N_9898,N_9450,N_9439);
nor U9899 (N_9899,N_9394,N_9558);
or U9900 (N_9900,N_9806,N_9720);
nor U9901 (N_9901,N_9781,N_9654);
nand U9902 (N_9902,N_9602,N_9621);
nand U9903 (N_9903,N_9729,N_9872);
nand U9904 (N_9904,N_9680,N_9627);
and U9905 (N_9905,N_9681,N_9874);
nor U9906 (N_9906,N_9869,N_9657);
and U9907 (N_9907,N_9826,N_9718);
or U9908 (N_9908,N_9810,N_9619);
xnor U9909 (N_9909,N_9883,N_9618);
nand U9910 (N_9910,N_9751,N_9867);
nand U9911 (N_9911,N_9827,N_9802);
and U9912 (N_9912,N_9835,N_9607);
or U9913 (N_9913,N_9811,N_9648);
or U9914 (N_9914,N_9812,N_9818);
or U9915 (N_9915,N_9755,N_9773);
nand U9916 (N_9916,N_9899,N_9660);
and U9917 (N_9917,N_9787,N_9875);
or U9918 (N_9918,N_9622,N_9858);
or U9919 (N_9919,N_9888,N_9746);
and U9920 (N_9920,N_9739,N_9682);
nand U9921 (N_9921,N_9647,N_9713);
and U9922 (N_9922,N_9631,N_9757);
or U9923 (N_9923,N_9782,N_9700);
xor U9924 (N_9924,N_9662,N_9674);
nor U9925 (N_9925,N_9603,N_9701);
or U9926 (N_9926,N_9889,N_9708);
or U9927 (N_9927,N_9721,N_9873);
or U9928 (N_9928,N_9877,N_9849);
nor U9929 (N_9929,N_9897,N_9684);
nor U9930 (N_9930,N_9679,N_9742);
nor U9931 (N_9931,N_9853,N_9797);
or U9932 (N_9932,N_9691,N_9604);
nor U9933 (N_9933,N_9821,N_9860);
xnor U9934 (N_9934,N_9642,N_9846);
nor U9935 (N_9935,N_9832,N_9756);
and U9936 (N_9936,N_9633,N_9879);
nor U9937 (N_9937,N_9666,N_9809);
nand U9938 (N_9938,N_9876,N_9763);
or U9939 (N_9939,N_9683,N_9878);
nor U9940 (N_9940,N_9722,N_9606);
nor U9941 (N_9941,N_9749,N_9840);
xnor U9942 (N_9942,N_9772,N_9778);
nor U9943 (N_9943,N_9706,N_9789);
nor U9944 (N_9944,N_9791,N_9608);
nor U9945 (N_9945,N_9712,N_9779);
nand U9946 (N_9946,N_9637,N_9824);
xnor U9947 (N_9947,N_9898,N_9696);
or U9948 (N_9948,N_9850,N_9728);
nand U9949 (N_9949,N_9752,N_9732);
or U9950 (N_9950,N_9687,N_9833);
nand U9951 (N_9951,N_9842,N_9725);
xor U9952 (N_9952,N_9704,N_9645);
or U9953 (N_9953,N_9766,N_9675);
and U9954 (N_9954,N_9617,N_9776);
nand U9955 (N_9955,N_9774,N_9890);
or U9956 (N_9956,N_9671,N_9771);
nor U9957 (N_9957,N_9887,N_9893);
or U9958 (N_9958,N_9768,N_9765);
nor U9959 (N_9959,N_9726,N_9616);
nor U9960 (N_9960,N_9646,N_9839);
or U9961 (N_9961,N_9609,N_9730);
xor U9962 (N_9962,N_9624,N_9620);
and U9963 (N_9963,N_9894,N_9798);
nand U9964 (N_9964,N_9881,N_9868);
nand U9965 (N_9965,N_9834,N_9688);
xnor U9966 (N_9966,N_9717,N_9855);
and U9967 (N_9967,N_9822,N_9856);
nor U9968 (N_9968,N_9817,N_9828);
and U9969 (N_9969,N_9775,N_9611);
nor U9970 (N_9970,N_9767,N_9814);
nand U9971 (N_9971,N_9659,N_9851);
xnor U9972 (N_9972,N_9692,N_9673);
or U9973 (N_9973,N_9885,N_9644);
xor U9974 (N_9974,N_9769,N_9747);
or U9975 (N_9975,N_9841,N_9760);
nor U9976 (N_9976,N_9629,N_9678);
and U9977 (N_9977,N_9805,N_9650);
or U9978 (N_9978,N_9823,N_9825);
nand U9979 (N_9979,N_9643,N_9723);
or U9980 (N_9980,N_9649,N_9784);
and U9981 (N_9981,N_9697,N_9731);
xor U9982 (N_9982,N_9702,N_9820);
nand U9983 (N_9983,N_9754,N_9830);
and U9984 (N_9984,N_9735,N_9777);
nor U9985 (N_9985,N_9785,N_9790);
xor U9986 (N_9986,N_9625,N_9896);
or U9987 (N_9987,N_9663,N_9891);
nor U9988 (N_9988,N_9669,N_9819);
nand U9989 (N_9989,N_9800,N_9623);
nor U9990 (N_9990,N_9614,N_9750);
xor U9991 (N_9991,N_9610,N_9848);
nor U9992 (N_9992,N_9711,N_9753);
and U9993 (N_9993,N_9719,N_9799);
or U9994 (N_9994,N_9761,N_9698);
and U9995 (N_9995,N_9600,N_9656);
or U9996 (N_9996,N_9852,N_9804);
nor U9997 (N_9997,N_9664,N_9738);
or U9998 (N_9998,N_9714,N_9759);
xnor U9999 (N_9999,N_9892,N_9831);
and U10000 (N_10000,N_9686,N_9745);
or U10001 (N_10001,N_9859,N_9737);
nand U10002 (N_10002,N_9667,N_9715);
nand U10003 (N_10003,N_9668,N_9676);
and U10004 (N_10004,N_9863,N_9634);
nor U10005 (N_10005,N_9640,N_9808);
nor U10006 (N_10006,N_9854,N_9727);
xnor U10007 (N_10007,N_9792,N_9685);
xnor U10008 (N_10008,N_9838,N_9635);
nand U10009 (N_10009,N_9628,N_9709);
nand U10010 (N_10010,N_9794,N_9864);
or U10011 (N_10011,N_9845,N_9880);
or U10012 (N_10012,N_9707,N_9882);
xor U10013 (N_10013,N_9612,N_9801);
xnor U10014 (N_10014,N_9886,N_9651);
nor U10015 (N_10015,N_9716,N_9693);
or U10016 (N_10016,N_9615,N_9703);
nand U10017 (N_10017,N_9843,N_9870);
or U10018 (N_10018,N_9857,N_9748);
xor U10019 (N_10019,N_9672,N_9670);
nor U10020 (N_10020,N_9665,N_9639);
nor U10021 (N_10021,N_9744,N_9652);
nor U10022 (N_10022,N_9795,N_9783);
nand U10023 (N_10023,N_9694,N_9895);
or U10024 (N_10024,N_9689,N_9638);
nand U10025 (N_10025,N_9695,N_9605);
nor U10026 (N_10026,N_9630,N_9803);
nand U10027 (N_10027,N_9788,N_9758);
or U10028 (N_10028,N_9641,N_9743);
nor U10029 (N_10029,N_9871,N_9865);
and U10030 (N_10030,N_9813,N_9632);
nand U10031 (N_10031,N_9653,N_9636);
nor U10032 (N_10032,N_9793,N_9780);
and U10033 (N_10033,N_9740,N_9847);
nor U10034 (N_10034,N_9661,N_9862);
xor U10035 (N_10035,N_9613,N_9866);
nand U10036 (N_10036,N_9815,N_9741);
nor U10037 (N_10037,N_9724,N_9733);
xnor U10038 (N_10038,N_9677,N_9861);
or U10039 (N_10039,N_9626,N_9658);
nand U10040 (N_10040,N_9705,N_9770);
nor U10041 (N_10041,N_9816,N_9710);
nand U10042 (N_10042,N_9601,N_9734);
nand U10043 (N_10043,N_9844,N_9836);
or U10044 (N_10044,N_9796,N_9786);
nor U10045 (N_10045,N_9807,N_9829);
xor U10046 (N_10046,N_9690,N_9655);
or U10047 (N_10047,N_9762,N_9736);
xor U10048 (N_10048,N_9837,N_9884);
nand U10049 (N_10049,N_9699,N_9764);
and U10050 (N_10050,N_9627,N_9890);
nand U10051 (N_10051,N_9836,N_9602);
nand U10052 (N_10052,N_9799,N_9673);
nand U10053 (N_10053,N_9796,N_9888);
nor U10054 (N_10054,N_9873,N_9821);
nand U10055 (N_10055,N_9759,N_9847);
or U10056 (N_10056,N_9660,N_9896);
nor U10057 (N_10057,N_9701,N_9780);
nand U10058 (N_10058,N_9632,N_9816);
or U10059 (N_10059,N_9662,N_9695);
or U10060 (N_10060,N_9639,N_9845);
or U10061 (N_10061,N_9737,N_9776);
xnor U10062 (N_10062,N_9647,N_9886);
xor U10063 (N_10063,N_9786,N_9821);
and U10064 (N_10064,N_9706,N_9784);
and U10065 (N_10065,N_9795,N_9687);
and U10066 (N_10066,N_9671,N_9759);
or U10067 (N_10067,N_9771,N_9885);
nor U10068 (N_10068,N_9715,N_9882);
and U10069 (N_10069,N_9656,N_9690);
or U10070 (N_10070,N_9644,N_9894);
nor U10071 (N_10071,N_9782,N_9726);
nand U10072 (N_10072,N_9836,N_9815);
or U10073 (N_10073,N_9709,N_9760);
nand U10074 (N_10074,N_9643,N_9684);
nor U10075 (N_10075,N_9838,N_9663);
or U10076 (N_10076,N_9757,N_9781);
xor U10077 (N_10077,N_9763,N_9607);
or U10078 (N_10078,N_9664,N_9749);
nor U10079 (N_10079,N_9635,N_9717);
and U10080 (N_10080,N_9780,N_9748);
nor U10081 (N_10081,N_9778,N_9677);
nor U10082 (N_10082,N_9774,N_9819);
nor U10083 (N_10083,N_9658,N_9809);
and U10084 (N_10084,N_9729,N_9697);
nand U10085 (N_10085,N_9631,N_9751);
and U10086 (N_10086,N_9817,N_9616);
xnor U10087 (N_10087,N_9664,N_9886);
nor U10088 (N_10088,N_9815,N_9899);
or U10089 (N_10089,N_9811,N_9768);
nor U10090 (N_10090,N_9672,N_9705);
nor U10091 (N_10091,N_9745,N_9880);
xnor U10092 (N_10092,N_9728,N_9803);
nor U10093 (N_10093,N_9692,N_9799);
and U10094 (N_10094,N_9737,N_9674);
nand U10095 (N_10095,N_9748,N_9779);
and U10096 (N_10096,N_9723,N_9787);
or U10097 (N_10097,N_9855,N_9695);
or U10098 (N_10098,N_9871,N_9699);
nor U10099 (N_10099,N_9827,N_9647);
nor U10100 (N_10100,N_9761,N_9779);
nand U10101 (N_10101,N_9617,N_9879);
or U10102 (N_10102,N_9745,N_9810);
or U10103 (N_10103,N_9784,N_9818);
xor U10104 (N_10104,N_9793,N_9618);
nor U10105 (N_10105,N_9687,N_9890);
nor U10106 (N_10106,N_9636,N_9659);
xnor U10107 (N_10107,N_9813,N_9809);
nand U10108 (N_10108,N_9759,N_9889);
nor U10109 (N_10109,N_9724,N_9845);
and U10110 (N_10110,N_9646,N_9812);
nor U10111 (N_10111,N_9645,N_9636);
xor U10112 (N_10112,N_9844,N_9804);
nor U10113 (N_10113,N_9772,N_9654);
and U10114 (N_10114,N_9634,N_9800);
and U10115 (N_10115,N_9646,N_9671);
nand U10116 (N_10116,N_9813,N_9886);
xor U10117 (N_10117,N_9836,N_9811);
or U10118 (N_10118,N_9810,N_9809);
and U10119 (N_10119,N_9808,N_9675);
or U10120 (N_10120,N_9738,N_9625);
and U10121 (N_10121,N_9621,N_9795);
nor U10122 (N_10122,N_9652,N_9660);
nor U10123 (N_10123,N_9802,N_9684);
or U10124 (N_10124,N_9897,N_9723);
xnor U10125 (N_10125,N_9684,N_9872);
xor U10126 (N_10126,N_9677,N_9736);
nand U10127 (N_10127,N_9635,N_9700);
nor U10128 (N_10128,N_9731,N_9784);
xnor U10129 (N_10129,N_9835,N_9829);
xnor U10130 (N_10130,N_9708,N_9764);
nor U10131 (N_10131,N_9887,N_9736);
or U10132 (N_10132,N_9650,N_9632);
nand U10133 (N_10133,N_9799,N_9894);
and U10134 (N_10134,N_9852,N_9645);
or U10135 (N_10135,N_9853,N_9889);
nand U10136 (N_10136,N_9840,N_9872);
nand U10137 (N_10137,N_9639,N_9745);
xnor U10138 (N_10138,N_9773,N_9810);
nor U10139 (N_10139,N_9678,N_9709);
xor U10140 (N_10140,N_9884,N_9612);
and U10141 (N_10141,N_9772,N_9638);
nand U10142 (N_10142,N_9682,N_9681);
nand U10143 (N_10143,N_9848,N_9810);
and U10144 (N_10144,N_9662,N_9796);
nand U10145 (N_10145,N_9664,N_9682);
and U10146 (N_10146,N_9626,N_9701);
or U10147 (N_10147,N_9749,N_9697);
nor U10148 (N_10148,N_9738,N_9644);
and U10149 (N_10149,N_9726,N_9679);
xnor U10150 (N_10150,N_9652,N_9686);
or U10151 (N_10151,N_9826,N_9691);
nor U10152 (N_10152,N_9807,N_9682);
or U10153 (N_10153,N_9734,N_9887);
nor U10154 (N_10154,N_9840,N_9877);
xor U10155 (N_10155,N_9711,N_9821);
nand U10156 (N_10156,N_9609,N_9694);
nand U10157 (N_10157,N_9716,N_9835);
xor U10158 (N_10158,N_9663,N_9745);
nor U10159 (N_10159,N_9751,N_9807);
nand U10160 (N_10160,N_9868,N_9875);
or U10161 (N_10161,N_9630,N_9804);
nand U10162 (N_10162,N_9603,N_9767);
xnor U10163 (N_10163,N_9811,N_9664);
nor U10164 (N_10164,N_9832,N_9781);
or U10165 (N_10165,N_9816,N_9883);
or U10166 (N_10166,N_9778,N_9866);
nand U10167 (N_10167,N_9839,N_9722);
nor U10168 (N_10168,N_9691,N_9661);
nand U10169 (N_10169,N_9745,N_9854);
nand U10170 (N_10170,N_9867,N_9821);
or U10171 (N_10171,N_9763,N_9712);
nor U10172 (N_10172,N_9839,N_9693);
xor U10173 (N_10173,N_9898,N_9812);
or U10174 (N_10174,N_9754,N_9604);
nor U10175 (N_10175,N_9737,N_9768);
and U10176 (N_10176,N_9740,N_9683);
and U10177 (N_10177,N_9747,N_9745);
nand U10178 (N_10178,N_9680,N_9865);
nand U10179 (N_10179,N_9872,N_9725);
and U10180 (N_10180,N_9830,N_9633);
or U10181 (N_10181,N_9894,N_9811);
or U10182 (N_10182,N_9809,N_9700);
xor U10183 (N_10183,N_9775,N_9632);
or U10184 (N_10184,N_9824,N_9615);
nand U10185 (N_10185,N_9603,N_9795);
xor U10186 (N_10186,N_9819,N_9899);
and U10187 (N_10187,N_9849,N_9639);
xnor U10188 (N_10188,N_9750,N_9735);
xor U10189 (N_10189,N_9746,N_9739);
nand U10190 (N_10190,N_9731,N_9820);
nand U10191 (N_10191,N_9844,N_9742);
nand U10192 (N_10192,N_9723,N_9861);
or U10193 (N_10193,N_9775,N_9742);
xnor U10194 (N_10194,N_9752,N_9884);
and U10195 (N_10195,N_9770,N_9680);
nand U10196 (N_10196,N_9783,N_9832);
nor U10197 (N_10197,N_9704,N_9710);
or U10198 (N_10198,N_9826,N_9897);
nor U10199 (N_10199,N_9811,N_9765);
nand U10200 (N_10200,N_10121,N_10083);
or U10201 (N_10201,N_10140,N_10127);
xnor U10202 (N_10202,N_9917,N_9947);
nor U10203 (N_10203,N_10177,N_10053);
nand U10204 (N_10204,N_9919,N_10014);
or U10205 (N_10205,N_10024,N_10156);
xor U10206 (N_10206,N_10038,N_10139);
nand U10207 (N_10207,N_9937,N_9991);
xnor U10208 (N_10208,N_10176,N_10187);
nand U10209 (N_10209,N_10167,N_9972);
xnor U10210 (N_10210,N_10085,N_10133);
xor U10211 (N_10211,N_10065,N_10044);
nor U10212 (N_10212,N_10021,N_9964);
or U10213 (N_10213,N_9990,N_10166);
nand U10214 (N_10214,N_10050,N_9946);
nor U10215 (N_10215,N_10143,N_9995);
nor U10216 (N_10216,N_9989,N_9963);
nor U10217 (N_10217,N_10054,N_10055);
xor U10218 (N_10218,N_9904,N_10049);
nand U10219 (N_10219,N_10040,N_10197);
nor U10220 (N_10220,N_9936,N_9997);
nand U10221 (N_10221,N_9986,N_10154);
nand U10222 (N_10222,N_10094,N_9978);
nor U10223 (N_10223,N_9902,N_10129);
and U10224 (N_10224,N_10060,N_10070);
or U10225 (N_10225,N_10087,N_10198);
nor U10226 (N_10226,N_10010,N_10191);
and U10227 (N_10227,N_9925,N_10086);
nor U10228 (N_10228,N_10036,N_9970);
or U10229 (N_10229,N_9903,N_10150);
xnor U10230 (N_10230,N_10076,N_10131);
nand U10231 (N_10231,N_9958,N_10062);
xnor U10232 (N_10232,N_10093,N_9907);
or U10233 (N_10233,N_9980,N_10001);
xnor U10234 (N_10234,N_10162,N_10046);
nand U10235 (N_10235,N_10136,N_10034);
xnor U10236 (N_10236,N_9954,N_10102);
or U10237 (N_10237,N_10068,N_9967);
and U10238 (N_10238,N_10193,N_10137);
nor U10239 (N_10239,N_9996,N_10020);
and U10240 (N_10240,N_9938,N_10132);
or U10241 (N_10241,N_10059,N_9924);
nand U10242 (N_10242,N_10158,N_10116);
or U10243 (N_10243,N_10066,N_9935);
nand U10244 (N_10244,N_10023,N_9953);
nand U10245 (N_10245,N_9960,N_10035);
nor U10246 (N_10246,N_9928,N_10006);
nand U10247 (N_10247,N_10032,N_10003);
or U10248 (N_10248,N_10141,N_10189);
nand U10249 (N_10249,N_10153,N_10015);
nor U10250 (N_10250,N_10002,N_10027);
or U10251 (N_10251,N_10179,N_9944);
nor U10252 (N_10252,N_9971,N_10120);
xor U10253 (N_10253,N_10045,N_10199);
xor U10254 (N_10254,N_9920,N_10122);
or U10255 (N_10255,N_9932,N_9942);
and U10256 (N_10256,N_10170,N_10125);
nand U10257 (N_10257,N_10119,N_10090);
nor U10258 (N_10258,N_10134,N_10042);
nand U10259 (N_10259,N_10145,N_9941);
or U10260 (N_10260,N_9968,N_10175);
xor U10261 (N_10261,N_9984,N_10089);
nand U10262 (N_10262,N_9922,N_9927);
nand U10263 (N_10263,N_10097,N_10067);
nand U10264 (N_10264,N_10112,N_10004);
nand U10265 (N_10265,N_9988,N_9987);
and U10266 (N_10266,N_10165,N_9952);
nor U10267 (N_10267,N_10123,N_9999);
xor U10268 (N_10268,N_9966,N_10009);
or U10269 (N_10269,N_9961,N_9905);
nor U10270 (N_10270,N_10181,N_10157);
nand U10271 (N_10271,N_9985,N_10180);
xor U10272 (N_10272,N_10168,N_10071);
nor U10273 (N_10273,N_10100,N_10106);
or U10274 (N_10274,N_10057,N_9949);
or U10275 (N_10275,N_10016,N_10194);
xnor U10276 (N_10276,N_9913,N_10185);
nand U10277 (N_10277,N_9992,N_10000);
xor U10278 (N_10278,N_10135,N_10118);
and U10279 (N_10279,N_10190,N_10064);
and U10280 (N_10280,N_9950,N_10149);
or U10281 (N_10281,N_10161,N_10029);
nand U10282 (N_10282,N_10113,N_10084);
nor U10283 (N_10283,N_9945,N_10017);
or U10284 (N_10284,N_10103,N_10026);
and U10285 (N_10285,N_9948,N_10078);
nor U10286 (N_10286,N_9933,N_9957);
or U10287 (N_10287,N_10098,N_9915);
nor U10288 (N_10288,N_10186,N_10108);
nor U10289 (N_10289,N_10144,N_10095);
or U10290 (N_10290,N_10183,N_10048);
xor U10291 (N_10291,N_9979,N_9969);
nor U10292 (N_10292,N_10013,N_10148);
and U10293 (N_10293,N_10081,N_10072);
or U10294 (N_10294,N_10130,N_10043);
nand U10295 (N_10295,N_10110,N_10164);
xor U10296 (N_10296,N_9910,N_9981);
and U10297 (N_10297,N_10160,N_10138);
and U10298 (N_10298,N_9916,N_10041);
nand U10299 (N_10299,N_9976,N_10088);
xnor U10300 (N_10300,N_10056,N_10092);
nor U10301 (N_10301,N_10058,N_10174);
xor U10302 (N_10302,N_9931,N_9901);
xor U10303 (N_10303,N_10128,N_10028);
nor U10304 (N_10304,N_9974,N_10114);
xor U10305 (N_10305,N_10047,N_10079);
xor U10306 (N_10306,N_10159,N_9923);
or U10307 (N_10307,N_9951,N_10061);
nor U10308 (N_10308,N_10151,N_10091);
nand U10309 (N_10309,N_9918,N_9940);
or U10310 (N_10310,N_10051,N_10008);
xor U10311 (N_10311,N_9982,N_9962);
and U10312 (N_10312,N_10005,N_10052);
and U10313 (N_10313,N_10196,N_9911);
nor U10314 (N_10314,N_9929,N_10096);
or U10315 (N_10315,N_10074,N_9908);
nand U10316 (N_10316,N_10037,N_10011);
or U10317 (N_10317,N_10155,N_10031);
or U10318 (N_10318,N_9914,N_10107);
nor U10319 (N_10319,N_10195,N_9993);
nor U10320 (N_10320,N_10109,N_10188);
nand U10321 (N_10321,N_10104,N_9998);
xnor U10322 (N_10322,N_10030,N_9977);
nor U10323 (N_10323,N_9959,N_10172);
xor U10324 (N_10324,N_10022,N_9975);
or U10325 (N_10325,N_10018,N_10069);
or U10326 (N_10326,N_10152,N_10073);
and U10327 (N_10327,N_10192,N_9930);
and U10328 (N_10328,N_9965,N_10163);
nor U10329 (N_10329,N_9956,N_10099);
xnor U10330 (N_10330,N_9939,N_9909);
nand U10331 (N_10331,N_9906,N_10063);
nand U10332 (N_10332,N_10075,N_10101);
xnor U10333 (N_10333,N_9973,N_10012);
nand U10334 (N_10334,N_10019,N_9983);
or U10335 (N_10335,N_9934,N_10105);
and U10336 (N_10336,N_10126,N_10182);
nor U10337 (N_10337,N_9943,N_10173);
and U10338 (N_10338,N_10080,N_9912);
nor U10339 (N_10339,N_10111,N_10082);
xor U10340 (N_10340,N_9955,N_10169);
nand U10341 (N_10341,N_10007,N_10124);
nor U10342 (N_10342,N_10033,N_10077);
or U10343 (N_10343,N_10171,N_9926);
and U10344 (N_10344,N_10142,N_9900);
and U10345 (N_10345,N_9994,N_10039);
nand U10346 (N_10346,N_10147,N_10115);
or U10347 (N_10347,N_10117,N_10146);
or U10348 (N_10348,N_9921,N_10025);
nor U10349 (N_10349,N_10178,N_10184);
nor U10350 (N_10350,N_9926,N_10176);
xnor U10351 (N_10351,N_9920,N_10069);
nand U10352 (N_10352,N_10196,N_9985);
xnor U10353 (N_10353,N_10114,N_9943);
or U10354 (N_10354,N_10033,N_9968);
xor U10355 (N_10355,N_10146,N_10094);
nand U10356 (N_10356,N_10043,N_10184);
and U10357 (N_10357,N_9964,N_10046);
or U10358 (N_10358,N_9954,N_10073);
nor U10359 (N_10359,N_9926,N_10165);
xor U10360 (N_10360,N_10006,N_10056);
nor U10361 (N_10361,N_10004,N_10013);
and U10362 (N_10362,N_10166,N_10084);
or U10363 (N_10363,N_10165,N_10110);
xnor U10364 (N_10364,N_9976,N_10194);
nor U10365 (N_10365,N_10051,N_10157);
or U10366 (N_10366,N_10066,N_10181);
nor U10367 (N_10367,N_10045,N_10103);
nor U10368 (N_10368,N_10150,N_9995);
nor U10369 (N_10369,N_9919,N_9921);
or U10370 (N_10370,N_9976,N_10132);
nand U10371 (N_10371,N_9988,N_10184);
or U10372 (N_10372,N_9981,N_9930);
or U10373 (N_10373,N_9931,N_10118);
and U10374 (N_10374,N_9983,N_10080);
and U10375 (N_10375,N_10082,N_10049);
xnor U10376 (N_10376,N_10102,N_10163);
nand U10377 (N_10377,N_10006,N_10149);
xnor U10378 (N_10378,N_10099,N_9910);
or U10379 (N_10379,N_10077,N_10133);
or U10380 (N_10380,N_10074,N_10063);
xor U10381 (N_10381,N_10001,N_10198);
nor U10382 (N_10382,N_10167,N_10129);
or U10383 (N_10383,N_10185,N_10101);
or U10384 (N_10384,N_10130,N_10107);
nor U10385 (N_10385,N_10188,N_9923);
and U10386 (N_10386,N_10002,N_10192);
xnor U10387 (N_10387,N_10190,N_9969);
xnor U10388 (N_10388,N_9954,N_10132);
nor U10389 (N_10389,N_9900,N_10054);
nor U10390 (N_10390,N_10120,N_9989);
xor U10391 (N_10391,N_9953,N_9996);
and U10392 (N_10392,N_10193,N_10149);
xor U10393 (N_10393,N_9917,N_10117);
or U10394 (N_10394,N_9970,N_9967);
or U10395 (N_10395,N_10075,N_10063);
nor U10396 (N_10396,N_9925,N_10182);
and U10397 (N_10397,N_9945,N_9990);
and U10398 (N_10398,N_9948,N_10044);
nand U10399 (N_10399,N_10023,N_10155);
nor U10400 (N_10400,N_10048,N_10054);
and U10401 (N_10401,N_10103,N_10152);
nand U10402 (N_10402,N_9974,N_10141);
or U10403 (N_10403,N_9984,N_9974);
nand U10404 (N_10404,N_10014,N_10106);
nand U10405 (N_10405,N_10173,N_10192);
and U10406 (N_10406,N_9967,N_10126);
and U10407 (N_10407,N_9949,N_10107);
and U10408 (N_10408,N_10055,N_10003);
nand U10409 (N_10409,N_10127,N_9908);
or U10410 (N_10410,N_10179,N_9945);
nand U10411 (N_10411,N_9962,N_9980);
and U10412 (N_10412,N_10134,N_10198);
or U10413 (N_10413,N_10053,N_10063);
xor U10414 (N_10414,N_10144,N_10034);
or U10415 (N_10415,N_9913,N_10014);
xor U10416 (N_10416,N_9926,N_10081);
or U10417 (N_10417,N_9968,N_9981);
nand U10418 (N_10418,N_9956,N_10191);
nand U10419 (N_10419,N_10026,N_10193);
or U10420 (N_10420,N_10056,N_9902);
nand U10421 (N_10421,N_10047,N_10030);
nor U10422 (N_10422,N_10087,N_10060);
nand U10423 (N_10423,N_9911,N_9913);
and U10424 (N_10424,N_10193,N_10116);
nor U10425 (N_10425,N_9967,N_10135);
or U10426 (N_10426,N_10069,N_10057);
and U10427 (N_10427,N_10172,N_10054);
xnor U10428 (N_10428,N_10170,N_9971);
nor U10429 (N_10429,N_9907,N_10036);
nor U10430 (N_10430,N_10049,N_10012);
xor U10431 (N_10431,N_10012,N_10032);
or U10432 (N_10432,N_10177,N_10199);
xnor U10433 (N_10433,N_10122,N_10051);
or U10434 (N_10434,N_10089,N_10057);
xnor U10435 (N_10435,N_9947,N_10097);
nand U10436 (N_10436,N_10014,N_10052);
xnor U10437 (N_10437,N_10184,N_10174);
and U10438 (N_10438,N_10016,N_10191);
and U10439 (N_10439,N_10191,N_9900);
and U10440 (N_10440,N_10047,N_9970);
nand U10441 (N_10441,N_10091,N_10046);
nand U10442 (N_10442,N_9954,N_10095);
nor U10443 (N_10443,N_9966,N_10096);
or U10444 (N_10444,N_10082,N_10137);
or U10445 (N_10445,N_9925,N_10171);
xor U10446 (N_10446,N_10003,N_10199);
or U10447 (N_10447,N_10120,N_10113);
nand U10448 (N_10448,N_10126,N_9986);
nand U10449 (N_10449,N_10191,N_9931);
nand U10450 (N_10450,N_10048,N_10017);
nand U10451 (N_10451,N_10098,N_9952);
nor U10452 (N_10452,N_10169,N_9917);
xnor U10453 (N_10453,N_9966,N_9990);
and U10454 (N_10454,N_10131,N_10165);
or U10455 (N_10455,N_10112,N_10025);
xnor U10456 (N_10456,N_10041,N_9934);
nor U10457 (N_10457,N_9962,N_10138);
xnor U10458 (N_10458,N_10143,N_10100);
xnor U10459 (N_10459,N_9938,N_10136);
or U10460 (N_10460,N_10176,N_10046);
and U10461 (N_10461,N_9979,N_9985);
xnor U10462 (N_10462,N_9972,N_10149);
xnor U10463 (N_10463,N_10089,N_9979);
nor U10464 (N_10464,N_10101,N_9941);
xnor U10465 (N_10465,N_10059,N_9984);
and U10466 (N_10466,N_10094,N_10023);
nand U10467 (N_10467,N_9945,N_10158);
nand U10468 (N_10468,N_9985,N_10019);
xnor U10469 (N_10469,N_10192,N_10140);
xnor U10470 (N_10470,N_10124,N_10019);
and U10471 (N_10471,N_9913,N_9901);
xor U10472 (N_10472,N_9984,N_9921);
xnor U10473 (N_10473,N_9996,N_10175);
and U10474 (N_10474,N_10036,N_10177);
and U10475 (N_10475,N_9937,N_10038);
nor U10476 (N_10476,N_10199,N_10001);
xor U10477 (N_10477,N_10130,N_9976);
nand U10478 (N_10478,N_10176,N_10011);
or U10479 (N_10479,N_10036,N_10140);
or U10480 (N_10480,N_10122,N_10084);
and U10481 (N_10481,N_10025,N_10152);
nor U10482 (N_10482,N_9947,N_10185);
and U10483 (N_10483,N_10145,N_10175);
nor U10484 (N_10484,N_10057,N_9952);
xnor U10485 (N_10485,N_10024,N_9924);
or U10486 (N_10486,N_10140,N_10156);
nor U10487 (N_10487,N_10187,N_9990);
nand U10488 (N_10488,N_10187,N_9957);
or U10489 (N_10489,N_10122,N_9967);
nor U10490 (N_10490,N_10126,N_10165);
nor U10491 (N_10491,N_10072,N_9957);
and U10492 (N_10492,N_9937,N_10074);
or U10493 (N_10493,N_9984,N_9933);
xor U10494 (N_10494,N_9977,N_10047);
nand U10495 (N_10495,N_10182,N_10107);
nand U10496 (N_10496,N_10095,N_10122);
nor U10497 (N_10497,N_10119,N_10129);
nand U10498 (N_10498,N_10115,N_10117);
nor U10499 (N_10499,N_10010,N_10038);
and U10500 (N_10500,N_10331,N_10434);
nor U10501 (N_10501,N_10394,N_10294);
nand U10502 (N_10502,N_10412,N_10232);
nor U10503 (N_10503,N_10417,N_10353);
nand U10504 (N_10504,N_10268,N_10439);
xnor U10505 (N_10505,N_10465,N_10222);
or U10506 (N_10506,N_10468,N_10457);
nand U10507 (N_10507,N_10459,N_10399);
and U10508 (N_10508,N_10273,N_10248);
or U10509 (N_10509,N_10435,N_10244);
nand U10510 (N_10510,N_10471,N_10321);
xor U10511 (N_10511,N_10252,N_10253);
and U10512 (N_10512,N_10343,N_10396);
xor U10513 (N_10513,N_10267,N_10272);
or U10514 (N_10514,N_10354,N_10256);
or U10515 (N_10515,N_10275,N_10236);
and U10516 (N_10516,N_10350,N_10372);
or U10517 (N_10517,N_10277,N_10442);
and U10518 (N_10518,N_10328,N_10498);
nor U10519 (N_10519,N_10438,N_10488);
and U10520 (N_10520,N_10373,N_10473);
and U10521 (N_10521,N_10274,N_10392);
or U10522 (N_10522,N_10271,N_10255);
or U10523 (N_10523,N_10241,N_10458);
nor U10524 (N_10524,N_10299,N_10485);
nand U10525 (N_10525,N_10254,N_10482);
and U10526 (N_10526,N_10213,N_10289);
nand U10527 (N_10527,N_10344,N_10281);
nor U10528 (N_10528,N_10381,N_10445);
nand U10529 (N_10529,N_10363,N_10407);
and U10530 (N_10530,N_10234,N_10284);
xnor U10531 (N_10531,N_10409,N_10245);
or U10532 (N_10532,N_10400,N_10243);
xnor U10533 (N_10533,N_10413,N_10237);
or U10534 (N_10534,N_10246,N_10379);
nor U10535 (N_10535,N_10216,N_10415);
xnor U10536 (N_10536,N_10228,N_10359);
nand U10537 (N_10537,N_10305,N_10214);
xnor U10538 (N_10538,N_10329,N_10269);
or U10539 (N_10539,N_10423,N_10447);
nor U10540 (N_10540,N_10239,N_10318);
nand U10541 (N_10541,N_10395,N_10332);
and U10542 (N_10542,N_10365,N_10341);
nand U10543 (N_10543,N_10349,N_10431);
nor U10544 (N_10544,N_10325,N_10364);
or U10545 (N_10545,N_10355,N_10462);
xnor U10546 (N_10546,N_10259,N_10390);
or U10547 (N_10547,N_10258,N_10319);
xnor U10548 (N_10548,N_10358,N_10205);
and U10549 (N_10549,N_10327,N_10429);
or U10550 (N_10550,N_10295,N_10202);
xnor U10551 (N_10551,N_10410,N_10476);
and U10552 (N_10552,N_10416,N_10334);
and U10553 (N_10553,N_10496,N_10201);
and U10554 (N_10554,N_10310,N_10302);
or U10555 (N_10555,N_10322,N_10283);
or U10556 (N_10556,N_10368,N_10315);
or U10557 (N_10557,N_10309,N_10491);
or U10558 (N_10558,N_10314,N_10389);
and U10559 (N_10559,N_10215,N_10495);
xor U10560 (N_10560,N_10219,N_10377);
nor U10561 (N_10561,N_10304,N_10427);
and U10562 (N_10562,N_10432,N_10478);
or U10563 (N_10563,N_10265,N_10339);
and U10564 (N_10564,N_10260,N_10367);
xnor U10565 (N_10565,N_10419,N_10278);
or U10566 (N_10566,N_10348,N_10200);
nor U10567 (N_10567,N_10472,N_10208);
nor U10568 (N_10568,N_10440,N_10204);
nor U10569 (N_10569,N_10221,N_10420);
xor U10570 (N_10570,N_10437,N_10424);
nand U10571 (N_10571,N_10446,N_10264);
xor U10572 (N_10572,N_10499,N_10317);
nand U10573 (N_10573,N_10231,N_10337);
or U10574 (N_10574,N_10371,N_10210);
or U10575 (N_10575,N_10441,N_10418);
nor U10576 (N_10576,N_10378,N_10230);
nand U10577 (N_10577,N_10320,N_10207);
nand U10578 (N_10578,N_10477,N_10203);
and U10579 (N_10579,N_10292,N_10298);
and U10580 (N_10580,N_10481,N_10455);
and U10581 (N_10581,N_10217,N_10357);
xnor U10582 (N_10582,N_10405,N_10335);
nor U10583 (N_10583,N_10483,N_10301);
and U10584 (N_10584,N_10209,N_10374);
nand U10585 (N_10585,N_10262,N_10474);
nor U10586 (N_10586,N_10489,N_10312);
and U10587 (N_10587,N_10360,N_10324);
xor U10588 (N_10588,N_10475,N_10376);
nand U10589 (N_10589,N_10452,N_10280);
and U10590 (N_10590,N_10282,N_10307);
or U10591 (N_10591,N_10285,N_10351);
and U10592 (N_10592,N_10287,N_10497);
xor U10593 (N_10593,N_10492,N_10362);
and U10594 (N_10594,N_10387,N_10456);
xnor U10595 (N_10595,N_10464,N_10336);
and U10596 (N_10596,N_10296,N_10463);
and U10597 (N_10597,N_10242,N_10257);
nor U10598 (N_10598,N_10369,N_10421);
and U10599 (N_10599,N_10469,N_10225);
nor U10600 (N_10600,N_10227,N_10430);
or U10601 (N_10601,N_10466,N_10453);
xnor U10602 (N_10602,N_10385,N_10286);
nor U10603 (N_10603,N_10323,N_10352);
xnor U10604 (N_10604,N_10490,N_10233);
nand U10605 (N_10605,N_10300,N_10450);
and U10606 (N_10606,N_10249,N_10338);
nand U10607 (N_10607,N_10206,N_10484);
nor U10608 (N_10608,N_10345,N_10397);
nor U10609 (N_10609,N_10479,N_10311);
nor U10610 (N_10610,N_10238,N_10370);
or U10611 (N_10611,N_10375,N_10380);
or U10612 (N_10612,N_10470,N_10218);
nand U10613 (N_10613,N_10461,N_10414);
nor U10614 (N_10614,N_10288,N_10487);
or U10615 (N_10615,N_10486,N_10467);
nand U10616 (N_10616,N_10428,N_10290);
and U10617 (N_10617,N_10451,N_10401);
nand U10618 (N_10618,N_10293,N_10443);
and U10619 (N_10619,N_10454,N_10333);
or U10620 (N_10620,N_10211,N_10436);
and U10621 (N_10621,N_10250,N_10361);
nand U10622 (N_10622,N_10384,N_10340);
and U10623 (N_10623,N_10326,N_10403);
xor U10624 (N_10624,N_10313,N_10356);
nor U10625 (N_10625,N_10425,N_10291);
and U10626 (N_10626,N_10346,N_10406);
or U10627 (N_10627,N_10276,N_10460);
xor U10628 (N_10628,N_10383,N_10261);
xor U10629 (N_10629,N_10297,N_10404);
nand U10630 (N_10630,N_10270,N_10251);
and U10631 (N_10631,N_10433,N_10480);
or U10632 (N_10632,N_10279,N_10388);
nand U10633 (N_10633,N_10266,N_10223);
and U10634 (N_10634,N_10493,N_10247);
xor U10635 (N_10635,N_10402,N_10224);
and U10636 (N_10636,N_10220,N_10303);
xnor U10637 (N_10637,N_10316,N_10308);
or U10638 (N_10638,N_10330,N_10494);
or U10639 (N_10639,N_10382,N_10448);
or U10640 (N_10640,N_10306,N_10347);
and U10641 (N_10641,N_10226,N_10235);
nor U10642 (N_10642,N_10398,N_10408);
or U10643 (N_10643,N_10386,N_10212);
nor U10644 (N_10644,N_10229,N_10342);
and U10645 (N_10645,N_10366,N_10393);
and U10646 (N_10646,N_10411,N_10422);
and U10647 (N_10647,N_10240,N_10444);
nor U10648 (N_10648,N_10263,N_10391);
and U10649 (N_10649,N_10426,N_10449);
or U10650 (N_10650,N_10314,N_10286);
nand U10651 (N_10651,N_10278,N_10294);
nand U10652 (N_10652,N_10499,N_10266);
and U10653 (N_10653,N_10338,N_10346);
xor U10654 (N_10654,N_10213,N_10312);
nor U10655 (N_10655,N_10254,N_10242);
and U10656 (N_10656,N_10406,N_10480);
and U10657 (N_10657,N_10471,N_10279);
and U10658 (N_10658,N_10498,N_10409);
and U10659 (N_10659,N_10345,N_10440);
nor U10660 (N_10660,N_10487,N_10375);
nor U10661 (N_10661,N_10395,N_10404);
nor U10662 (N_10662,N_10406,N_10493);
xor U10663 (N_10663,N_10384,N_10325);
and U10664 (N_10664,N_10483,N_10201);
or U10665 (N_10665,N_10212,N_10316);
or U10666 (N_10666,N_10387,N_10321);
and U10667 (N_10667,N_10243,N_10436);
or U10668 (N_10668,N_10489,N_10402);
xnor U10669 (N_10669,N_10367,N_10207);
xnor U10670 (N_10670,N_10372,N_10358);
or U10671 (N_10671,N_10376,N_10270);
nand U10672 (N_10672,N_10254,N_10405);
or U10673 (N_10673,N_10201,N_10249);
and U10674 (N_10674,N_10226,N_10416);
and U10675 (N_10675,N_10284,N_10344);
xor U10676 (N_10676,N_10410,N_10467);
nor U10677 (N_10677,N_10265,N_10345);
or U10678 (N_10678,N_10358,N_10430);
nand U10679 (N_10679,N_10374,N_10221);
nand U10680 (N_10680,N_10411,N_10384);
nor U10681 (N_10681,N_10293,N_10244);
nand U10682 (N_10682,N_10421,N_10420);
nor U10683 (N_10683,N_10257,N_10235);
nand U10684 (N_10684,N_10340,N_10488);
nor U10685 (N_10685,N_10314,N_10461);
xnor U10686 (N_10686,N_10468,N_10221);
nor U10687 (N_10687,N_10454,N_10320);
nand U10688 (N_10688,N_10487,N_10484);
nor U10689 (N_10689,N_10465,N_10293);
and U10690 (N_10690,N_10370,N_10494);
nor U10691 (N_10691,N_10228,N_10406);
nor U10692 (N_10692,N_10247,N_10409);
xnor U10693 (N_10693,N_10333,N_10221);
or U10694 (N_10694,N_10333,N_10386);
nand U10695 (N_10695,N_10402,N_10266);
nand U10696 (N_10696,N_10357,N_10401);
xor U10697 (N_10697,N_10317,N_10468);
and U10698 (N_10698,N_10300,N_10282);
xor U10699 (N_10699,N_10434,N_10401);
nor U10700 (N_10700,N_10336,N_10380);
nand U10701 (N_10701,N_10457,N_10455);
nor U10702 (N_10702,N_10492,N_10271);
xor U10703 (N_10703,N_10491,N_10408);
and U10704 (N_10704,N_10399,N_10395);
nor U10705 (N_10705,N_10421,N_10375);
xor U10706 (N_10706,N_10220,N_10209);
and U10707 (N_10707,N_10346,N_10461);
and U10708 (N_10708,N_10203,N_10483);
or U10709 (N_10709,N_10204,N_10304);
nor U10710 (N_10710,N_10296,N_10362);
or U10711 (N_10711,N_10267,N_10371);
and U10712 (N_10712,N_10263,N_10407);
and U10713 (N_10713,N_10429,N_10271);
nand U10714 (N_10714,N_10449,N_10287);
or U10715 (N_10715,N_10352,N_10331);
nand U10716 (N_10716,N_10346,N_10289);
nor U10717 (N_10717,N_10300,N_10215);
xor U10718 (N_10718,N_10358,N_10280);
nand U10719 (N_10719,N_10365,N_10292);
xor U10720 (N_10720,N_10274,N_10458);
or U10721 (N_10721,N_10395,N_10440);
or U10722 (N_10722,N_10333,N_10335);
nand U10723 (N_10723,N_10374,N_10383);
xor U10724 (N_10724,N_10373,N_10204);
nand U10725 (N_10725,N_10234,N_10255);
xor U10726 (N_10726,N_10227,N_10426);
nor U10727 (N_10727,N_10304,N_10271);
nand U10728 (N_10728,N_10225,N_10353);
or U10729 (N_10729,N_10382,N_10377);
or U10730 (N_10730,N_10419,N_10407);
xnor U10731 (N_10731,N_10349,N_10252);
nand U10732 (N_10732,N_10434,N_10358);
or U10733 (N_10733,N_10296,N_10378);
nand U10734 (N_10734,N_10210,N_10299);
or U10735 (N_10735,N_10370,N_10392);
nor U10736 (N_10736,N_10347,N_10205);
xor U10737 (N_10737,N_10248,N_10381);
or U10738 (N_10738,N_10375,N_10258);
and U10739 (N_10739,N_10335,N_10475);
or U10740 (N_10740,N_10351,N_10241);
or U10741 (N_10741,N_10392,N_10462);
or U10742 (N_10742,N_10361,N_10329);
nand U10743 (N_10743,N_10269,N_10282);
xor U10744 (N_10744,N_10406,N_10462);
nand U10745 (N_10745,N_10268,N_10302);
and U10746 (N_10746,N_10350,N_10232);
xor U10747 (N_10747,N_10482,N_10430);
xor U10748 (N_10748,N_10377,N_10404);
and U10749 (N_10749,N_10252,N_10207);
or U10750 (N_10750,N_10306,N_10402);
xnor U10751 (N_10751,N_10448,N_10342);
nand U10752 (N_10752,N_10417,N_10389);
nor U10753 (N_10753,N_10355,N_10203);
nand U10754 (N_10754,N_10204,N_10365);
nor U10755 (N_10755,N_10260,N_10381);
and U10756 (N_10756,N_10239,N_10376);
nand U10757 (N_10757,N_10495,N_10372);
nor U10758 (N_10758,N_10381,N_10206);
and U10759 (N_10759,N_10360,N_10418);
nor U10760 (N_10760,N_10465,N_10388);
nor U10761 (N_10761,N_10331,N_10367);
nand U10762 (N_10762,N_10242,N_10488);
xor U10763 (N_10763,N_10451,N_10293);
nand U10764 (N_10764,N_10216,N_10277);
and U10765 (N_10765,N_10250,N_10330);
or U10766 (N_10766,N_10433,N_10321);
and U10767 (N_10767,N_10392,N_10460);
or U10768 (N_10768,N_10244,N_10308);
and U10769 (N_10769,N_10239,N_10275);
xor U10770 (N_10770,N_10281,N_10217);
nand U10771 (N_10771,N_10417,N_10292);
nor U10772 (N_10772,N_10290,N_10362);
and U10773 (N_10773,N_10476,N_10216);
nor U10774 (N_10774,N_10229,N_10259);
or U10775 (N_10775,N_10367,N_10483);
xor U10776 (N_10776,N_10276,N_10304);
nand U10777 (N_10777,N_10373,N_10428);
nand U10778 (N_10778,N_10293,N_10310);
nand U10779 (N_10779,N_10319,N_10221);
nor U10780 (N_10780,N_10274,N_10402);
or U10781 (N_10781,N_10416,N_10289);
xnor U10782 (N_10782,N_10387,N_10486);
and U10783 (N_10783,N_10400,N_10386);
xnor U10784 (N_10784,N_10254,N_10322);
nand U10785 (N_10785,N_10495,N_10477);
nand U10786 (N_10786,N_10457,N_10303);
or U10787 (N_10787,N_10479,N_10271);
nand U10788 (N_10788,N_10267,N_10486);
xnor U10789 (N_10789,N_10436,N_10233);
nand U10790 (N_10790,N_10206,N_10412);
nand U10791 (N_10791,N_10343,N_10340);
nand U10792 (N_10792,N_10373,N_10200);
and U10793 (N_10793,N_10329,N_10219);
xnor U10794 (N_10794,N_10404,N_10476);
nor U10795 (N_10795,N_10225,N_10403);
nand U10796 (N_10796,N_10330,N_10235);
nand U10797 (N_10797,N_10453,N_10290);
or U10798 (N_10798,N_10483,N_10310);
nor U10799 (N_10799,N_10259,N_10399);
and U10800 (N_10800,N_10668,N_10525);
nand U10801 (N_10801,N_10763,N_10604);
nand U10802 (N_10802,N_10594,N_10683);
and U10803 (N_10803,N_10646,N_10635);
and U10804 (N_10804,N_10709,N_10545);
or U10805 (N_10805,N_10643,N_10723);
nand U10806 (N_10806,N_10760,N_10516);
and U10807 (N_10807,N_10622,N_10618);
and U10808 (N_10808,N_10770,N_10510);
and U10809 (N_10809,N_10722,N_10680);
nand U10810 (N_10810,N_10521,N_10685);
xnor U10811 (N_10811,N_10675,N_10582);
nor U10812 (N_10812,N_10662,N_10543);
nand U10813 (N_10813,N_10515,N_10684);
or U10814 (N_10814,N_10529,N_10676);
and U10815 (N_10815,N_10728,N_10737);
xor U10816 (N_10816,N_10561,N_10562);
and U10817 (N_10817,N_10745,N_10798);
xor U10818 (N_10818,N_10551,N_10747);
xnor U10819 (N_10819,N_10508,N_10780);
and U10820 (N_10820,N_10678,N_10611);
nor U10821 (N_10821,N_10571,N_10575);
nor U10822 (N_10822,N_10522,N_10593);
and U10823 (N_10823,N_10524,N_10795);
xor U10824 (N_10824,N_10659,N_10653);
xnor U10825 (N_10825,N_10616,N_10679);
nor U10826 (N_10826,N_10632,N_10609);
and U10827 (N_10827,N_10619,N_10540);
nor U10828 (N_10828,N_10563,N_10781);
and U10829 (N_10829,N_10667,N_10577);
and U10830 (N_10830,N_10520,N_10782);
nor U10831 (N_10831,N_10740,N_10692);
or U10832 (N_10832,N_10603,N_10509);
nand U10833 (N_10833,N_10537,N_10691);
nor U10834 (N_10834,N_10787,N_10598);
or U10835 (N_10835,N_10584,N_10559);
nand U10836 (N_10836,N_10757,N_10707);
nor U10837 (N_10837,N_10642,N_10704);
nor U10838 (N_10838,N_10710,N_10518);
nand U10839 (N_10839,N_10553,N_10601);
and U10840 (N_10840,N_10505,N_10673);
or U10841 (N_10841,N_10706,N_10533);
xnor U10842 (N_10842,N_10771,N_10719);
nor U10843 (N_10843,N_10556,N_10519);
nand U10844 (N_10844,N_10753,N_10777);
nor U10845 (N_10845,N_10565,N_10587);
and U10846 (N_10846,N_10568,N_10758);
and U10847 (N_10847,N_10630,N_10769);
nor U10848 (N_10848,N_10738,N_10644);
xor U10849 (N_10849,N_10681,N_10569);
or U10850 (N_10850,N_10656,N_10796);
xnor U10851 (N_10851,N_10712,N_10666);
xnor U10852 (N_10852,N_10754,N_10655);
nor U10853 (N_10853,N_10726,N_10661);
or U10854 (N_10854,N_10602,N_10547);
and U10855 (N_10855,N_10744,N_10645);
nor U10856 (N_10856,N_10688,N_10640);
and U10857 (N_10857,N_10576,N_10589);
nand U10858 (N_10858,N_10654,N_10535);
and U10859 (N_10859,N_10658,N_10773);
nand U10860 (N_10860,N_10652,N_10698);
xnor U10861 (N_10861,N_10513,N_10793);
nor U10862 (N_10862,N_10566,N_10720);
xor U10863 (N_10863,N_10702,N_10665);
nor U10864 (N_10864,N_10752,N_10613);
and U10865 (N_10865,N_10549,N_10765);
nor U10866 (N_10866,N_10605,N_10558);
nor U10867 (N_10867,N_10610,N_10620);
or U10868 (N_10868,N_10623,N_10625);
or U10869 (N_10869,N_10785,N_10799);
or U10870 (N_10870,N_10790,N_10621);
and U10871 (N_10871,N_10748,N_10682);
nor U10872 (N_10872,N_10732,N_10607);
nand U10873 (N_10873,N_10523,N_10669);
or U10874 (N_10874,N_10541,N_10786);
nor U10875 (N_10875,N_10555,N_10542);
xor U10876 (N_10876,N_10671,N_10767);
or U10877 (N_10877,N_10651,N_10731);
nand U10878 (N_10878,N_10701,N_10727);
nand U10879 (N_10879,N_10742,N_10538);
and U10880 (N_10880,N_10664,N_10776);
xnor U10881 (N_10881,N_10660,N_10534);
xor U10882 (N_10882,N_10511,N_10628);
nand U10883 (N_10883,N_10591,N_10638);
or U10884 (N_10884,N_10670,N_10705);
nor U10885 (N_10885,N_10637,N_10531);
nand U10886 (N_10886,N_10590,N_10581);
and U10887 (N_10887,N_10749,N_10716);
nor U10888 (N_10888,N_10764,N_10755);
nand U10889 (N_10889,N_10506,N_10703);
xor U10890 (N_10890,N_10759,N_10750);
nor U10891 (N_10891,N_10708,N_10648);
nor U10892 (N_10892,N_10746,N_10714);
and U10893 (N_10893,N_10774,N_10768);
xnor U10894 (N_10894,N_10629,N_10624);
xnor U10895 (N_10895,N_10532,N_10500);
and U10896 (N_10896,N_10792,N_10606);
or U10897 (N_10897,N_10564,N_10557);
or U10898 (N_10898,N_10588,N_10784);
or U10899 (N_10899,N_10762,N_10528);
or U10900 (N_10900,N_10689,N_10633);
and U10901 (N_10901,N_10583,N_10677);
or U10902 (N_10902,N_10711,N_10779);
nand U10903 (N_10903,N_10687,N_10626);
nand U10904 (N_10904,N_10733,N_10717);
and U10905 (N_10905,N_10695,N_10578);
nor U10906 (N_10906,N_10579,N_10503);
nand U10907 (N_10907,N_10736,N_10592);
xor U10908 (N_10908,N_10586,N_10512);
nor U10909 (N_10909,N_10696,N_10686);
and U10910 (N_10910,N_10693,N_10791);
or U10911 (N_10911,N_10788,N_10674);
nor U10912 (N_10912,N_10504,N_10572);
nor U10913 (N_10913,N_10649,N_10734);
nor U10914 (N_10914,N_10690,N_10548);
nand U10915 (N_10915,N_10721,N_10550);
nor U10916 (N_10916,N_10599,N_10725);
xor U10917 (N_10917,N_10650,N_10775);
xor U10918 (N_10918,N_10614,N_10766);
xnor U10919 (N_10919,N_10608,N_10789);
xor U10920 (N_10920,N_10597,N_10718);
and U10921 (N_10921,N_10517,N_10552);
nor U10922 (N_10922,N_10697,N_10539);
nand U10923 (N_10923,N_10596,N_10699);
and U10924 (N_10924,N_10570,N_10729);
and U10925 (N_10925,N_10595,N_10600);
xnor U10926 (N_10926,N_10730,N_10527);
nand U10927 (N_10927,N_10617,N_10772);
nor U10928 (N_10928,N_10634,N_10739);
xor U10929 (N_10929,N_10526,N_10530);
and U10930 (N_10930,N_10636,N_10514);
xnor U10931 (N_10931,N_10778,N_10544);
and U10932 (N_10932,N_10797,N_10713);
nand U10933 (N_10933,N_10672,N_10724);
and U10934 (N_10934,N_10700,N_10756);
nor U10935 (N_10935,N_10647,N_10546);
xnor U10936 (N_10936,N_10761,N_10641);
nor U10937 (N_10937,N_10536,N_10735);
or U10938 (N_10938,N_10580,N_10567);
and U10939 (N_10939,N_10615,N_10783);
or U10940 (N_10940,N_10794,N_10573);
xnor U10941 (N_10941,N_10627,N_10631);
or U10942 (N_10942,N_10657,N_10507);
xor U10943 (N_10943,N_10560,N_10501);
and U10944 (N_10944,N_10715,N_10554);
xnor U10945 (N_10945,N_10743,N_10502);
xnor U10946 (N_10946,N_10694,N_10741);
or U10947 (N_10947,N_10663,N_10574);
nand U10948 (N_10948,N_10751,N_10612);
or U10949 (N_10949,N_10639,N_10585);
xnor U10950 (N_10950,N_10571,N_10762);
or U10951 (N_10951,N_10595,N_10695);
nor U10952 (N_10952,N_10773,N_10669);
and U10953 (N_10953,N_10767,N_10525);
and U10954 (N_10954,N_10768,N_10578);
xnor U10955 (N_10955,N_10748,N_10517);
or U10956 (N_10956,N_10747,N_10510);
and U10957 (N_10957,N_10566,N_10741);
nor U10958 (N_10958,N_10754,N_10639);
xnor U10959 (N_10959,N_10522,N_10516);
nand U10960 (N_10960,N_10738,N_10521);
nor U10961 (N_10961,N_10529,N_10715);
xor U10962 (N_10962,N_10631,N_10738);
and U10963 (N_10963,N_10650,N_10777);
nor U10964 (N_10964,N_10659,N_10687);
and U10965 (N_10965,N_10535,N_10780);
nand U10966 (N_10966,N_10615,N_10530);
xnor U10967 (N_10967,N_10584,N_10742);
and U10968 (N_10968,N_10523,N_10688);
nand U10969 (N_10969,N_10752,N_10611);
nand U10970 (N_10970,N_10774,N_10682);
and U10971 (N_10971,N_10654,N_10522);
or U10972 (N_10972,N_10734,N_10629);
nand U10973 (N_10973,N_10678,N_10658);
xnor U10974 (N_10974,N_10716,N_10579);
xnor U10975 (N_10975,N_10783,N_10719);
and U10976 (N_10976,N_10659,N_10729);
xnor U10977 (N_10977,N_10745,N_10693);
or U10978 (N_10978,N_10541,N_10603);
nor U10979 (N_10979,N_10601,N_10755);
or U10980 (N_10980,N_10602,N_10566);
or U10981 (N_10981,N_10554,N_10622);
nand U10982 (N_10982,N_10553,N_10515);
and U10983 (N_10983,N_10684,N_10557);
and U10984 (N_10984,N_10592,N_10727);
xor U10985 (N_10985,N_10666,N_10575);
or U10986 (N_10986,N_10621,N_10729);
and U10987 (N_10987,N_10559,N_10798);
xnor U10988 (N_10988,N_10507,N_10662);
nor U10989 (N_10989,N_10549,N_10733);
or U10990 (N_10990,N_10730,N_10608);
and U10991 (N_10991,N_10741,N_10592);
and U10992 (N_10992,N_10740,N_10729);
nand U10993 (N_10993,N_10659,N_10675);
nand U10994 (N_10994,N_10633,N_10535);
nor U10995 (N_10995,N_10594,N_10634);
nor U10996 (N_10996,N_10609,N_10784);
or U10997 (N_10997,N_10719,N_10787);
or U10998 (N_10998,N_10651,N_10557);
nor U10999 (N_10999,N_10605,N_10623);
xnor U11000 (N_11000,N_10707,N_10606);
and U11001 (N_11001,N_10730,N_10722);
nand U11002 (N_11002,N_10731,N_10539);
xor U11003 (N_11003,N_10694,N_10660);
nor U11004 (N_11004,N_10605,N_10765);
xnor U11005 (N_11005,N_10665,N_10552);
and U11006 (N_11006,N_10713,N_10664);
nor U11007 (N_11007,N_10624,N_10610);
nand U11008 (N_11008,N_10630,N_10643);
xor U11009 (N_11009,N_10632,N_10506);
nor U11010 (N_11010,N_10560,N_10791);
xor U11011 (N_11011,N_10593,N_10617);
nand U11012 (N_11012,N_10662,N_10671);
nand U11013 (N_11013,N_10723,N_10677);
xor U11014 (N_11014,N_10602,N_10717);
xnor U11015 (N_11015,N_10724,N_10676);
or U11016 (N_11016,N_10569,N_10589);
xor U11017 (N_11017,N_10623,N_10757);
and U11018 (N_11018,N_10607,N_10581);
or U11019 (N_11019,N_10564,N_10530);
nor U11020 (N_11020,N_10592,N_10694);
or U11021 (N_11021,N_10595,N_10526);
nand U11022 (N_11022,N_10512,N_10603);
nor U11023 (N_11023,N_10678,N_10574);
nor U11024 (N_11024,N_10512,N_10744);
nand U11025 (N_11025,N_10730,N_10783);
and U11026 (N_11026,N_10510,N_10740);
or U11027 (N_11027,N_10764,N_10778);
xnor U11028 (N_11028,N_10746,N_10768);
nor U11029 (N_11029,N_10733,N_10714);
and U11030 (N_11030,N_10500,N_10787);
or U11031 (N_11031,N_10603,N_10722);
nand U11032 (N_11032,N_10563,N_10678);
nor U11033 (N_11033,N_10641,N_10661);
or U11034 (N_11034,N_10679,N_10595);
and U11035 (N_11035,N_10619,N_10526);
nor U11036 (N_11036,N_10718,N_10642);
and U11037 (N_11037,N_10728,N_10782);
or U11038 (N_11038,N_10676,N_10581);
xnor U11039 (N_11039,N_10651,N_10500);
nor U11040 (N_11040,N_10556,N_10761);
xor U11041 (N_11041,N_10536,N_10751);
xnor U11042 (N_11042,N_10578,N_10663);
nor U11043 (N_11043,N_10690,N_10711);
xnor U11044 (N_11044,N_10572,N_10577);
nor U11045 (N_11045,N_10781,N_10585);
or U11046 (N_11046,N_10501,N_10727);
or U11047 (N_11047,N_10701,N_10616);
or U11048 (N_11048,N_10783,N_10614);
nand U11049 (N_11049,N_10775,N_10730);
xor U11050 (N_11050,N_10618,N_10769);
and U11051 (N_11051,N_10798,N_10561);
nand U11052 (N_11052,N_10561,N_10613);
nand U11053 (N_11053,N_10740,N_10769);
nand U11054 (N_11054,N_10658,N_10755);
nand U11055 (N_11055,N_10619,N_10545);
xnor U11056 (N_11056,N_10507,N_10771);
or U11057 (N_11057,N_10724,N_10634);
xnor U11058 (N_11058,N_10798,N_10572);
nor U11059 (N_11059,N_10531,N_10668);
xor U11060 (N_11060,N_10617,N_10693);
nand U11061 (N_11061,N_10640,N_10676);
nand U11062 (N_11062,N_10774,N_10750);
nor U11063 (N_11063,N_10760,N_10762);
nand U11064 (N_11064,N_10583,N_10590);
or U11065 (N_11065,N_10584,N_10528);
nor U11066 (N_11066,N_10540,N_10678);
or U11067 (N_11067,N_10648,N_10549);
or U11068 (N_11068,N_10509,N_10571);
nor U11069 (N_11069,N_10608,N_10580);
nor U11070 (N_11070,N_10759,N_10621);
nand U11071 (N_11071,N_10501,N_10509);
nand U11072 (N_11072,N_10652,N_10629);
nor U11073 (N_11073,N_10558,N_10713);
nor U11074 (N_11074,N_10610,N_10637);
or U11075 (N_11075,N_10583,N_10627);
xor U11076 (N_11076,N_10712,N_10751);
xor U11077 (N_11077,N_10538,N_10610);
nand U11078 (N_11078,N_10548,N_10568);
nor U11079 (N_11079,N_10688,N_10612);
nor U11080 (N_11080,N_10610,N_10550);
nor U11081 (N_11081,N_10541,N_10581);
and U11082 (N_11082,N_10759,N_10611);
xor U11083 (N_11083,N_10652,N_10760);
xnor U11084 (N_11084,N_10732,N_10637);
nand U11085 (N_11085,N_10685,N_10635);
nand U11086 (N_11086,N_10779,N_10699);
or U11087 (N_11087,N_10542,N_10575);
nand U11088 (N_11088,N_10794,N_10798);
or U11089 (N_11089,N_10784,N_10726);
nand U11090 (N_11090,N_10538,N_10519);
and U11091 (N_11091,N_10679,N_10699);
nand U11092 (N_11092,N_10793,N_10709);
or U11093 (N_11093,N_10665,N_10717);
or U11094 (N_11094,N_10748,N_10663);
or U11095 (N_11095,N_10634,N_10735);
xnor U11096 (N_11096,N_10676,N_10685);
or U11097 (N_11097,N_10530,N_10563);
and U11098 (N_11098,N_10796,N_10662);
nor U11099 (N_11099,N_10787,N_10771);
or U11100 (N_11100,N_11038,N_10824);
and U11101 (N_11101,N_10979,N_10896);
or U11102 (N_11102,N_10935,N_10906);
or U11103 (N_11103,N_11055,N_10870);
nand U11104 (N_11104,N_10818,N_10868);
xor U11105 (N_11105,N_11019,N_11075);
xnor U11106 (N_11106,N_11007,N_11014);
or U11107 (N_11107,N_11042,N_11064);
and U11108 (N_11108,N_11067,N_11023);
nor U11109 (N_11109,N_10848,N_11018);
nand U11110 (N_11110,N_10968,N_11054);
and U11111 (N_11111,N_10965,N_11086);
nand U11112 (N_11112,N_10852,N_10922);
xor U11113 (N_11113,N_10980,N_11028);
xnor U11114 (N_11114,N_10994,N_10806);
nand U11115 (N_11115,N_10856,N_11081);
xor U11116 (N_11116,N_10850,N_10819);
and U11117 (N_11117,N_11000,N_10891);
xnor U11118 (N_11118,N_11003,N_11099);
nand U11119 (N_11119,N_11010,N_10944);
or U11120 (N_11120,N_11070,N_10826);
or U11121 (N_11121,N_10854,N_10992);
xor U11122 (N_11122,N_10801,N_10936);
nor U11123 (N_11123,N_10961,N_10841);
nand U11124 (N_11124,N_11068,N_10836);
and U11125 (N_11125,N_10957,N_11059);
xnor U11126 (N_11126,N_10902,N_11091);
and U11127 (N_11127,N_10978,N_10910);
or U11128 (N_11128,N_10873,N_10828);
or U11129 (N_11129,N_11058,N_10898);
nor U11130 (N_11130,N_10872,N_10915);
or U11131 (N_11131,N_10901,N_11006);
or U11132 (N_11132,N_10827,N_10977);
nand U11133 (N_11133,N_11036,N_10830);
nand U11134 (N_11134,N_10812,N_11088);
nor U11135 (N_11135,N_10934,N_11008);
nand U11136 (N_11136,N_11078,N_10807);
xnor U11137 (N_11137,N_11049,N_11044);
or U11138 (N_11138,N_10859,N_10986);
nand U11139 (N_11139,N_10863,N_10843);
nor U11140 (N_11140,N_10838,N_10820);
nor U11141 (N_11141,N_10948,N_11097);
xor U11142 (N_11142,N_10970,N_10943);
and U11143 (N_11143,N_10991,N_10800);
nor U11144 (N_11144,N_10908,N_11009);
or U11145 (N_11145,N_10881,N_10969);
nand U11146 (N_11146,N_10962,N_11056);
nand U11147 (N_11147,N_11062,N_11074);
and U11148 (N_11148,N_10884,N_10972);
or U11149 (N_11149,N_11022,N_10844);
xor U11150 (N_11150,N_11061,N_10993);
nor U11151 (N_11151,N_10967,N_10833);
xnor U11152 (N_11152,N_10938,N_11098);
nand U11153 (N_11153,N_10846,N_11015);
nand U11154 (N_11154,N_10897,N_10959);
nand U11155 (N_11155,N_11095,N_11071);
nand U11156 (N_11156,N_11005,N_10858);
nand U11157 (N_11157,N_10855,N_10914);
nand U11158 (N_11158,N_10808,N_11065);
xnor U11159 (N_11159,N_10995,N_11030);
or U11160 (N_11160,N_11013,N_10887);
and U11161 (N_11161,N_11024,N_11096);
xnor U11162 (N_11162,N_10921,N_10939);
nand U11163 (N_11163,N_11020,N_11077);
and U11164 (N_11164,N_10817,N_10883);
xor U11165 (N_11165,N_10917,N_10985);
or U11166 (N_11166,N_10952,N_11052);
nand U11167 (N_11167,N_10950,N_10842);
or U11168 (N_11168,N_10880,N_11035);
xnor U11169 (N_11169,N_10871,N_11087);
nor U11170 (N_11170,N_10916,N_11080);
nor U11171 (N_11171,N_11089,N_11051);
xnor U11172 (N_11172,N_10821,N_10953);
xor U11173 (N_11173,N_11079,N_11083);
nor U11174 (N_11174,N_10971,N_10892);
nand U11175 (N_11175,N_10853,N_10927);
nand U11176 (N_11176,N_10814,N_10882);
nand U11177 (N_11177,N_10813,N_11039);
nand U11178 (N_11178,N_11053,N_10857);
and U11179 (N_11179,N_10829,N_10894);
or U11180 (N_11180,N_10890,N_10928);
and U11181 (N_11181,N_11031,N_10816);
xor U11182 (N_11182,N_11040,N_10989);
or U11183 (N_11183,N_11085,N_10941);
xor U11184 (N_11184,N_11043,N_10864);
nor U11185 (N_11185,N_11076,N_10840);
nand U11186 (N_11186,N_11029,N_10832);
or U11187 (N_11187,N_10929,N_10924);
and U11188 (N_11188,N_10988,N_10946);
nand U11189 (N_11189,N_11084,N_11001);
or U11190 (N_11190,N_10925,N_10804);
and U11191 (N_11191,N_10974,N_10923);
nand U11192 (N_11192,N_10876,N_10920);
and U11193 (N_11193,N_11002,N_10885);
or U11194 (N_11194,N_11026,N_10956);
nand U11195 (N_11195,N_11063,N_10899);
nand U11196 (N_11196,N_10918,N_10895);
nor U11197 (N_11197,N_10987,N_11004);
and U11198 (N_11198,N_10937,N_11066);
nand U11199 (N_11199,N_11073,N_10886);
nor U11200 (N_11200,N_10849,N_10942);
xnor U11201 (N_11201,N_10867,N_10866);
nor U11202 (N_11202,N_10878,N_10805);
xor U11203 (N_11203,N_10837,N_10976);
and U11204 (N_11204,N_11045,N_11069);
and U11205 (N_11205,N_10905,N_10879);
nand U11206 (N_11206,N_11057,N_10975);
nor U11207 (N_11207,N_11092,N_10984);
and U11208 (N_11208,N_10964,N_10932);
nand U11209 (N_11209,N_11032,N_11047);
nand U11210 (N_11210,N_11021,N_11025);
nand U11211 (N_11211,N_10823,N_10982);
nand U11212 (N_11212,N_10825,N_10990);
nor U11213 (N_11213,N_10909,N_10945);
nor U11214 (N_11214,N_10874,N_11046);
and U11215 (N_11215,N_10913,N_10877);
or U11216 (N_11216,N_10926,N_10809);
nor U11217 (N_11217,N_10822,N_10940);
nor U11218 (N_11218,N_10889,N_11094);
xor U11219 (N_11219,N_11093,N_10810);
nor U11220 (N_11220,N_10834,N_11050);
and U11221 (N_11221,N_11060,N_11041);
or U11222 (N_11222,N_10860,N_10861);
or U11223 (N_11223,N_10947,N_11090);
and U11224 (N_11224,N_10900,N_11016);
or U11225 (N_11225,N_10997,N_10893);
nand U11226 (N_11226,N_10862,N_11082);
and U11227 (N_11227,N_11034,N_10903);
or U11228 (N_11228,N_10803,N_10931);
and U11229 (N_11229,N_10869,N_10839);
or U11230 (N_11230,N_11011,N_10981);
and U11231 (N_11231,N_11037,N_10963);
and U11232 (N_11232,N_10847,N_11072);
or U11233 (N_11233,N_10949,N_10888);
xnor U11234 (N_11234,N_11033,N_11017);
xnor U11235 (N_11235,N_10904,N_10815);
nor U11236 (N_11236,N_10875,N_11012);
xor U11237 (N_11237,N_10831,N_10933);
xnor U11238 (N_11238,N_10951,N_10851);
xor U11239 (N_11239,N_10996,N_10983);
xor U11240 (N_11240,N_10998,N_10912);
nor U11241 (N_11241,N_10865,N_10973);
nand U11242 (N_11242,N_10930,N_10960);
nand U11243 (N_11243,N_10845,N_10911);
nor U11244 (N_11244,N_10966,N_10955);
nor U11245 (N_11245,N_10907,N_10954);
xnor U11246 (N_11246,N_10802,N_11027);
or U11247 (N_11247,N_10811,N_10958);
nor U11248 (N_11248,N_10999,N_10835);
nand U11249 (N_11249,N_10919,N_11048);
xnor U11250 (N_11250,N_10927,N_10896);
and U11251 (N_11251,N_10993,N_11041);
or U11252 (N_11252,N_10886,N_10815);
xor U11253 (N_11253,N_10972,N_10870);
xnor U11254 (N_11254,N_11074,N_10807);
nor U11255 (N_11255,N_10810,N_10963);
nand U11256 (N_11256,N_11092,N_11022);
or U11257 (N_11257,N_11049,N_10813);
nor U11258 (N_11258,N_10893,N_11043);
or U11259 (N_11259,N_10877,N_10963);
or U11260 (N_11260,N_10953,N_11088);
nor U11261 (N_11261,N_11021,N_10827);
xor U11262 (N_11262,N_11082,N_10979);
nand U11263 (N_11263,N_11096,N_10873);
xor U11264 (N_11264,N_10810,N_10828);
or U11265 (N_11265,N_10951,N_10816);
nand U11266 (N_11266,N_11076,N_11090);
nor U11267 (N_11267,N_10919,N_10933);
xnor U11268 (N_11268,N_10950,N_10957);
xor U11269 (N_11269,N_10956,N_10996);
nand U11270 (N_11270,N_10886,N_10979);
or U11271 (N_11271,N_10929,N_11066);
nand U11272 (N_11272,N_10873,N_11043);
nand U11273 (N_11273,N_11007,N_11095);
or U11274 (N_11274,N_11057,N_10864);
nand U11275 (N_11275,N_10867,N_10908);
xor U11276 (N_11276,N_11047,N_11043);
and U11277 (N_11277,N_10964,N_10839);
nand U11278 (N_11278,N_10871,N_11085);
and U11279 (N_11279,N_10838,N_10912);
or U11280 (N_11280,N_10975,N_10912);
and U11281 (N_11281,N_10973,N_10990);
xor U11282 (N_11282,N_10862,N_10919);
or U11283 (N_11283,N_10833,N_10839);
xnor U11284 (N_11284,N_10967,N_10906);
xor U11285 (N_11285,N_10957,N_10993);
and U11286 (N_11286,N_10858,N_10823);
nor U11287 (N_11287,N_10949,N_10985);
xor U11288 (N_11288,N_10954,N_10983);
or U11289 (N_11289,N_10812,N_10942);
or U11290 (N_11290,N_11099,N_10907);
nand U11291 (N_11291,N_11026,N_10954);
and U11292 (N_11292,N_10910,N_10887);
nor U11293 (N_11293,N_10822,N_11054);
nand U11294 (N_11294,N_11089,N_11063);
xnor U11295 (N_11295,N_10809,N_10871);
nand U11296 (N_11296,N_10946,N_11092);
and U11297 (N_11297,N_10839,N_10981);
nor U11298 (N_11298,N_11082,N_10814);
nor U11299 (N_11299,N_10836,N_10970);
nor U11300 (N_11300,N_10923,N_10882);
xnor U11301 (N_11301,N_10900,N_10960);
xnor U11302 (N_11302,N_10877,N_11045);
nand U11303 (N_11303,N_10890,N_10932);
or U11304 (N_11304,N_11001,N_11060);
nor U11305 (N_11305,N_11013,N_10943);
or U11306 (N_11306,N_10801,N_10859);
or U11307 (N_11307,N_10880,N_10910);
and U11308 (N_11308,N_10940,N_10987);
nor U11309 (N_11309,N_10837,N_11048);
nand U11310 (N_11310,N_11009,N_10856);
and U11311 (N_11311,N_10892,N_11052);
or U11312 (N_11312,N_11067,N_11079);
nand U11313 (N_11313,N_11074,N_10844);
xor U11314 (N_11314,N_11055,N_10986);
and U11315 (N_11315,N_10961,N_10990);
nand U11316 (N_11316,N_10959,N_11068);
nor U11317 (N_11317,N_10821,N_10935);
or U11318 (N_11318,N_10957,N_11008);
nor U11319 (N_11319,N_11043,N_10889);
xnor U11320 (N_11320,N_11047,N_10800);
nor U11321 (N_11321,N_11098,N_10817);
and U11322 (N_11322,N_11031,N_11062);
nor U11323 (N_11323,N_10948,N_11082);
nand U11324 (N_11324,N_10802,N_10926);
xnor U11325 (N_11325,N_11030,N_10858);
or U11326 (N_11326,N_11073,N_11037);
xnor U11327 (N_11327,N_11054,N_10902);
and U11328 (N_11328,N_10828,N_10869);
xnor U11329 (N_11329,N_10833,N_11017);
xor U11330 (N_11330,N_11087,N_10982);
xor U11331 (N_11331,N_10804,N_10885);
nor U11332 (N_11332,N_10844,N_10910);
and U11333 (N_11333,N_11074,N_11069);
and U11334 (N_11334,N_11086,N_11051);
nand U11335 (N_11335,N_10873,N_10867);
or U11336 (N_11336,N_10823,N_10873);
nand U11337 (N_11337,N_10817,N_10844);
nand U11338 (N_11338,N_10880,N_10922);
nor U11339 (N_11339,N_11087,N_10858);
nor U11340 (N_11340,N_11030,N_11057);
or U11341 (N_11341,N_10984,N_10915);
nand U11342 (N_11342,N_10990,N_11049);
nand U11343 (N_11343,N_10934,N_11025);
xnor U11344 (N_11344,N_11089,N_10935);
nor U11345 (N_11345,N_10956,N_10905);
xor U11346 (N_11346,N_10832,N_10835);
xor U11347 (N_11347,N_10821,N_10964);
nand U11348 (N_11348,N_11025,N_10947);
or U11349 (N_11349,N_11009,N_11058);
and U11350 (N_11350,N_10946,N_11047);
and U11351 (N_11351,N_10899,N_10971);
and U11352 (N_11352,N_11064,N_10806);
and U11353 (N_11353,N_11023,N_10938);
or U11354 (N_11354,N_10848,N_10821);
and U11355 (N_11355,N_10909,N_11015);
or U11356 (N_11356,N_11040,N_10951);
nor U11357 (N_11357,N_11059,N_11070);
nor U11358 (N_11358,N_10851,N_10976);
and U11359 (N_11359,N_10807,N_11032);
or U11360 (N_11360,N_11094,N_11077);
nand U11361 (N_11361,N_10955,N_10833);
xnor U11362 (N_11362,N_10903,N_10836);
and U11363 (N_11363,N_11071,N_10807);
nand U11364 (N_11364,N_10868,N_11098);
xor U11365 (N_11365,N_11087,N_10884);
nor U11366 (N_11366,N_10846,N_10847);
nand U11367 (N_11367,N_11095,N_10884);
and U11368 (N_11368,N_10903,N_10929);
nor U11369 (N_11369,N_11036,N_10980);
nor U11370 (N_11370,N_11086,N_10984);
or U11371 (N_11371,N_10924,N_10855);
xnor U11372 (N_11372,N_10991,N_10969);
nor U11373 (N_11373,N_11048,N_10884);
nor U11374 (N_11374,N_11096,N_10818);
nand U11375 (N_11375,N_11014,N_11079);
nand U11376 (N_11376,N_10923,N_11059);
nand U11377 (N_11377,N_11037,N_10833);
nor U11378 (N_11378,N_11026,N_10865);
and U11379 (N_11379,N_10870,N_10853);
and U11380 (N_11380,N_10880,N_10931);
and U11381 (N_11381,N_10922,N_10947);
nand U11382 (N_11382,N_10836,N_10873);
nand U11383 (N_11383,N_10950,N_10919);
nand U11384 (N_11384,N_11041,N_11026);
and U11385 (N_11385,N_11045,N_11067);
or U11386 (N_11386,N_10803,N_11009);
xnor U11387 (N_11387,N_10908,N_10996);
xnor U11388 (N_11388,N_11044,N_10938);
nand U11389 (N_11389,N_10912,N_10970);
xnor U11390 (N_11390,N_10935,N_11017);
nand U11391 (N_11391,N_10951,N_10902);
nor U11392 (N_11392,N_11005,N_10931);
nand U11393 (N_11393,N_10997,N_11039);
xnor U11394 (N_11394,N_10824,N_10802);
nand U11395 (N_11395,N_11070,N_10929);
or U11396 (N_11396,N_10988,N_10927);
xnor U11397 (N_11397,N_10950,N_10820);
nand U11398 (N_11398,N_11010,N_11003);
and U11399 (N_11399,N_10888,N_10807);
xor U11400 (N_11400,N_11297,N_11303);
nor U11401 (N_11401,N_11395,N_11361);
nor U11402 (N_11402,N_11381,N_11370);
and U11403 (N_11403,N_11138,N_11274);
nand U11404 (N_11404,N_11286,N_11136);
nor U11405 (N_11405,N_11283,N_11252);
and U11406 (N_11406,N_11238,N_11234);
and U11407 (N_11407,N_11383,N_11174);
nor U11408 (N_11408,N_11233,N_11117);
xor U11409 (N_11409,N_11363,N_11251);
or U11410 (N_11410,N_11351,N_11280);
or U11411 (N_11411,N_11256,N_11154);
nand U11412 (N_11412,N_11108,N_11336);
and U11413 (N_11413,N_11321,N_11359);
xor U11414 (N_11414,N_11319,N_11206);
or U11415 (N_11415,N_11374,N_11307);
nor U11416 (N_11416,N_11196,N_11128);
nor U11417 (N_11417,N_11120,N_11171);
nor U11418 (N_11418,N_11141,N_11343);
and U11419 (N_11419,N_11394,N_11158);
and U11420 (N_11420,N_11342,N_11105);
xor U11421 (N_11421,N_11115,N_11201);
nand U11422 (N_11422,N_11209,N_11130);
nand U11423 (N_11423,N_11241,N_11191);
and U11424 (N_11424,N_11228,N_11194);
nand U11425 (N_11425,N_11264,N_11239);
xnor U11426 (N_11426,N_11382,N_11355);
or U11427 (N_11427,N_11184,N_11119);
nand U11428 (N_11428,N_11213,N_11326);
nor U11429 (N_11429,N_11155,N_11334);
and U11430 (N_11430,N_11293,N_11193);
xor U11431 (N_11431,N_11327,N_11306);
and U11432 (N_11432,N_11204,N_11371);
nor U11433 (N_11433,N_11142,N_11160);
nor U11434 (N_11434,N_11183,N_11311);
xnor U11435 (N_11435,N_11110,N_11161);
xnor U11436 (N_11436,N_11388,N_11353);
nor U11437 (N_11437,N_11302,N_11169);
xnor U11438 (N_11438,N_11140,N_11111);
nor U11439 (N_11439,N_11122,N_11102);
nor U11440 (N_11440,N_11377,N_11159);
nand U11441 (N_11441,N_11348,N_11369);
or U11442 (N_11442,N_11247,N_11282);
nand U11443 (N_11443,N_11143,N_11266);
nand U11444 (N_11444,N_11253,N_11254);
or U11445 (N_11445,N_11230,N_11118);
and U11446 (N_11446,N_11344,N_11367);
and U11447 (N_11447,N_11277,N_11269);
and U11448 (N_11448,N_11273,N_11203);
nand U11449 (N_11449,N_11229,N_11219);
xor U11450 (N_11450,N_11322,N_11275);
nand U11451 (N_11451,N_11153,N_11179);
xnor U11452 (N_11452,N_11245,N_11346);
nand U11453 (N_11453,N_11259,N_11258);
or U11454 (N_11454,N_11166,N_11398);
nand U11455 (N_11455,N_11231,N_11340);
or U11456 (N_11456,N_11187,N_11197);
or U11457 (N_11457,N_11341,N_11216);
nor U11458 (N_11458,N_11250,N_11123);
and U11459 (N_11459,N_11390,N_11214);
nand U11460 (N_11460,N_11185,N_11320);
or U11461 (N_11461,N_11354,N_11207);
xnor U11462 (N_11462,N_11223,N_11186);
nor U11463 (N_11463,N_11132,N_11202);
nand U11464 (N_11464,N_11150,N_11385);
nand U11465 (N_11465,N_11272,N_11325);
and U11466 (N_11466,N_11249,N_11284);
xnor U11467 (N_11467,N_11106,N_11198);
nand U11468 (N_11468,N_11267,N_11181);
or U11469 (N_11469,N_11396,N_11255);
nor U11470 (N_11470,N_11188,N_11289);
nand U11471 (N_11471,N_11350,N_11215);
or U11472 (N_11472,N_11335,N_11152);
and U11473 (N_11473,N_11205,N_11107);
or U11474 (N_11474,N_11232,N_11177);
nor U11475 (N_11475,N_11162,N_11244);
xor U11476 (N_11476,N_11109,N_11295);
and U11477 (N_11477,N_11133,N_11313);
xor U11478 (N_11478,N_11349,N_11263);
nand U11479 (N_11479,N_11278,N_11195);
nand U11480 (N_11480,N_11113,N_11240);
xnor U11481 (N_11481,N_11182,N_11131);
nand U11482 (N_11482,N_11242,N_11305);
and U11483 (N_11483,N_11391,N_11208);
and U11484 (N_11484,N_11221,N_11200);
nand U11485 (N_11485,N_11288,N_11121);
nor U11486 (N_11486,N_11165,N_11285);
nor U11487 (N_11487,N_11309,N_11294);
and U11488 (N_11488,N_11199,N_11366);
xor U11489 (N_11489,N_11290,N_11308);
or U11490 (N_11490,N_11149,N_11301);
xnor U11491 (N_11491,N_11167,N_11147);
nand U11492 (N_11492,N_11243,N_11246);
xor U11493 (N_11493,N_11339,N_11129);
nor U11494 (N_11494,N_11368,N_11237);
nor U11495 (N_11495,N_11324,N_11338);
xor U11496 (N_11496,N_11314,N_11330);
nor U11497 (N_11497,N_11298,N_11218);
or U11498 (N_11498,N_11172,N_11137);
or U11499 (N_11499,N_11329,N_11281);
nand U11500 (N_11500,N_11127,N_11164);
or U11501 (N_11501,N_11360,N_11227);
xor U11502 (N_11502,N_11176,N_11151);
xor U11503 (N_11503,N_11101,N_11210);
or U11504 (N_11504,N_11226,N_11260);
and U11505 (N_11505,N_11271,N_11386);
nand U11506 (N_11506,N_11399,N_11144);
xnor U11507 (N_11507,N_11393,N_11362);
nand U11508 (N_11508,N_11296,N_11318);
xnor U11509 (N_11509,N_11392,N_11261);
nand U11510 (N_11510,N_11389,N_11291);
and U11511 (N_11511,N_11315,N_11316);
nor U11512 (N_11512,N_11332,N_11178);
nand U11513 (N_11513,N_11379,N_11265);
nor U11514 (N_11514,N_11358,N_11257);
nor U11515 (N_11515,N_11365,N_11212);
nor U11516 (N_11516,N_11114,N_11262);
xnor U11517 (N_11517,N_11268,N_11135);
xor U11518 (N_11518,N_11323,N_11190);
nand U11519 (N_11519,N_11248,N_11299);
xnor U11520 (N_11520,N_11125,N_11337);
xnor U11521 (N_11521,N_11170,N_11364);
and U11522 (N_11522,N_11372,N_11376);
nand U11523 (N_11523,N_11116,N_11126);
or U11524 (N_11524,N_11189,N_11145);
and U11525 (N_11525,N_11112,N_11387);
nor U11526 (N_11526,N_11192,N_11270);
nor U11527 (N_11527,N_11304,N_11373);
or U11528 (N_11528,N_11378,N_11173);
or U11529 (N_11529,N_11312,N_11375);
nor U11530 (N_11530,N_11146,N_11276);
nand U11531 (N_11531,N_11397,N_11287);
nand U11532 (N_11532,N_11220,N_11134);
or U11533 (N_11533,N_11225,N_11317);
and U11534 (N_11534,N_11100,N_11222);
or U11535 (N_11535,N_11333,N_11380);
xnor U11536 (N_11536,N_11347,N_11163);
nor U11537 (N_11537,N_11310,N_11157);
and U11538 (N_11538,N_11356,N_11175);
and U11539 (N_11539,N_11224,N_11292);
or U11540 (N_11540,N_11345,N_11168);
and U11541 (N_11541,N_11217,N_11384);
nand U11542 (N_11542,N_11180,N_11279);
or U11543 (N_11543,N_11148,N_11328);
nand U11544 (N_11544,N_11104,N_11235);
nand U11545 (N_11545,N_11236,N_11211);
xnor U11546 (N_11546,N_11300,N_11139);
xnor U11547 (N_11547,N_11156,N_11124);
or U11548 (N_11548,N_11103,N_11331);
nor U11549 (N_11549,N_11357,N_11352);
nor U11550 (N_11550,N_11314,N_11285);
nor U11551 (N_11551,N_11221,N_11308);
and U11552 (N_11552,N_11141,N_11291);
nor U11553 (N_11553,N_11270,N_11228);
nand U11554 (N_11554,N_11293,N_11218);
nor U11555 (N_11555,N_11213,N_11283);
nand U11556 (N_11556,N_11139,N_11124);
nor U11557 (N_11557,N_11137,N_11312);
or U11558 (N_11558,N_11123,N_11300);
nor U11559 (N_11559,N_11247,N_11392);
nor U11560 (N_11560,N_11117,N_11395);
or U11561 (N_11561,N_11228,N_11366);
xnor U11562 (N_11562,N_11213,N_11137);
nor U11563 (N_11563,N_11292,N_11166);
or U11564 (N_11564,N_11208,N_11262);
and U11565 (N_11565,N_11356,N_11212);
or U11566 (N_11566,N_11166,N_11176);
xnor U11567 (N_11567,N_11284,N_11261);
nand U11568 (N_11568,N_11227,N_11316);
nand U11569 (N_11569,N_11367,N_11365);
xnor U11570 (N_11570,N_11279,N_11208);
nor U11571 (N_11571,N_11324,N_11315);
or U11572 (N_11572,N_11265,N_11164);
nand U11573 (N_11573,N_11362,N_11377);
nor U11574 (N_11574,N_11312,N_11320);
or U11575 (N_11575,N_11121,N_11144);
nor U11576 (N_11576,N_11240,N_11151);
nor U11577 (N_11577,N_11276,N_11387);
nor U11578 (N_11578,N_11139,N_11383);
nand U11579 (N_11579,N_11256,N_11272);
or U11580 (N_11580,N_11383,N_11130);
nor U11581 (N_11581,N_11163,N_11311);
nand U11582 (N_11582,N_11399,N_11280);
and U11583 (N_11583,N_11122,N_11244);
nand U11584 (N_11584,N_11311,N_11263);
and U11585 (N_11585,N_11232,N_11204);
or U11586 (N_11586,N_11140,N_11300);
nand U11587 (N_11587,N_11120,N_11251);
and U11588 (N_11588,N_11107,N_11277);
nand U11589 (N_11589,N_11212,N_11154);
nand U11590 (N_11590,N_11296,N_11188);
and U11591 (N_11591,N_11344,N_11333);
and U11592 (N_11592,N_11232,N_11200);
xor U11593 (N_11593,N_11358,N_11283);
nand U11594 (N_11594,N_11148,N_11202);
and U11595 (N_11595,N_11255,N_11368);
xor U11596 (N_11596,N_11306,N_11349);
xnor U11597 (N_11597,N_11145,N_11356);
nor U11598 (N_11598,N_11288,N_11357);
nand U11599 (N_11599,N_11386,N_11245);
and U11600 (N_11600,N_11308,N_11196);
nor U11601 (N_11601,N_11357,N_11259);
or U11602 (N_11602,N_11224,N_11284);
or U11603 (N_11603,N_11325,N_11112);
and U11604 (N_11604,N_11336,N_11338);
and U11605 (N_11605,N_11221,N_11309);
and U11606 (N_11606,N_11165,N_11200);
xor U11607 (N_11607,N_11178,N_11186);
nor U11608 (N_11608,N_11158,N_11194);
and U11609 (N_11609,N_11366,N_11359);
xor U11610 (N_11610,N_11330,N_11128);
and U11611 (N_11611,N_11390,N_11367);
xnor U11612 (N_11612,N_11187,N_11266);
nand U11613 (N_11613,N_11380,N_11271);
nand U11614 (N_11614,N_11363,N_11270);
and U11615 (N_11615,N_11223,N_11189);
nand U11616 (N_11616,N_11169,N_11205);
or U11617 (N_11617,N_11260,N_11202);
nand U11618 (N_11618,N_11280,N_11358);
nand U11619 (N_11619,N_11346,N_11196);
nor U11620 (N_11620,N_11178,N_11176);
nor U11621 (N_11621,N_11163,N_11165);
xor U11622 (N_11622,N_11358,N_11162);
nor U11623 (N_11623,N_11121,N_11320);
nor U11624 (N_11624,N_11389,N_11315);
and U11625 (N_11625,N_11305,N_11168);
nor U11626 (N_11626,N_11190,N_11321);
nor U11627 (N_11627,N_11382,N_11197);
or U11628 (N_11628,N_11273,N_11294);
nand U11629 (N_11629,N_11366,N_11394);
and U11630 (N_11630,N_11113,N_11100);
or U11631 (N_11631,N_11351,N_11199);
and U11632 (N_11632,N_11152,N_11282);
xnor U11633 (N_11633,N_11104,N_11277);
or U11634 (N_11634,N_11266,N_11224);
nor U11635 (N_11635,N_11156,N_11134);
and U11636 (N_11636,N_11172,N_11192);
xnor U11637 (N_11637,N_11341,N_11370);
xor U11638 (N_11638,N_11381,N_11192);
and U11639 (N_11639,N_11201,N_11136);
xor U11640 (N_11640,N_11376,N_11275);
xor U11641 (N_11641,N_11272,N_11193);
nand U11642 (N_11642,N_11146,N_11240);
or U11643 (N_11643,N_11113,N_11371);
nand U11644 (N_11644,N_11171,N_11206);
xor U11645 (N_11645,N_11265,N_11276);
or U11646 (N_11646,N_11390,N_11219);
and U11647 (N_11647,N_11175,N_11314);
nand U11648 (N_11648,N_11242,N_11340);
and U11649 (N_11649,N_11139,N_11120);
and U11650 (N_11650,N_11105,N_11398);
and U11651 (N_11651,N_11112,N_11277);
xor U11652 (N_11652,N_11263,N_11336);
nor U11653 (N_11653,N_11317,N_11248);
nor U11654 (N_11654,N_11327,N_11335);
and U11655 (N_11655,N_11362,N_11207);
nor U11656 (N_11656,N_11201,N_11346);
xnor U11657 (N_11657,N_11205,N_11324);
or U11658 (N_11658,N_11152,N_11135);
or U11659 (N_11659,N_11228,N_11243);
xor U11660 (N_11660,N_11174,N_11237);
or U11661 (N_11661,N_11239,N_11270);
xnor U11662 (N_11662,N_11176,N_11386);
nand U11663 (N_11663,N_11388,N_11306);
nand U11664 (N_11664,N_11184,N_11120);
or U11665 (N_11665,N_11349,N_11288);
and U11666 (N_11666,N_11205,N_11297);
nor U11667 (N_11667,N_11148,N_11308);
nand U11668 (N_11668,N_11331,N_11215);
xor U11669 (N_11669,N_11154,N_11359);
or U11670 (N_11670,N_11265,N_11250);
and U11671 (N_11671,N_11277,N_11166);
and U11672 (N_11672,N_11347,N_11199);
and U11673 (N_11673,N_11132,N_11206);
nand U11674 (N_11674,N_11327,N_11311);
nor U11675 (N_11675,N_11320,N_11248);
nor U11676 (N_11676,N_11218,N_11165);
nor U11677 (N_11677,N_11155,N_11276);
and U11678 (N_11678,N_11321,N_11322);
nor U11679 (N_11679,N_11202,N_11104);
or U11680 (N_11680,N_11371,N_11353);
xnor U11681 (N_11681,N_11163,N_11287);
xnor U11682 (N_11682,N_11112,N_11138);
or U11683 (N_11683,N_11351,N_11379);
nand U11684 (N_11684,N_11185,N_11354);
nand U11685 (N_11685,N_11192,N_11324);
nand U11686 (N_11686,N_11249,N_11314);
or U11687 (N_11687,N_11210,N_11337);
nor U11688 (N_11688,N_11235,N_11220);
xnor U11689 (N_11689,N_11208,N_11360);
and U11690 (N_11690,N_11390,N_11298);
xnor U11691 (N_11691,N_11279,N_11351);
and U11692 (N_11692,N_11134,N_11357);
xnor U11693 (N_11693,N_11200,N_11207);
or U11694 (N_11694,N_11147,N_11134);
xor U11695 (N_11695,N_11229,N_11214);
or U11696 (N_11696,N_11377,N_11231);
nand U11697 (N_11697,N_11371,N_11303);
nor U11698 (N_11698,N_11362,N_11214);
xnor U11699 (N_11699,N_11145,N_11387);
xnor U11700 (N_11700,N_11656,N_11473);
nand U11701 (N_11701,N_11419,N_11447);
and U11702 (N_11702,N_11658,N_11558);
and U11703 (N_11703,N_11482,N_11483);
nand U11704 (N_11704,N_11415,N_11510);
nor U11705 (N_11705,N_11580,N_11521);
nor U11706 (N_11706,N_11696,N_11573);
and U11707 (N_11707,N_11631,N_11517);
or U11708 (N_11708,N_11461,N_11405);
nand U11709 (N_11709,N_11552,N_11684);
xor U11710 (N_11710,N_11470,N_11424);
nand U11711 (N_11711,N_11599,N_11548);
nor U11712 (N_11712,N_11619,N_11591);
xnor U11713 (N_11713,N_11571,N_11425);
nor U11714 (N_11714,N_11423,N_11603);
nor U11715 (N_11715,N_11481,N_11633);
xor U11716 (N_11716,N_11575,N_11453);
or U11717 (N_11717,N_11454,N_11437);
nor U11718 (N_11718,N_11641,N_11478);
xor U11719 (N_11719,N_11611,N_11653);
nand U11720 (N_11720,N_11593,N_11418);
or U11721 (N_11721,N_11597,N_11568);
nor U11722 (N_11722,N_11657,N_11460);
and U11723 (N_11723,N_11496,N_11432);
nand U11724 (N_11724,N_11673,N_11562);
nor U11725 (N_11725,N_11636,N_11649);
nand U11726 (N_11726,N_11678,N_11578);
or U11727 (N_11727,N_11477,N_11472);
nor U11728 (N_11728,N_11550,N_11404);
nand U11729 (N_11729,N_11488,N_11539);
xor U11730 (N_11730,N_11540,N_11694);
xnor U11731 (N_11731,N_11479,N_11601);
nor U11732 (N_11732,N_11566,N_11624);
nand U11733 (N_11733,N_11574,N_11588);
and U11734 (N_11734,N_11498,N_11639);
nor U11735 (N_11735,N_11468,N_11660);
and U11736 (N_11736,N_11598,N_11590);
nor U11737 (N_11737,N_11589,N_11449);
nand U11738 (N_11738,N_11541,N_11495);
xnor U11739 (N_11739,N_11570,N_11665);
and U11740 (N_11740,N_11697,N_11625);
and U11741 (N_11741,N_11687,N_11560);
xnor U11742 (N_11742,N_11576,N_11497);
nand U11743 (N_11743,N_11563,N_11690);
nand U11744 (N_11744,N_11484,N_11620);
or U11745 (N_11745,N_11466,N_11410);
nand U11746 (N_11746,N_11531,N_11503);
nor U11747 (N_11747,N_11606,N_11522);
and U11748 (N_11748,N_11676,N_11512);
or U11749 (N_11749,N_11680,N_11544);
xnor U11750 (N_11750,N_11400,N_11529);
xor U11751 (N_11751,N_11407,N_11693);
xnor U11752 (N_11752,N_11485,N_11632);
and U11753 (N_11753,N_11507,N_11450);
xor U11754 (N_11754,N_11621,N_11448);
xor U11755 (N_11755,N_11523,N_11698);
or U11756 (N_11756,N_11644,N_11586);
xor U11757 (N_11757,N_11467,N_11542);
nand U11758 (N_11758,N_11637,N_11567);
or U11759 (N_11759,N_11408,N_11608);
or U11760 (N_11760,N_11577,N_11465);
nand U11761 (N_11761,N_11416,N_11643);
and U11762 (N_11762,N_11431,N_11582);
nor U11763 (N_11763,N_11434,N_11555);
or U11764 (N_11764,N_11647,N_11505);
or U11765 (N_11765,N_11442,N_11452);
and U11766 (N_11766,N_11439,N_11602);
nand U11767 (N_11767,N_11520,N_11493);
nand U11768 (N_11768,N_11534,N_11671);
and U11769 (N_11769,N_11422,N_11436);
nor U11770 (N_11770,N_11545,N_11682);
nand U11771 (N_11771,N_11561,N_11516);
xnor U11772 (N_11772,N_11699,N_11683);
nand U11773 (N_11773,N_11646,N_11557);
and U11774 (N_11774,N_11451,N_11413);
and U11775 (N_11775,N_11519,N_11463);
and U11776 (N_11776,N_11500,N_11513);
xnor U11777 (N_11777,N_11622,N_11536);
and U11778 (N_11778,N_11433,N_11675);
and U11779 (N_11779,N_11648,N_11421);
nor U11780 (N_11780,N_11506,N_11514);
nor U11781 (N_11781,N_11492,N_11695);
or U11782 (N_11782,N_11677,N_11650);
or U11783 (N_11783,N_11501,N_11672);
nand U11784 (N_11784,N_11596,N_11428);
or U11785 (N_11785,N_11471,N_11614);
or U11786 (N_11786,N_11579,N_11455);
and U11787 (N_11787,N_11547,N_11426);
or U11788 (N_11788,N_11659,N_11654);
or U11789 (N_11789,N_11628,N_11435);
nand U11790 (N_11790,N_11564,N_11689);
nor U11791 (N_11791,N_11612,N_11685);
nor U11792 (N_11792,N_11499,N_11559);
nor U11793 (N_11793,N_11670,N_11508);
xor U11794 (N_11794,N_11487,N_11525);
or U11795 (N_11795,N_11615,N_11686);
and U11796 (N_11796,N_11556,N_11688);
xnor U11797 (N_11797,N_11651,N_11592);
nor U11798 (N_11798,N_11515,N_11652);
xnor U11799 (N_11799,N_11551,N_11618);
nand U11800 (N_11800,N_11475,N_11669);
and U11801 (N_11801,N_11509,N_11610);
and U11802 (N_11802,N_11494,N_11402);
and U11803 (N_11803,N_11462,N_11655);
nand U11804 (N_11804,N_11480,N_11569);
nand U11805 (N_11805,N_11617,N_11663);
nor U11806 (N_11806,N_11429,N_11518);
nand U11807 (N_11807,N_11661,N_11604);
nor U11808 (N_11808,N_11681,N_11464);
or U11809 (N_11809,N_11430,N_11444);
nand U11810 (N_11810,N_11489,N_11443);
nor U11811 (N_11811,N_11585,N_11613);
and U11812 (N_11812,N_11533,N_11511);
nor U11813 (N_11813,N_11490,N_11459);
or U11814 (N_11814,N_11630,N_11546);
and U11815 (N_11815,N_11565,N_11491);
nand U11816 (N_11816,N_11412,N_11524);
xnor U11817 (N_11817,N_11623,N_11474);
xor U11818 (N_11818,N_11581,N_11530);
and U11819 (N_11819,N_11420,N_11666);
and U11820 (N_11820,N_11645,N_11664);
nor U11821 (N_11821,N_11458,N_11427);
nor U11822 (N_11822,N_11629,N_11456);
xnor U11823 (N_11823,N_11406,N_11554);
xnor U11824 (N_11824,N_11627,N_11616);
nand U11825 (N_11825,N_11595,N_11609);
and U11826 (N_11826,N_11692,N_11457);
nor U11827 (N_11827,N_11640,N_11583);
nand U11828 (N_11828,N_11642,N_11440);
nor U11829 (N_11829,N_11553,N_11662);
xnor U11830 (N_11830,N_11409,N_11527);
or U11831 (N_11831,N_11607,N_11635);
nand U11832 (N_11832,N_11532,N_11401);
and U11833 (N_11833,N_11667,N_11638);
nand U11834 (N_11834,N_11537,N_11543);
and U11835 (N_11835,N_11668,N_11438);
nand U11836 (N_11836,N_11502,N_11446);
xnor U11837 (N_11837,N_11605,N_11403);
or U11838 (N_11838,N_11584,N_11528);
nor U11839 (N_11839,N_11535,N_11441);
nand U11840 (N_11840,N_11526,N_11445);
nor U11841 (N_11841,N_11538,N_11504);
nand U11842 (N_11842,N_11600,N_11549);
xor U11843 (N_11843,N_11587,N_11486);
and U11844 (N_11844,N_11674,N_11634);
nand U11845 (N_11845,N_11417,N_11469);
nor U11846 (N_11846,N_11414,N_11679);
and U11847 (N_11847,N_11411,N_11691);
and U11848 (N_11848,N_11572,N_11626);
and U11849 (N_11849,N_11476,N_11594);
or U11850 (N_11850,N_11640,N_11599);
nand U11851 (N_11851,N_11628,N_11578);
nor U11852 (N_11852,N_11491,N_11609);
xnor U11853 (N_11853,N_11530,N_11452);
nor U11854 (N_11854,N_11501,N_11449);
nand U11855 (N_11855,N_11606,N_11647);
or U11856 (N_11856,N_11485,N_11435);
nand U11857 (N_11857,N_11499,N_11631);
and U11858 (N_11858,N_11655,N_11681);
and U11859 (N_11859,N_11443,N_11520);
nand U11860 (N_11860,N_11507,N_11542);
nor U11861 (N_11861,N_11627,N_11619);
or U11862 (N_11862,N_11671,N_11400);
nor U11863 (N_11863,N_11578,N_11539);
nand U11864 (N_11864,N_11625,N_11524);
or U11865 (N_11865,N_11520,N_11401);
nand U11866 (N_11866,N_11628,N_11658);
nor U11867 (N_11867,N_11536,N_11614);
and U11868 (N_11868,N_11410,N_11522);
xnor U11869 (N_11869,N_11424,N_11560);
xnor U11870 (N_11870,N_11464,N_11439);
and U11871 (N_11871,N_11641,N_11565);
and U11872 (N_11872,N_11538,N_11512);
or U11873 (N_11873,N_11530,N_11560);
nand U11874 (N_11874,N_11458,N_11483);
or U11875 (N_11875,N_11519,N_11498);
nor U11876 (N_11876,N_11414,N_11682);
nand U11877 (N_11877,N_11475,N_11400);
and U11878 (N_11878,N_11626,N_11430);
and U11879 (N_11879,N_11655,N_11639);
xor U11880 (N_11880,N_11505,N_11544);
xor U11881 (N_11881,N_11613,N_11473);
nor U11882 (N_11882,N_11483,N_11576);
xnor U11883 (N_11883,N_11425,N_11494);
nand U11884 (N_11884,N_11409,N_11509);
xor U11885 (N_11885,N_11642,N_11509);
nor U11886 (N_11886,N_11601,N_11491);
or U11887 (N_11887,N_11452,N_11467);
nor U11888 (N_11888,N_11549,N_11478);
nand U11889 (N_11889,N_11568,N_11406);
nand U11890 (N_11890,N_11455,N_11422);
and U11891 (N_11891,N_11601,N_11677);
xor U11892 (N_11892,N_11463,N_11516);
nor U11893 (N_11893,N_11648,N_11577);
nand U11894 (N_11894,N_11503,N_11647);
nand U11895 (N_11895,N_11404,N_11681);
nand U11896 (N_11896,N_11597,N_11409);
nor U11897 (N_11897,N_11612,N_11482);
xnor U11898 (N_11898,N_11526,N_11580);
nand U11899 (N_11899,N_11561,N_11552);
nor U11900 (N_11900,N_11520,N_11606);
or U11901 (N_11901,N_11406,N_11546);
xnor U11902 (N_11902,N_11421,N_11466);
nor U11903 (N_11903,N_11534,N_11589);
nand U11904 (N_11904,N_11633,N_11636);
and U11905 (N_11905,N_11661,N_11594);
nand U11906 (N_11906,N_11417,N_11698);
and U11907 (N_11907,N_11472,N_11693);
nand U11908 (N_11908,N_11448,N_11525);
and U11909 (N_11909,N_11543,N_11419);
xnor U11910 (N_11910,N_11414,N_11538);
xnor U11911 (N_11911,N_11456,N_11457);
nand U11912 (N_11912,N_11603,N_11619);
xor U11913 (N_11913,N_11518,N_11531);
xor U11914 (N_11914,N_11647,N_11438);
and U11915 (N_11915,N_11567,N_11540);
nor U11916 (N_11916,N_11608,N_11524);
or U11917 (N_11917,N_11469,N_11489);
nand U11918 (N_11918,N_11509,N_11518);
and U11919 (N_11919,N_11417,N_11557);
or U11920 (N_11920,N_11575,N_11447);
nor U11921 (N_11921,N_11402,N_11556);
nand U11922 (N_11922,N_11603,N_11475);
xor U11923 (N_11923,N_11639,N_11688);
nand U11924 (N_11924,N_11419,N_11407);
or U11925 (N_11925,N_11665,N_11657);
nand U11926 (N_11926,N_11405,N_11603);
and U11927 (N_11927,N_11538,N_11557);
nand U11928 (N_11928,N_11525,N_11674);
nand U11929 (N_11929,N_11490,N_11542);
xor U11930 (N_11930,N_11558,N_11429);
xor U11931 (N_11931,N_11492,N_11633);
nand U11932 (N_11932,N_11645,N_11468);
or U11933 (N_11933,N_11627,N_11493);
or U11934 (N_11934,N_11606,N_11508);
xnor U11935 (N_11935,N_11697,N_11683);
xnor U11936 (N_11936,N_11588,N_11431);
nor U11937 (N_11937,N_11465,N_11695);
xnor U11938 (N_11938,N_11523,N_11674);
xnor U11939 (N_11939,N_11491,N_11603);
or U11940 (N_11940,N_11454,N_11650);
and U11941 (N_11941,N_11474,N_11486);
or U11942 (N_11942,N_11668,N_11510);
xnor U11943 (N_11943,N_11453,N_11580);
nand U11944 (N_11944,N_11462,N_11454);
nand U11945 (N_11945,N_11678,N_11671);
xnor U11946 (N_11946,N_11573,N_11626);
and U11947 (N_11947,N_11668,N_11412);
nand U11948 (N_11948,N_11554,N_11562);
xor U11949 (N_11949,N_11456,N_11536);
xor U11950 (N_11950,N_11678,N_11679);
or U11951 (N_11951,N_11448,N_11566);
xnor U11952 (N_11952,N_11668,N_11415);
nor U11953 (N_11953,N_11460,N_11420);
nand U11954 (N_11954,N_11408,N_11416);
nand U11955 (N_11955,N_11427,N_11691);
nand U11956 (N_11956,N_11484,N_11605);
and U11957 (N_11957,N_11518,N_11512);
nand U11958 (N_11958,N_11402,N_11492);
or U11959 (N_11959,N_11638,N_11517);
xor U11960 (N_11960,N_11563,N_11448);
xor U11961 (N_11961,N_11433,N_11490);
xnor U11962 (N_11962,N_11680,N_11589);
and U11963 (N_11963,N_11529,N_11651);
xnor U11964 (N_11964,N_11646,N_11484);
or U11965 (N_11965,N_11615,N_11506);
nand U11966 (N_11966,N_11670,N_11565);
xor U11967 (N_11967,N_11481,N_11569);
nor U11968 (N_11968,N_11432,N_11438);
or U11969 (N_11969,N_11459,N_11534);
xor U11970 (N_11970,N_11577,N_11451);
nor U11971 (N_11971,N_11699,N_11514);
nor U11972 (N_11972,N_11420,N_11520);
xnor U11973 (N_11973,N_11694,N_11642);
nor U11974 (N_11974,N_11698,N_11637);
nor U11975 (N_11975,N_11645,N_11515);
or U11976 (N_11976,N_11567,N_11465);
xnor U11977 (N_11977,N_11605,N_11634);
xor U11978 (N_11978,N_11534,N_11568);
xor U11979 (N_11979,N_11609,N_11463);
or U11980 (N_11980,N_11610,N_11539);
xnor U11981 (N_11981,N_11644,N_11530);
nor U11982 (N_11982,N_11482,N_11520);
nand U11983 (N_11983,N_11691,N_11486);
or U11984 (N_11984,N_11663,N_11407);
nand U11985 (N_11985,N_11579,N_11430);
and U11986 (N_11986,N_11439,N_11470);
nor U11987 (N_11987,N_11698,N_11588);
and U11988 (N_11988,N_11546,N_11604);
nand U11989 (N_11989,N_11603,N_11502);
nand U11990 (N_11990,N_11600,N_11540);
xnor U11991 (N_11991,N_11645,N_11462);
and U11992 (N_11992,N_11428,N_11677);
nand U11993 (N_11993,N_11544,N_11416);
xnor U11994 (N_11994,N_11406,N_11512);
and U11995 (N_11995,N_11694,N_11568);
and U11996 (N_11996,N_11586,N_11453);
nor U11997 (N_11997,N_11507,N_11690);
nand U11998 (N_11998,N_11606,N_11566);
nor U11999 (N_11999,N_11699,N_11569);
or U12000 (N_12000,N_11765,N_11901);
nand U12001 (N_12001,N_11742,N_11813);
or U12002 (N_12002,N_11754,N_11888);
or U12003 (N_12003,N_11810,N_11815);
xor U12004 (N_12004,N_11811,N_11749);
or U12005 (N_12005,N_11827,N_11971);
xor U12006 (N_12006,N_11764,N_11892);
or U12007 (N_12007,N_11798,N_11862);
nor U12008 (N_12008,N_11883,N_11780);
and U12009 (N_12009,N_11936,N_11783);
and U12010 (N_12010,N_11807,N_11730);
xor U12011 (N_12011,N_11766,N_11791);
nor U12012 (N_12012,N_11816,N_11882);
xnor U12013 (N_12013,N_11894,N_11880);
or U12014 (N_12014,N_11729,N_11781);
nand U12015 (N_12015,N_11714,N_11757);
xnor U12016 (N_12016,N_11859,N_11831);
xnor U12017 (N_12017,N_11863,N_11884);
xnor U12018 (N_12018,N_11899,N_11994);
or U12019 (N_12019,N_11785,N_11981);
xor U12020 (N_12020,N_11896,N_11715);
and U12021 (N_12021,N_11837,N_11910);
or U12022 (N_12022,N_11747,N_11849);
and U12023 (N_12023,N_11728,N_11777);
nand U12024 (N_12024,N_11900,N_11871);
nand U12025 (N_12025,N_11858,N_11834);
nand U12026 (N_12026,N_11977,N_11952);
or U12027 (N_12027,N_11890,N_11943);
and U12028 (N_12028,N_11778,N_11756);
xor U12029 (N_12029,N_11864,N_11857);
or U12030 (N_12030,N_11877,N_11794);
nand U12031 (N_12031,N_11948,N_11712);
nand U12032 (N_12032,N_11898,N_11741);
xor U12033 (N_12033,N_11821,N_11851);
or U12034 (N_12034,N_11760,N_11946);
and U12035 (N_12035,N_11972,N_11879);
nand U12036 (N_12036,N_11969,N_11845);
xor U12037 (N_12037,N_11724,N_11716);
nand U12038 (N_12038,N_11840,N_11875);
nor U12039 (N_12039,N_11993,N_11953);
xnor U12040 (N_12040,N_11842,N_11873);
nor U12041 (N_12041,N_11828,N_11839);
nor U12042 (N_12042,N_11999,N_11947);
or U12043 (N_12043,N_11922,N_11852);
and U12044 (N_12044,N_11767,N_11720);
and U12045 (N_12045,N_11793,N_11738);
xnor U12046 (N_12046,N_11867,N_11963);
nor U12047 (N_12047,N_11758,N_11819);
xnor U12048 (N_12048,N_11773,N_11796);
nor U12049 (N_12049,N_11872,N_11717);
or U12050 (N_12050,N_11995,N_11992);
nand U12051 (N_12051,N_11893,N_11700);
nor U12052 (N_12052,N_11824,N_11832);
xnor U12053 (N_12053,N_11823,N_11762);
and U12054 (N_12054,N_11833,N_11985);
and U12055 (N_12055,N_11753,N_11775);
nor U12056 (N_12056,N_11902,N_11903);
nand U12057 (N_12057,N_11782,N_11907);
or U12058 (N_12058,N_11869,N_11812);
nand U12059 (N_12059,N_11913,N_11960);
nor U12060 (N_12060,N_11743,N_11889);
nand U12061 (N_12061,N_11909,N_11841);
or U12062 (N_12062,N_11731,N_11966);
and U12063 (N_12063,N_11848,N_11850);
and U12064 (N_12064,N_11727,N_11725);
nand U12065 (N_12065,N_11853,N_11868);
and U12066 (N_12066,N_11957,N_11881);
or U12067 (N_12067,N_11708,N_11740);
nor U12068 (N_12068,N_11951,N_11751);
nor U12069 (N_12069,N_11870,N_11710);
nand U12070 (N_12070,N_11924,N_11918);
or U12071 (N_12071,N_11808,N_11925);
and U12072 (N_12072,N_11876,N_11788);
nand U12073 (N_12073,N_11745,N_11945);
xnor U12074 (N_12074,N_11790,N_11904);
nor U12075 (N_12075,N_11774,N_11784);
nand U12076 (N_12076,N_11949,N_11802);
nand U12077 (N_12077,N_11974,N_11961);
and U12078 (N_12078,N_11905,N_11734);
nand U12079 (N_12079,N_11755,N_11847);
or U12080 (N_12080,N_11826,N_11732);
or U12081 (N_12081,N_11886,N_11703);
and U12082 (N_12082,N_11804,N_11865);
or U12083 (N_12083,N_11706,N_11761);
nor U12084 (N_12084,N_11855,N_11926);
xnor U12085 (N_12085,N_11705,N_11895);
and U12086 (N_12086,N_11932,N_11934);
nand U12087 (N_12087,N_11805,N_11763);
nand U12088 (N_12088,N_11962,N_11702);
and U12089 (N_12089,N_11792,N_11983);
or U12090 (N_12090,N_11830,N_11861);
or U12091 (N_12091,N_11987,N_11944);
xnor U12092 (N_12092,N_11984,N_11744);
nand U12093 (N_12093,N_11990,N_11933);
nand U12094 (N_12094,N_11988,N_11954);
xor U12095 (N_12095,N_11776,N_11856);
and U12096 (N_12096,N_11935,N_11996);
and U12097 (N_12097,N_11941,N_11814);
nor U12098 (N_12098,N_11726,N_11860);
xor U12099 (N_12099,N_11719,N_11959);
and U12100 (N_12100,N_11975,N_11911);
nand U12101 (N_12101,N_11787,N_11797);
nand U12102 (N_12102,N_11940,N_11866);
or U12103 (N_12103,N_11739,N_11916);
xnor U12104 (N_12104,N_11736,N_11722);
nand U12105 (N_12105,N_11919,N_11942);
or U12106 (N_12106,N_11806,N_11750);
nor U12107 (N_12107,N_11908,N_11914);
nor U12108 (N_12108,N_11927,N_11772);
and U12109 (N_12109,N_11973,N_11920);
nand U12110 (N_12110,N_11836,N_11770);
nor U12111 (N_12111,N_11854,N_11829);
nor U12112 (N_12112,N_11733,N_11789);
or U12113 (N_12113,N_11878,N_11923);
or U12114 (N_12114,N_11906,N_11915);
xnor U12115 (N_12115,N_11759,N_11950);
nor U12116 (N_12116,N_11939,N_11980);
xor U12117 (N_12117,N_11769,N_11748);
nand U12118 (N_12118,N_11997,N_11885);
and U12119 (N_12119,N_11820,N_11709);
nand U12120 (N_12120,N_11818,N_11735);
and U12121 (N_12121,N_11917,N_11838);
nand U12122 (N_12122,N_11930,N_11978);
or U12123 (N_12123,N_11752,N_11912);
and U12124 (N_12124,N_11843,N_11795);
nand U12125 (N_12125,N_11737,N_11846);
nor U12126 (N_12126,N_11968,N_11723);
and U12127 (N_12127,N_11701,N_11825);
nor U12128 (N_12128,N_11970,N_11817);
nand U12129 (N_12129,N_11771,N_11801);
nor U12130 (N_12130,N_11989,N_11707);
and U12131 (N_12131,N_11965,N_11809);
nor U12132 (N_12132,N_11835,N_11897);
nor U12133 (N_12133,N_11822,N_11786);
and U12134 (N_12134,N_11991,N_11979);
xor U12135 (N_12135,N_11929,N_11928);
nand U12136 (N_12136,N_11967,N_11958);
and U12137 (N_12137,N_11976,N_11711);
nor U12138 (N_12138,N_11874,N_11891);
nor U12139 (N_12139,N_11887,N_11803);
nand U12140 (N_12140,N_11982,N_11986);
nor U12141 (N_12141,N_11938,N_11768);
xnor U12142 (N_12142,N_11956,N_11937);
or U12143 (N_12143,N_11779,N_11964);
nand U12144 (N_12144,N_11800,N_11721);
nand U12145 (N_12145,N_11998,N_11931);
nor U12146 (N_12146,N_11713,N_11718);
nor U12147 (N_12147,N_11799,N_11955);
or U12148 (N_12148,N_11921,N_11746);
nand U12149 (N_12149,N_11704,N_11844);
nand U12150 (N_12150,N_11837,N_11977);
xor U12151 (N_12151,N_11738,N_11863);
or U12152 (N_12152,N_11826,N_11715);
nor U12153 (N_12153,N_11872,N_11723);
xor U12154 (N_12154,N_11928,N_11719);
or U12155 (N_12155,N_11914,N_11904);
or U12156 (N_12156,N_11995,N_11775);
nand U12157 (N_12157,N_11853,N_11765);
xor U12158 (N_12158,N_11714,N_11940);
nand U12159 (N_12159,N_11924,N_11835);
or U12160 (N_12160,N_11701,N_11930);
xnor U12161 (N_12161,N_11989,N_11828);
or U12162 (N_12162,N_11700,N_11860);
nand U12163 (N_12163,N_11947,N_11863);
or U12164 (N_12164,N_11881,N_11964);
nand U12165 (N_12165,N_11929,N_11768);
nor U12166 (N_12166,N_11753,N_11951);
and U12167 (N_12167,N_11723,N_11729);
or U12168 (N_12168,N_11950,N_11948);
or U12169 (N_12169,N_11817,N_11902);
nand U12170 (N_12170,N_11716,N_11889);
or U12171 (N_12171,N_11935,N_11708);
nor U12172 (N_12172,N_11770,N_11864);
or U12173 (N_12173,N_11983,N_11815);
nor U12174 (N_12174,N_11919,N_11817);
nand U12175 (N_12175,N_11824,N_11948);
nand U12176 (N_12176,N_11913,N_11702);
or U12177 (N_12177,N_11987,N_11722);
xor U12178 (N_12178,N_11936,N_11901);
xnor U12179 (N_12179,N_11893,N_11912);
nor U12180 (N_12180,N_11800,N_11848);
xor U12181 (N_12181,N_11927,N_11900);
nor U12182 (N_12182,N_11869,N_11782);
and U12183 (N_12183,N_11880,N_11982);
or U12184 (N_12184,N_11778,N_11842);
xnor U12185 (N_12185,N_11942,N_11773);
or U12186 (N_12186,N_11894,N_11998);
nor U12187 (N_12187,N_11949,N_11892);
xnor U12188 (N_12188,N_11960,N_11881);
nor U12189 (N_12189,N_11787,N_11908);
and U12190 (N_12190,N_11701,N_11974);
nand U12191 (N_12191,N_11726,N_11834);
nand U12192 (N_12192,N_11908,N_11902);
nor U12193 (N_12193,N_11727,N_11823);
and U12194 (N_12194,N_11844,N_11784);
and U12195 (N_12195,N_11865,N_11961);
or U12196 (N_12196,N_11725,N_11723);
and U12197 (N_12197,N_11853,N_11757);
or U12198 (N_12198,N_11791,N_11821);
nor U12199 (N_12199,N_11757,N_11924);
nand U12200 (N_12200,N_11950,N_11775);
nor U12201 (N_12201,N_11822,N_11910);
and U12202 (N_12202,N_11995,N_11777);
xnor U12203 (N_12203,N_11938,N_11703);
and U12204 (N_12204,N_11944,N_11828);
or U12205 (N_12205,N_11965,N_11805);
nor U12206 (N_12206,N_11994,N_11848);
xor U12207 (N_12207,N_11883,N_11764);
nand U12208 (N_12208,N_11824,N_11827);
nand U12209 (N_12209,N_11843,N_11927);
nor U12210 (N_12210,N_11772,N_11985);
xnor U12211 (N_12211,N_11888,N_11782);
nand U12212 (N_12212,N_11941,N_11761);
or U12213 (N_12213,N_11836,N_11889);
and U12214 (N_12214,N_11860,N_11707);
nand U12215 (N_12215,N_11909,N_11788);
nand U12216 (N_12216,N_11787,N_11818);
and U12217 (N_12217,N_11993,N_11925);
xor U12218 (N_12218,N_11945,N_11982);
or U12219 (N_12219,N_11927,N_11780);
nor U12220 (N_12220,N_11743,N_11735);
xor U12221 (N_12221,N_11903,N_11835);
xor U12222 (N_12222,N_11746,N_11959);
nor U12223 (N_12223,N_11801,N_11957);
nand U12224 (N_12224,N_11988,N_11888);
nor U12225 (N_12225,N_11709,N_11770);
and U12226 (N_12226,N_11829,N_11778);
xor U12227 (N_12227,N_11852,N_11934);
and U12228 (N_12228,N_11911,N_11871);
nand U12229 (N_12229,N_11943,N_11965);
and U12230 (N_12230,N_11900,N_11843);
nor U12231 (N_12231,N_11838,N_11888);
nor U12232 (N_12232,N_11835,N_11925);
xor U12233 (N_12233,N_11972,N_11726);
and U12234 (N_12234,N_11833,N_11782);
nor U12235 (N_12235,N_11853,N_11743);
and U12236 (N_12236,N_11871,N_11964);
nand U12237 (N_12237,N_11999,N_11742);
and U12238 (N_12238,N_11893,N_11885);
and U12239 (N_12239,N_11931,N_11773);
xor U12240 (N_12240,N_11815,N_11830);
nand U12241 (N_12241,N_11870,N_11897);
or U12242 (N_12242,N_11851,N_11725);
nor U12243 (N_12243,N_11793,N_11978);
nand U12244 (N_12244,N_11911,N_11764);
and U12245 (N_12245,N_11745,N_11752);
and U12246 (N_12246,N_11889,N_11791);
or U12247 (N_12247,N_11856,N_11846);
nand U12248 (N_12248,N_11891,N_11983);
nand U12249 (N_12249,N_11719,N_11705);
nor U12250 (N_12250,N_11964,N_11823);
and U12251 (N_12251,N_11833,N_11944);
or U12252 (N_12252,N_11704,N_11854);
or U12253 (N_12253,N_11845,N_11916);
and U12254 (N_12254,N_11914,N_11946);
nand U12255 (N_12255,N_11801,N_11947);
or U12256 (N_12256,N_11845,N_11840);
nand U12257 (N_12257,N_11944,N_11951);
and U12258 (N_12258,N_11712,N_11809);
and U12259 (N_12259,N_11967,N_11711);
xnor U12260 (N_12260,N_11716,N_11762);
and U12261 (N_12261,N_11921,N_11820);
or U12262 (N_12262,N_11776,N_11874);
and U12263 (N_12263,N_11752,N_11832);
and U12264 (N_12264,N_11878,N_11748);
and U12265 (N_12265,N_11729,N_11985);
xnor U12266 (N_12266,N_11887,N_11806);
nand U12267 (N_12267,N_11741,N_11754);
nor U12268 (N_12268,N_11706,N_11959);
xnor U12269 (N_12269,N_11929,N_11957);
or U12270 (N_12270,N_11744,N_11848);
xnor U12271 (N_12271,N_11725,N_11874);
xor U12272 (N_12272,N_11709,N_11826);
or U12273 (N_12273,N_11774,N_11878);
xor U12274 (N_12274,N_11884,N_11773);
nand U12275 (N_12275,N_11836,N_11993);
nand U12276 (N_12276,N_11923,N_11937);
and U12277 (N_12277,N_11997,N_11715);
xnor U12278 (N_12278,N_11731,N_11748);
and U12279 (N_12279,N_11906,N_11877);
nor U12280 (N_12280,N_11851,N_11970);
nor U12281 (N_12281,N_11785,N_11942);
xor U12282 (N_12282,N_11739,N_11804);
and U12283 (N_12283,N_11968,N_11905);
nand U12284 (N_12284,N_11935,N_11979);
nand U12285 (N_12285,N_11909,N_11859);
xor U12286 (N_12286,N_11791,N_11723);
nand U12287 (N_12287,N_11870,N_11947);
xor U12288 (N_12288,N_11922,N_11788);
and U12289 (N_12289,N_11724,N_11893);
and U12290 (N_12290,N_11798,N_11724);
nand U12291 (N_12291,N_11868,N_11903);
xor U12292 (N_12292,N_11840,N_11876);
nand U12293 (N_12293,N_11759,N_11764);
nor U12294 (N_12294,N_11906,N_11969);
and U12295 (N_12295,N_11793,N_11999);
xnor U12296 (N_12296,N_11796,N_11983);
xor U12297 (N_12297,N_11836,N_11771);
nor U12298 (N_12298,N_11882,N_11910);
nand U12299 (N_12299,N_11735,N_11848);
and U12300 (N_12300,N_12124,N_12058);
xnor U12301 (N_12301,N_12051,N_12090);
nand U12302 (N_12302,N_12020,N_12096);
or U12303 (N_12303,N_12137,N_12221);
and U12304 (N_12304,N_12295,N_12179);
nand U12305 (N_12305,N_12046,N_12012);
nand U12306 (N_12306,N_12088,N_12174);
xor U12307 (N_12307,N_12173,N_12224);
or U12308 (N_12308,N_12119,N_12035);
xnor U12309 (N_12309,N_12198,N_12235);
nor U12310 (N_12310,N_12265,N_12134);
nor U12311 (N_12311,N_12187,N_12192);
nor U12312 (N_12312,N_12227,N_12209);
nor U12313 (N_12313,N_12256,N_12066);
nand U12314 (N_12314,N_12142,N_12052);
xnor U12315 (N_12315,N_12261,N_12118);
nor U12316 (N_12316,N_12022,N_12070);
nor U12317 (N_12317,N_12234,N_12128);
nand U12318 (N_12318,N_12230,N_12279);
or U12319 (N_12319,N_12037,N_12113);
xor U12320 (N_12320,N_12262,N_12018);
nand U12321 (N_12321,N_12283,N_12156);
nor U12322 (N_12322,N_12293,N_12285);
or U12323 (N_12323,N_12165,N_12087);
nand U12324 (N_12324,N_12040,N_12007);
xor U12325 (N_12325,N_12178,N_12114);
xnor U12326 (N_12326,N_12086,N_12299);
nor U12327 (N_12327,N_12218,N_12084);
xnor U12328 (N_12328,N_12225,N_12255);
or U12329 (N_12329,N_12250,N_12059);
or U12330 (N_12330,N_12145,N_12009);
xor U12331 (N_12331,N_12195,N_12243);
nand U12332 (N_12332,N_12238,N_12032);
and U12333 (N_12333,N_12122,N_12284);
nor U12334 (N_12334,N_12267,N_12212);
xor U12335 (N_12335,N_12213,N_12109);
nor U12336 (N_12336,N_12127,N_12260);
nor U12337 (N_12337,N_12002,N_12103);
nor U12338 (N_12338,N_12130,N_12199);
or U12339 (N_12339,N_12120,N_12186);
and U12340 (N_12340,N_12278,N_12148);
nor U12341 (N_12341,N_12141,N_12024);
and U12342 (N_12342,N_12085,N_12170);
and U12343 (N_12343,N_12194,N_12296);
nand U12344 (N_12344,N_12060,N_12294);
xnor U12345 (N_12345,N_12168,N_12044);
and U12346 (N_12346,N_12136,N_12143);
nand U12347 (N_12347,N_12244,N_12126);
and U12348 (N_12348,N_12251,N_12207);
or U12349 (N_12349,N_12107,N_12298);
xnor U12350 (N_12350,N_12117,N_12184);
nand U12351 (N_12351,N_12016,N_12031);
and U12352 (N_12352,N_12286,N_12079);
nor U12353 (N_12353,N_12264,N_12161);
and U12354 (N_12354,N_12001,N_12211);
or U12355 (N_12355,N_12166,N_12259);
xor U12356 (N_12356,N_12258,N_12006);
or U12357 (N_12357,N_12133,N_12280);
nor U12358 (N_12358,N_12281,N_12093);
xor U12359 (N_12359,N_12135,N_12236);
xor U12360 (N_12360,N_12138,N_12222);
and U12361 (N_12361,N_12078,N_12277);
xor U12362 (N_12362,N_12275,N_12241);
nand U12363 (N_12363,N_12062,N_12223);
xor U12364 (N_12364,N_12057,N_12248);
or U12365 (N_12365,N_12181,N_12038);
nand U12366 (N_12366,N_12152,N_12054);
nand U12367 (N_12367,N_12027,N_12067);
nor U12368 (N_12368,N_12131,N_12164);
and U12369 (N_12369,N_12081,N_12169);
and U12370 (N_12370,N_12121,N_12202);
and U12371 (N_12371,N_12182,N_12253);
or U12372 (N_12372,N_12091,N_12125);
nand U12373 (N_12373,N_12077,N_12157);
and U12374 (N_12374,N_12112,N_12063);
nand U12375 (N_12375,N_12036,N_12185);
xor U12376 (N_12376,N_12028,N_12014);
or U12377 (N_12377,N_12247,N_12104);
nand U12378 (N_12378,N_12158,N_12039);
nor U12379 (N_12379,N_12197,N_12110);
nor U12380 (N_12380,N_12056,N_12159);
xnor U12381 (N_12381,N_12228,N_12106);
xnor U12382 (N_12382,N_12167,N_12095);
nor U12383 (N_12383,N_12074,N_12061);
and U12384 (N_12384,N_12071,N_12191);
xnor U12385 (N_12385,N_12151,N_12089);
and U12386 (N_12386,N_12276,N_12033);
or U12387 (N_12387,N_12053,N_12023);
xor U12388 (N_12388,N_12162,N_12010);
nand U12389 (N_12389,N_12263,N_12252);
and U12390 (N_12390,N_12208,N_12019);
nand U12391 (N_12391,N_12232,N_12080);
nand U12392 (N_12392,N_12108,N_12291);
nor U12393 (N_12393,N_12196,N_12217);
nor U12394 (N_12394,N_12257,N_12011);
or U12395 (N_12395,N_12047,N_12034);
nand U12396 (N_12396,N_12189,N_12082);
or U12397 (N_12397,N_12204,N_12226);
nor U12398 (N_12398,N_12005,N_12043);
and U12399 (N_12399,N_12099,N_12176);
or U12400 (N_12400,N_12254,N_12073);
xor U12401 (N_12401,N_12271,N_12206);
nand U12402 (N_12402,N_12270,N_12075);
xnor U12403 (N_12403,N_12287,N_12026);
xor U12404 (N_12404,N_12154,N_12163);
nor U12405 (N_12405,N_12068,N_12055);
nor U12406 (N_12406,N_12245,N_12268);
nor U12407 (N_12407,N_12272,N_12269);
nand U12408 (N_12408,N_12190,N_12210);
and U12409 (N_12409,N_12144,N_12266);
nand U12410 (N_12410,N_12297,N_12177);
nand U12411 (N_12411,N_12288,N_12172);
nor U12412 (N_12412,N_12237,N_12097);
nand U12413 (N_12413,N_12025,N_12008);
nand U12414 (N_12414,N_12153,N_12042);
nand U12415 (N_12415,N_12003,N_12273);
and U12416 (N_12416,N_12239,N_12140);
and U12417 (N_12417,N_12289,N_12102);
and U12418 (N_12418,N_12050,N_12216);
nand U12419 (N_12419,N_12240,N_12150);
and U12420 (N_12420,N_12069,N_12282);
xnor U12421 (N_12421,N_12049,N_12160);
or U12422 (N_12422,N_12139,N_12205);
nor U12423 (N_12423,N_12015,N_12231);
or U12424 (N_12424,N_12220,N_12201);
nand U12425 (N_12425,N_12129,N_12180);
xnor U12426 (N_12426,N_12203,N_12123);
nand U12427 (N_12427,N_12246,N_12219);
nand U12428 (N_12428,N_12175,N_12155);
and U12429 (N_12429,N_12017,N_12029);
nand U12430 (N_12430,N_12111,N_12242);
nand U12431 (N_12431,N_12200,N_12249);
xnor U12432 (N_12432,N_12193,N_12013);
and U12433 (N_12433,N_12064,N_12098);
nand U12434 (N_12434,N_12030,N_12105);
and U12435 (N_12435,N_12233,N_12171);
nor U12436 (N_12436,N_12146,N_12092);
and U12437 (N_12437,N_12048,N_12290);
nor U12438 (N_12438,N_12116,N_12229);
nor U12439 (N_12439,N_12100,N_12132);
xor U12440 (N_12440,N_12115,N_12083);
or U12441 (N_12441,N_12041,N_12183);
or U12442 (N_12442,N_12000,N_12147);
nor U12443 (N_12443,N_12274,N_12004);
xor U12444 (N_12444,N_12076,N_12094);
nand U12445 (N_12445,N_12021,N_12149);
xnor U12446 (N_12446,N_12188,N_12214);
xnor U12447 (N_12447,N_12065,N_12101);
nand U12448 (N_12448,N_12072,N_12292);
nor U12449 (N_12449,N_12045,N_12215);
nor U12450 (N_12450,N_12092,N_12087);
and U12451 (N_12451,N_12072,N_12196);
or U12452 (N_12452,N_12247,N_12226);
xnor U12453 (N_12453,N_12272,N_12100);
nand U12454 (N_12454,N_12082,N_12076);
or U12455 (N_12455,N_12045,N_12222);
and U12456 (N_12456,N_12229,N_12171);
and U12457 (N_12457,N_12104,N_12122);
nor U12458 (N_12458,N_12200,N_12073);
or U12459 (N_12459,N_12234,N_12246);
and U12460 (N_12460,N_12045,N_12120);
or U12461 (N_12461,N_12045,N_12059);
nor U12462 (N_12462,N_12024,N_12041);
or U12463 (N_12463,N_12240,N_12129);
and U12464 (N_12464,N_12199,N_12209);
and U12465 (N_12465,N_12129,N_12102);
xnor U12466 (N_12466,N_12116,N_12055);
xor U12467 (N_12467,N_12295,N_12111);
nand U12468 (N_12468,N_12159,N_12063);
nand U12469 (N_12469,N_12192,N_12134);
nor U12470 (N_12470,N_12063,N_12069);
xor U12471 (N_12471,N_12077,N_12174);
nor U12472 (N_12472,N_12153,N_12255);
and U12473 (N_12473,N_12020,N_12288);
xnor U12474 (N_12474,N_12110,N_12025);
nand U12475 (N_12475,N_12175,N_12190);
nor U12476 (N_12476,N_12157,N_12264);
or U12477 (N_12477,N_12244,N_12274);
nor U12478 (N_12478,N_12111,N_12148);
nand U12479 (N_12479,N_12124,N_12148);
nor U12480 (N_12480,N_12236,N_12083);
xor U12481 (N_12481,N_12255,N_12107);
or U12482 (N_12482,N_12069,N_12104);
and U12483 (N_12483,N_12175,N_12110);
nand U12484 (N_12484,N_12026,N_12193);
xor U12485 (N_12485,N_12006,N_12247);
nor U12486 (N_12486,N_12240,N_12193);
nor U12487 (N_12487,N_12064,N_12039);
xnor U12488 (N_12488,N_12223,N_12033);
nand U12489 (N_12489,N_12224,N_12079);
or U12490 (N_12490,N_12061,N_12119);
nand U12491 (N_12491,N_12065,N_12114);
nand U12492 (N_12492,N_12017,N_12119);
nand U12493 (N_12493,N_12153,N_12068);
or U12494 (N_12494,N_12071,N_12039);
xnor U12495 (N_12495,N_12092,N_12205);
nand U12496 (N_12496,N_12244,N_12137);
or U12497 (N_12497,N_12028,N_12102);
or U12498 (N_12498,N_12178,N_12219);
or U12499 (N_12499,N_12295,N_12269);
nor U12500 (N_12500,N_12050,N_12173);
xnor U12501 (N_12501,N_12283,N_12260);
nor U12502 (N_12502,N_12234,N_12071);
or U12503 (N_12503,N_12128,N_12097);
and U12504 (N_12504,N_12078,N_12295);
xnor U12505 (N_12505,N_12030,N_12059);
xnor U12506 (N_12506,N_12290,N_12045);
and U12507 (N_12507,N_12289,N_12243);
or U12508 (N_12508,N_12050,N_12070);
nand U12509 (N_12509,N_12274,N_12034);
nor U12510 (N_12510,N_12147,N_12089);
nor U12511 (N_12511,N_12289,N_12119);
or U12512 (N_12512,N_12045,N_12265);
or U12513 (N_12513,N_12133,N_12278);
xnor U12514 (N_12514,N_12170,N_12113);
nand U12515 (N_12515,N_12220,N_12239);
and U12516 (N_12516,N_12254,N_12242);
or U12517 (N_12517,N_12100,N_12169);
or U12518 (N_12518,N_12115,N_12178);
or U12519 (N_12519,N_12121,N_12165);
xor U12520 (N_12520,N_12165,N_12021);
and U12521 (N_12521,N_12219,N_12001);
and U12522 (N_12522,N_12061,N_12101);
xnor U12523 (N_12523,N_12253,N_12296);
xor U12524 (N_12524,N_12074,N_12293);
nor U12525 (N_12525,N_12089,N_12234);
nor U12526 (N_12526,N_12141,N_12072);
nand U12527 (N_12527,N_12261,N_12125);
xor U12528 (N_12528,N_12023,N_12055);
nor U12529 (N_12529,N_12090,N_12162);
nor U12530 (N_12530,N_12139,N_12095);
xor U12531 (N_12531,N_12283,N_12014);
and U12532 (N_12532,N_12200,N_12287);
xnor U12533 (N_12533,N_12222,N_12030);
nand U12534 (N_12534,N_12182,N_12071);
nor U12535 (N_12535,N_12089,N_12241);
and U12536 (N_12536,N_12285,N_12102);
xor U12537 (N_12537,N_12115,N_12048);
and U12538 (N_12538,N_12179,N_12216);
nand U12539 (N_12539,N_12247,N_12071);
nor U12540 (N_12540,N_12007,N_12045);
or U12541 (N_12541,N_12045,N_12028);
nand U12542 (N_12542,N_12168,N_12297);
and U12543 (N_12543,N_12214,N_12179);
or U12544 (N_12544,N_12153,N_12291);
xor U12545 (N_12545,N_12196,N_12250);
nor U12546 (N_12546,N_12043,N_12213);
nor U12547 (N_12547,N_12191,N_12284);
nand U12548 (N_12548,N_12011,N_12151);
or U12549 (N_12549,N_12229,N_12246);
and U12550 (N_12550,N_12251,N_12155);
xnor U12551 (N_12551,N_12106,N_12191);
or U12552 (N_12552,N_12032,N_12086);
xor U12553 (N_12553,N_12102,N_12107);
nand U12554 (N_12554,N_12261,N_12293);
and U12555 (N_12555,N_12098,N_12203);
nor U12556 (N_12556,N_12035,N_12085);
xnor U12557 (N_12557,N_12126,N_12127);
nor U12558 (N_12558,N_12267,N_12298);
or U12559 (N_12559,N_12180,N_12246);
and U12560 (N_12560,N_12253,N_12085);
or U12561 (N_12561,N_12051,N_12151);
xnor U12562 (N_12562,N_12275,N_12205);
or U12563 (N_12563,N_12197,N_12255);
and U12564 (N_12564,N_12146,N_12132);
nand U12565 (N_12565,N_12139,N_12284);
nor U12566 (N_12566,N_12147,N_12183);
nor U12567 (N_12567,N_12131,N_12166);
xnor U12568 (N_12568,N_12045,N_12114);
or U12569 (N_12569,N_12248,N_12201);
and U12570 (N_12570,N_12005,N_12011);
nor U12571 (N_12571,N_12262,N_12205);
and U12572 (N_12572,N_12187,N_12273);
and U12573 (N_12573,N_12225,N_12193);
and U12574 (N_12574,N_12236,N_12299);
nor U12575 (N_12575,N_12115,N_12103);
or U12576 (N_12576,N_12200,N_12018);
and U12577 (N_12577,N_12060,N_12208);
nand U12578 (N_12578,N_12170,N_12295);
nand U12579 (N_12579,N_12205,N_12194);
nor U12580 (N_12580,N_12169,N_12025);
or U12581 (N_12581,N_12191,N_12017);
or U12582 (N_12582,N_12117,N_12294);
nor U12583 (N_12583,N_12031,N_12287);
nand U12584 (N_12584,N_12081,N_12108);
and U12585 (N_12585,N_12266,N_12038);
xor U12586 (N_12586,N_12133,N_12010);
or U12587 (N_12587,N_12011,N_12249);
nor U12588 (N_12588,N_12109,N_12075);
or U12589 (N_12589,N_12232,N_12120);
and U12590 (N_12590,N_12190,N_12151);
or U12591 (N_12591,N_12169,N_12098);
or U12592 (N_12592,N_12222,N_12253);
and U12593 (N_12593,N_12056,N_12242);
or U12594 (N_12594,N_12061,N_12207);
and U12595 (N_12595,N_12134,N_12286);
or U12596 (N_12596,N_12279,N_12269);
or U12597 (N_12597,N_12149,N_12011);
and U12598 (N_12598,N_12213,N_12169);
xor U12599 (N_12599,N_12138,N_12176);
nor U12600 (N_12600,N_12333,N_12405);
xnor U12601 (N_12601,N_12481,N_12519);
nor U12602 (N_12602,N_12570,N_12585);
or U12603 (N_12603,N_12401,N_12336);
nor U12604 (N_12604,N_12461,N_12334);
nand U12605 (N_12605,N_12531,N_12545);
xor U12606 (N_12606,N_12501,N_12568);
nor U12607 (N_12607,N_12534,N_12451);
nor U12608 (N_12608,N_12548,N_12458);
nor U12609 (N_12609,N_12495,N_12587);
nand U12610 (N_12610,N_12374,N_12423);
nand U12611 (N_12611,N_12470,N_12376);
or U12612 (N_12612,N_12300,N_12506);
xor U12613 (N_12613,N_12472,N_12464);
nand U12614 (N_12614,N_12566,N_12349);
or U12615 (N_12615,N_12473,N_12590);
nor U12616 (N_12616,N_12364,N_12434);
nor U12617 (N_12617,N_12459,N_12468);
or U12618 (N_12618,N_12354,N_12476);
nand U12619 (N_12619,N_12457,N_12445);
nor U12620 (N_12620,N_12450,N_12523);
and U12621 (N_12621,N_12555,N_12517);
nor U12622 (N_12622,N_12493,N_12303);
nand U12623 (N_12623,N_12508,N_12504);
or U12624 (N_12624,N_12496,N_12500);
or U12625 (N_12625,N_12417,N_12340);
nand U12626 (N_12626,N_12379,N_12331);
nand U12627 (N_12627,N_12572,N_12395);
or U12628 (N_12628,N_12484,N_12592);
nand U12629 (N_12629,N_12426,N_12528);
or U12630 (N_12630,N_12318,N_12507);
nor U12631 (N_12631,N_12540,N_12490);
nor U12632 (N_12632,N_12368,N_12521);
nand U12633 (N_12633,N_12448,N_12332);
and U12634 (N_12634,N_12360,N_12560);
xor U12635 (N_12635,N_12538,N_12554);
or U12636 (N_12636,N_12411,N_12339);
and U12637 (N_12637,N_12418,N_12357);
xor U12638 (N_12638,N_12378,N_12479);
xnor U12639 (N_12639,N_12584,N_12355);
xor U12640 (N_12640,N_12591,N_12322);
nor U12641 (N_12641,N_12467,N_12558);
or U12642 (N_12642,N_12463,N_12577);
nand U12643 (N_12643,N_12342,N_12377);
nand U12644 (N_12644,N_12466,N_12365);
nand U12645 (N_12645,N_12406,N_12326);
nand U12646 (N_12646,N_12361,N_12443);
or U12647 (N_12647,N_12565,N_12546);
nor U12648 (N_12648,N_12543,N_12449);
nand U12649 (N_12649,N_12578,N_12439);
and U12650 (N_12650,N_12593,N_12444);
or U12651 (N_12651,N_12414,N_12441);
and U12652 (N_12652,N_12310,N_12579);
and U12653 (N_12653,N_12351,N_12323);
nor U12654 (N_12654,N_12487,N_12460);
nand U12655 (N_12655,N_12419,N_12350);
xor U12656 (N_12656,N_12338,N_12583);
and U12657 (N_12657,N_12478,N_12574);
and U12658 (N_12658,N_12305,N_12391);
and U12659 (N_12659,N_12345,N_12569);
nand U12660 (N_12660,N_12327,N_12509);
nor U12661 (N_12661,N_12527,N_12375);
nand U12662 (N_12662,N_12409,N_12367);
or U12663 (N_12663,N_12399,N_12510);
nand U12664 (N_12664,N_12525,N_12488);
or U12665 (N_12665,N_12413,N_12304);
or U12666 (N_12666,N_12471,N_12561);
and U12667 (N_12667,N_12393,N_12422);
nand U12668 (N_12668,N_12522,N_12486);
xor U12669 (N_12669,N_12415,N_12370);
and U12670 (N_12670,N_12311,N_12314);
nand U12671 (N_12671,N_12524,N_12316);
xor U12672 (N_12672,N_12550,N_12547);
or U12673 (N_12673,N_12429,N_12541);
or U12674 (N_12674,N_12556,N_12384);
nand U12675 (N_12675,N_12456,N_12567);
nor U12676 (N_12676,N_12420,N_12313);
xnor U12677 (N_12677,N_12480,N_12483);
nand U12678 (N_12678,N_12412,N_12553);
nor U12679 (N_12679,N_12588,N_12343);
nor U12680 (N_12680,N_12482,N_12372);
xnor U12681 (N_12681,N_12398,N_12402);
nor U12682 (N_12682,N_12475,N_12396);
or U12683 (N_12683,N_12551,N_12386);
and U12684 (N_12684,N_12505,N_12542);
xnor U12685 (N_12685,N_12388,N_12576);
and U12686 (N_12686,N_12453,N_12537);
xnor U12687 (N_12687,N_12430,N_12529);
xor U12688 (N_12688,N_12492,N_12328);
xnor U12689 (N_12689,N_12474,N_12369);
xnor U12690 (N_12690,N_12516,N_12597);
nand U12691 (N_12691,N_12366,N_12544);
nand U12692 (N_12692,N_12321,N_12563);
xor U12693 (N_12693,N_12526,N_12301);
xnor U12694 (N_12694,N_12494,N_12440);
nor U12695 (N_12695,N_12389,N_12515);
nor U12696 (N_12696,N_12358,N_12337);
and U12697 (N_12697,N_12373,N_12595);
or U12698 (N_12698,N_12432,N_12329);
or U12699 (N_12699,N_12416,N_12433);
xnor U12700 (N_12700,N_12520,N_12539);
xnor U12701 (N_12701,N_12320,N_12477);
and U12702 (N_12702,N_12346,N_12573);
or U12703 (N_12703,N_12557,N_12594);
and U12704 (N_12704,N_12586,N_12307);
nand U12705 (N_12705,N_12497,N_12403);
or U12706 (N_12706,N_12552,N_12302);
and U12707 (N_12707,N_12599,N_12530);
nor U12708 (N_12708,N_12518,N_12344);
or U12709 (N_12709,N_12598,N_12353);
or U12710 (N_12710,N_12455,N_12571);
nor U12711 (N_12711,N_12380,N_12424);
nand U12712 (N_12712,N_12356,N_12581);
xnor U12713 (N_12713,N_12341,N_12462);
xnor U12714 (N_12714,N_12410,N_12408);
xor U12715 (N_12715,N_12363,N_12397);
and U12716 (N_12716,N_12315,N_12549);
nand U12717 (N_12717,N_12446,N_12306);
nor U12718 (N_12718,N_12511,N_12431);
or U12719 (N_12719,N_12512,N_12394);
nor U12720 (N_12720,N_12447,N_12324);
nand U12721 (N_12721,N_12404,N_12335);
xnor U12722 (N_12722,N_12442,N_12390);
xor U12723 (N_12723,N_12308,N_12359);
xor U12724 (N_12724,N_12564,N_12381);
or U12725 (N_12725,N_12428,N_12427);
xor U12726 (N_12726,N_12491,N_12536);
xor U12727 (N_12727,N_12352,N_12371);
xnor U12728 (N_12728,N_12348,N_12407);
xor U12729 (N_12729,N_12347,N_12382);
nor U12730 (N_12730,N_12514,N_12503);
nand U12731 (N_12731,N_12452,N_12383);
nor U12732 (N_12732,N_12400,N_12465);
or U12733 (N_12733,N_12454,N_12580);
or U12734 (N_12734,N_12330,N_12309);
nand U12735 (N_12735,N_12319,N_12596);
xor U12736 (N_12736,N_12532,N_12387);
xor U12737 (N_12737,N_12362,N_12421);
and U12738 (N_12738,N_12438,N_12469);
and U12739 (N_12739,N_12589,N_12559);
nand U12740 (N_12740,N_12425,N_12498);
or U12741 (N_12741,N_12513,N_12325);
and U12742 (N_12742,N_12499,N_12575);
or U12743 (N_12743,N_12437,N_12392);
nand U12744 (N_12744,N_12485,N_12385);
nor U12745 (N_12745,N_12317,N_12312);
nor U12746 (N_12746,N_12436,N_12502);
nor U12747 (N_12747,N_12562,N_12582);
xor U12748 (N_12748,N_12489,N_12535);
xor U12749 (N_12749,N_12435,N_12533);
nor U12750 (N_12750,N_12454,N_12551);
or U12751 (N_12751,N_12525,N_12435);
nand U12752 (N_12752,N_12349,N_12402);
nand U12753 (N_12753,N_12418,N_12501);
and U12754 (N_12754,N_12442,N_12515);
or U12755 (N_12755,N_12483,N_12563);
nor U12756 (N_12756,N_12377,N_12379);
or U12757 (N_12757,N_12352,N_12396);
nor U12758 (N_12758,N_12368,N_12450);
and U12759 (N_12759,N_12470,N_12367);
xnor U12760 (N_12760,N_12313,N_12599);
nand U12761 (N_12761,N_12353,N_12374);
and U12762 (N_12762,N_12342,N_12369);
nor U12763 (N_12763,N_12595,N_12407);
and U12764 (N_12764,N_12429,N_12425);
nor U12765 (N_12765,N_12412,N_12531);
nand U12766 (N_12766,N_12544,N_12384);
and U12767 (N_12767,N_12395,N_12472);
and U12768 (N_12768,N_12348,N_12301);
nor U12769 (N_12769,N_12454,N_12360);
xnor U12770 (N_12770,N_12416,N_12518);
or U12771 (N_12771,N_12336,N_12391);
nor U12772 (N_12772,N_12411,N_12343);
and U12773 (N_12773,N_12578,N_12482);
nor U12774 (N_12774,N_12471,N_12542);
nor U12775 (N_12775,N_12454,N_12337);
or U12776 (N_12776,N_12571,N_12376);
xor U12777 (N_12777,N_12416,N_12389);
or U12778 (N_12778,N_12520,N_12371);
nor U12779 (N_12779,N_12480,N_12558);
nand U12780 (N_12780,N_12534,N_12572);
and U12781 (N_12781,N_12371,N_12529);
or U12782 (N_12782,N_12447,N_12405);
nand U12783 (N_12783,N_12567,N_12479);
xor U12784 (N_12784,N_12517,N_12591);
nor U12785 (N_12785,N_12326,N_12385);
xor U12786 (N_12786,N_12556,N_12359);
and U12787 (N_12787,N_12327,N_12313);
xnor U12788 (N_12788,N_12396,N_12305);
nor U12789 (N_12789,N_12395,N_12328);
and U12790 (N_12790,N_12598,N_12323);
or U12791 (N_12791,N_12564,N_12419);
nand U12792 (N_12792,N_12347,N_12421);
or U12793 (N_12793,N_12425,N_12339);
xnor U12794 (N_12794,N_12592,N_12513);
nand U12795 (N_12795,N_12548,N_12487);
or U12796 (N_12796,N_12470,N_12441);
or U12797 (N_12797,N_12434,N_12468);
and U12798 (N_12798,N_12534,N_12569);
nor U12799 (N_12799,N_12311,N_12446);
nor U12800 (N_12800,N_12457,N_12549);
xnor U12801 (N_12801,N_12541,N_12538);
nor U12802 (N_12802,N_12326,N_12407);
or U12803 (N_12803,N_12402,N_12568);
nand U12804 (N_12804,N_12424,N_12389);
and U12805 (N_12805,N_12313,N_12382);
or U12806 (N_12806,N_12441,N_12462);
and U12807 (N_12807,N_12493,N_12486);
nand U12808 (N_12808,N_12406,N_12592);
and U12809 (N_12809,N_12349,N_12448);
nand U12810 (N_12810,N_12584,N_12411);
nor U12811 (N_12811,N_12478,N_12502);
nor U12812 (N_12812,N_12505,N_12495);
and U12813 (N_12813,N_12340,N_12549);
nor U12814 (N_12814,N_12362,N_12523);
nand U12815 (N_12815,N_12433,N_12536);
nor U12816 (N_12816,N_12586,N_12580);
and U12817 (N_12817,N_12441,N_12468);
and U12818 (N_12818,N_12327,N_12444);
and U12819 (N_12819,N_12467,N_12324);
or U12820 (N_12820,N_12327,N_12452);
and U12821 (N_12821,N_12345,N_12484);
and U12822 (N_12822,N_12584,N_12489);
or U12823 (N_12823,N_12428,N_12368);
nor U12824 (N_12824,N_12379,N_12367);
nand U12825 (N_12825,N_12359,N_12453);
nor U12826 (N_12826,N_12329,N_12488);
nor U12827 (N_12827,N_12499,N_12321);
xnor U12828 (N_12828,N_12479,N_12322);
nand U12829 (N_12829,N_12304,N_12428);
nor U12830 (N_12830,N_12351,N_12516);
and U12831 (N_12831,N_12474,N_12450);
nor U12832 (N_12832,N_12562,N_12312);
or U12833 (N_12833,N_12589,N_12433);
nor U12834 (N_12834,N_12361,N_12593);
or U12835 (N_12835,N_12502,N_12490);
nor U12836 (N_12836,N_12395,N_12342);
nand U12837 (N_12837,N_12462,N_12560);
and U12838 (N_12838,N_12303,N_12441);
xor U12839 (N_12839,N_12300,N_12424);
and U12840 (N_12840,N_12517,N_12478);
nand U12841 (N_12841,N_12513,N_12457);
xnor U12842 (N_12842,N_12493,N_12401);
and U12843 (N_12843,N_12587,N_12553);
and U12844 (N_12844,N_12595,N_12452);
nand U12845 (N_12845,N_12340,N_12320);
xnor U12846 (N_12846,N_12453,N_12307);
or U12847 (N_12847,N_12469,N_12332);
or U12848 (N_12848,N_12569,N_12320);
nor U12849 (N_12849,N_12550,N_12444);
and U12850 (N_12850,N_12437,N_12425);
and U12851 (N_12851,N_12331,N_12567);
xor U12852 (N_12852,N_12509,N_12454);
nand U12853 (N_12853,N_12470,N_12339);
nor U12854 (N_12854,N_12392,N_12407);
nor U12855 (N_12855,N_12544,N_12383);
xnor U12856 (N_12856,N_12535,N_12553);
nor U12857 (N_12857,N_12396,N_12409);
nand U12858 (N_12858,N_12394,N_12459);
xor U12859 (N_12859,N_12501,N_12433);
or U12860 (N_12860,N_12301,N_12550);
and U12861 (N_12861,N_12576,N_12488);
nor U12862 (N_12862,N_12333,N_12440);
and U12863 (N_12863,N_12322,N_12482);
xnor U12864 (N_12864,N_12583,N_12438);
nor U12865 (N_12865,N_12364,N_12542);
or U12866 (N_12866,N_12517,N_12563);
xnor U12867 (N_12867,N_12322,N_12390);
nand U12868 (N_12868,N_12304,N_12484);
xnor U12869 (N_12869,N_12412,N_12330);
nor U12870 (N_12870,N_12499,N_12473);
or U12871 (N_12871,N_12547,N_12527);
nor U12872 (N_12872,N_12359,N_12575);
or U12873 (N_12873,N_12485,N_12588);
and U12874 (N_12874,N_12385,N_12512);
nor U12875 (N_12875,N_12356,N_12348);
nor U12876 (N_12876,N_12370,N_12424);
nor U12877 (N_12877,N_12584,N_12312);
xor U12878 (N_12878,N_12551,N_12522);
nand U12879 (N_12879,N_12314,N_12591);
xnor U12880 (N_12880,N_12469,N_12365);
xor U12881 (N_12881,N_12400,N_12349);
or U12882 (N_12882,N_12549,N_12310);
nand U12883 (N_12883,N_12466,N_12454);
nand U12884 (N_12884,N_12321,N_12598);
and U12885 (N_12885,N_12440,N_12589);
xnor U12886 (N_12886,N_12402,N_12491);
nand U12887 (N_12887,N_12302,N_12424);
xnor U12888 (N_12888,N_12429,N_12340);
nor U12889 (N_12889,N_12353,N_12551);
or U12890 (N_12890,N_12357,N_12316);
nor U12891 (N_12891,N_12373,N_12313);
nand U12892 (N_12892,N_12373,N_12376);
nand U12893 (N_12893,N_12456,N_12506);
nor U12894 (N_12894,N_12440,N_12523);
nand U12895 (N_12895,N_12362,N_12376);
and U12896 (N_12896,N_12526,N_12335);
nand U12897 (N_12897,N_12449,N_12444);
nand U12898 (N_12898,N_12589,N_12317);
nor U12899 (N_12899,N_12510,N_12564);
nand U12900 (N_12900,N_12898,N_12840);
nand U12901 (N_12901,N_12658,N_12750);
xor U12902 (N_12902,N_12769,N_12804);
nor U12903 (N_12903,N_12762,N_12678);
and U12904 (N_12904,N_12827,N_12697);
nor U12905 (N_12905,N_12615,N_12691);
xor U12906 (N_12906,N_12708,N_12745);
nand U12907 (N_12907,N_12893,N_12705);
or U12908 (N_12908,N_12810,N_12754);
nor U12909 (N_12909,N_12880,N_12715);
nor U12910 (N_12910,N_12735,N_12857);
and U12911 (N_12911,N_12757,N_12849);
or U12912 (N_12912,N_12878,N_12694);
and U12913 (N_12913,N_12764,N_12797);
nor U12914 (N_12914,N_12700,N_12648);
and U12915 (N_12915,N_12679,N_12874);
xnor U12916 (N_12916,N_12741,N_12733);
nand U12917 (N_12917,N_12875,N_12825);
xnor U12918 (N_12918,N_12627,N_12839);
xor U12919 (N_12919,N_12714,N_12855);
or U12920 (N_12920,N_12752,N_12672);
nor U12921 (N_12921,N_12766,N_12685);
nand U12922 (N_12922,N_12725,N_12604);
nand U12923 (N_12923,N_12780,N_12701);
and U12924 (N_12924,N_12767,N_12748);
or U12925 (N_12925,N_12660,N_12768);
or U12926 (N_12926,N_12634,N_12652);
and U12927 (N_12927,N_12605,N_12883);
xnor U12928 (N_12928,N_12713,N_12772);
nor U12929 (N_12929,N_12644,N_12729);
or U12930 (N_12930,N_12837,N_12747);
nor U12931 (N_12931,N_12899,N_12770);
xnor U12932 (N_12932,N_12881,N_12868);
and U12933 (N_12933,N_12819,N_12765);
or U12934 (N_12934,N_12856,N_12812);
xor U12935 (N_12935,N_12854,N_12873);
xor U12936 (N_12936,N_12816,N_12844);
nand U12937 (N_12937,N_12782,N_12633);
or U12938 (N_12938,N_12800,N_12756);
or U12939 (N_12939,N_12609,N_12630);
nor U12940 (N_12940,N_12793,N_12641);
nor U12941 (N_12941,N_12711,N_12621);
nor U12942 (N_12942,N_12867,N_12744);
xnor U12943 (N_12943,N_12699,N_12818);
and U12944 (N_12944,N_12631,N_12677);
nor U12945 (N_12945,N_12753,N_12689);
xnor U12946 (N_12946,N_12673,N_12608);
and U12947 (N_12947,N_12692,N_12783);
xnor U12948 (N_12948,N_12826,N_12852);
and U12949 (N_12949,N_12718,N_12645);
xnor U12950 (N_12950,N_12730,N_12661);
or U12951 (N_12951,N_12734,N_12789);
nand U12952 (N_12952,N_12629,N_12619);
nor U12953 (N_12953,N_12610,N_12802);
and U12954 (N_12954,N_12879,N_12895);
and U12955 (N_12955,N_12832,N_12728);
and U12956 (N_12956,N_12727,N_12788);
and U12957 (N_12957,N_12654,N_12666);
nand U12958 (N_12958,N_12693,N_12636);
or U12959 (N_12959,N_12784,N_12801);
nor U12960 (N_12960,N_12822,N_12876);
or U12961 (N_12961,N_12862,N_12670);
xnor U12962 (N_12962,N_12732,N_12817);
or U12963 (N_12963,N_12760,N_12842);
or U12964 (N_12964,N_12871,N_12829);
and U12965 (N_12965,N_12647,N_12758);
nand U12966 (N_12966,N_12888,N_12830);
nand U12967 (N_12967,N_12726,N_12649);
or U12968 (N_12968,N_12882,N_12743);
and U12969 (N_12969,N_12651,N_12877);
nand U12970 (N_12970,N_12795,N_12796);
xor U12971 (N_12971,N_12720,N_12785);
xnor U12972 (N_12972,N_12624,N_12847);
nand U12973 (N_12973,N_12731,N_12657);
or U12974 (N_12974,N_12653,N_12859);
nor U12975 (N_12975,N_12755,N_12884);
nand U12976 (N_12976,N_12845,N_12751);
nor U12977 (N_12977,N_12669,N_12712);
and U12978 (N_12978,N_12626,N_12864);
nor U12979 (N_12979,N_12646,N_12665);
nand U12980 (N_12980,N_12863,N_12777);
nor U12981 (N_12981,N_12828,N_12775);
xnor U12982 (N_12982,N_12815,N_12707);
or U12983 (N_12983,N_12637,N_12602);
nand U12984 (N_12984,N_12771,N_12601);
and U12985 (N_12985,N_12723,N_12890);
xnor U12986 (N_12986,N_12836,N_12886);
or U12987 (N_12987,N_12616,N_12695);
xor U12988 (N_12988,N_12639,N_12740);
nor U12989 (N_12989,N_12719,N_12716);
or U12990 (N_12990,N_12749,N_12709);
or U12991 (N_12991,N_12831,N_12787);
nor U12992 (N_12992,N_12702,N_12663);
and U12993 (N_12993,N_12617,N_12683);
nand U12994 (N_12994,N_12865,N_12682);
xor U12995 (N_12995,N_12778,N_12835);
xor U12996 (N_12996,N_12806,N_12791);
xor U12997 (N_12997,N_12834,N_12662);
and U12998 (N_12998,N_12671,N_12612);
nand U12999 (N_12999,N_12710,N_12640);
and U13000 (N_13000,N_12659,N_12870);
nor U13001 (N_13001,N_12623,N_12687);
nand U13002 (N_13002,N_12613,N_12736);
nor U13003 (N_13003,N_12739,N_12724);
nor U13004 (N_13004,N_12622,N_12696);
nor U13005 (N_13005,N_12869,N_12684);
xnor U13006 (N_13006,N_12607,N_12706);
nand U13007 (N_13007,N_12650,N_12896);
or U13008 (N_13008,N_12704,N_12635);
nor U13009 (N_13009,N_12858,N_12737);
xnor U13010 (N_13010,N_12638,N_12794);
or U13011 (N_13011,N_12798,N_12843);
nand U13012 (N_13012,N_12688,N_12675);
nor U13013 (N_13013,N_12820,N_12811);
and U13014 (N_13014,N_12807,N_12738);
xnor U13015 (N_13015,N_12632,N_12763);
nor U13016 (N_13016,N_12600,N_12773);
or U13017 (N_13017,N_12759,N_12643);
and U13018 (N_13018,N_12676,N_12860);
xnor U13019 (N_13019,N_12667,N_12866);
nand U13020 (N_13020,N_12897,N_12603);
xor U13021 (N_13021,N_12790,N_12885);
and U13022 (N_13022,N_12838,N_12618);
nand U13023 (N_13023,N_12681,N_12680);
and U13024 (N_13024,N_12887,N_12803);
nor U13025 (N_13025,N_12889,N_12722);
and U13026 (N_13026,N_12774,N_12853);
or U13027 (N_13027,N_12846,N_12655);
and U13028 (N_13028,N_12668,N_12628);
and U13029 (N_13029,N_12781,N_12642);
and U13030 (N_13030,N_12742,N_12779);
xnor U13031 (N_13031,N_12786,N_12656);
nor U13032 (N_13032,N_12674,N_12703);
and U13033 (N_13033,N_12761,N_12792);
nor U13034 (N_13034,N_12841,N_12809);
xnor U13035 (N_13035,N_12698,N_12833);
or U13036 (N_13036,N_12872,N_12620);
nand U13037 (N_13037,N_12606,N_12894);
nand U13038 (N_13038,N_12799,N_12861);
nor U13039 (N_13039,N_12813,N_12821);
and U13040 (N_13040,N_12611,N_12805);
xor U13041 (N_13041,N_12848,N_12823);
nand U13042 (N_13042,N_12808,N_12850);
xor U13043 (N_13043,N_12686,N_12625);
nor U13044 (N_13044,N_12824,N_12614);
and U13045 (N_13045,N_12776,N_12717);
xnor U13046 (N_13046,N_12664,N_12690);
and U13047 (N_13047,N_12721,N_12746);
or U13048 (N_13048,N_12814,N_12892);
and U13049 (N_13049,N_12851,N_12891);
xnor U13050 (N_13050,N_12660,N_12822);
and U13051 (N_13051,N_12880,N_12796);
nor U13052 (N_13052,N_12657,N_12711);
and U13053 (N_13053,N_12872,N_12678);
xor U13054 (N_13054,N_12806,N_12764);
nor U13055 (N_13055,N_12846,N_12706);
xnor U13056 (N_13056,N_12779,N_12606);
nand U13057 (N_13057,N_12624,N_12809);
xnor U13058 (N_13058,N_12624,N_12652);
nor U13059 (N_13059,N_12604,N_12636);
or U13060 (N_13060,N_12683,N_12885);
nor U13061 (N_13061,N_12696,N_12766);
nand U13062 (N_13062,N_12746,N_12645);
nor U13063 (N_13063,N_12751,N_12768);
xor U13064 (N_13064,N_12651,N_12708);
or U13065 (N_13065,N_12767,N_12632);
nand U13066 (N_13066,N_12815,N_12613);
or U13067 (N_13067,N_12773,N_12770);
nand U13068 (N_13068,N_12619,N_12756);
nand U13069 (N_13069,N_12611,N_12887);
xor U13070 (N_13070,N_12897,N_12844);
and U13071 (N_13071,N_12895,N_12626);
and U13072 (N_13072,N_12748,N_12803);
xnor U13073 (N_13073,N_12675,N_12891);
xnor U13074 (N_13074,N_12603,N_12614);
nand U13075 (N_13075,N_12719,N_12739);
nand U13076 (N_13076,N_12732,N_12844);
xnor U13077 (N_13077,N_12802,N_12637);
or U13078 (N_13078,N_12779,N_12845);
nand U13079 (N_13079,N_12780,N_12777);
or U13080 (N_13080,N_12637,N_12713);
or U13081 (N_13081,N_12832,N_12786);
nor U13082 (N_13082,N_12795,N_12830);
and U13083 (N_13083,N_12660,N_12669);
nand U13084 (N_13084,N_12868,N_12737);
and U13085 (N_13085,N_12623,N_12644);
xnor U13086 (N_13086,N_12798,N_12600);
nand U13087 (N_13087,N_12747,N_12702);
and U13088 (N_13088,N_12773,N_12624);
nand U13089 (N_13089,N_12678,N_12836);
xor U13090 (N_13090,N_12864,N_12781);
nor U13091 (N_13091,N_12777,N_12773);
nand U13092 (N_13092,N_12763,N_12617);
xor U13093 (N_13093,N_12689,N_12815);
xnor U13094 (N_13094,N_12804,N_12646);
and U13095 (N_13095,N_12732,N_12806);
nand U13096 (N_13096,N_12703,N_12769);
or U13097 (N_13097,N_12869,N_12602);
or U13098 (N_13098,N_12820,N_12652);
nand U13099 (N_13099,N_12846,N_12638);
xor U13100 (N_13100,N_12603,N_12767);
and U13101 (N_13101,N_12665,N_12781);
nand U13102 (N_13102,N_12705,N_12702);
xor U13103 (N_13103,N_12814,N_12890);
nand U13104 (N_13104,N_12614,N_12822);
or U13105 (N_13105,N_12849,N_12851);
and U13106 (N_13106,N_12706,N_12684);
and U13107 (N_13107,N_12683,N_12825);
nor U13108 (N_13108,N_12639,N_12791);
or U13109 (N_13109,N_12823,N_12815);
nand U13110 (N_13110,N_12637,N_12625);
and U13111 (N_13111,N_12761,N_12879);
or U13112 (N_13112,N_12763,N_12688);
nand U13113 (N_13113,N_12638,N_12772);
or U13114 (N_13114,N_12692,N_12689);
xor U13115 (N_13115,N_12622,N_12806);
and U13116 (N_13116,N_12884,N_12711);
or U13117 (N_13117,N_12870,N_12723);
or U13118 (N_13118,N_12670,N_12848);
nand U13119 (N_13119,N_12802,N_12765);
and U13120 (N_13120,N_12630,N_12671);
and U13121 (N_13121,N_12796,N_12789);
xor U13122 (N_13122,N_12869,N_12682);
nor U13123 (N_13123,N_12691,N_12805);
nand U13124 (N_13124,N_12814,N_12758);
or U13125 (N_13125,N_12729,N_12803);
nand U13126 (N_13126,N_12668,N_12759);
nor U13127 (N_13127,N_12773,N_12848);
nand U13128 (N_13128,N_12741,N_12866);
and U13129 (N_13129,N_12648,N_12897);
xor U13130 (N_13130,N_12712,N_12888);
nand U13131 (N_13131,N_12850,N_12613);
and U13132 (N_13132,N_12796,N_12810);
nand U13133 (N_13133,N_12874,N_12858);
nor U13134 (N_13134,N_12893,N_12697);
xor U13135 (N_13135,N_12859,N_12895);
nor U13136 (N_13136,N_12752,N_12611);
nor U13137 (N_13137,N_12758,N_12770);
and U13138 (N_13138,N_12762,N_12620);
nand U13139 (N_13139,N_12614,N_12694);
nand U13140 (N_13140,N_12800,N_12629);
nand U13141 (N_13141,N_12631,N_12791);
xnor U13142 (N_13142,N_12830,N_12878);
xor U13143 (N_13143,N_12611,N_12608);
xnor U13144 (N_13144,N_12693,N_12635);
nor U13145 (N_13145,N_12623,N_12750);
or U13146 (N_13146,N_12602,N_12614);
nand U13147 (N_13147,N_12717,N_12811);
nand U13148 (N_13148,N_12643,N_12750);
nor U13149 (N_13149,N_12799,N_12621);
and U13150 (N_13150,N_12833,N_12808);
nor U13151 (N_13151,N_12698,N_12672);
nor U13152 (N_13152,N_12685,N_12645);
nor U13153 (N_13153,N_12857,N_12788);
xnor U13154 (N_13154,N_12885,N_12762);
xor U13155 (N_13155,N_12611,N_12769);
or U13156 (N_13156,N_12848,N_12805);
xor U13157 (N_13157,N_12776,N_12606);
xor U13158 (N_13158,N_12753,N_12803);
nand U13159 (N_13159,N_12788,N_12634);
nor U13160 (N_13160,N_12777,N_12747);
or U13161 (N_13161,N_12659,N_12738);
xnor U13162 (N_13162,N_12833,N_12705);
xor U13163 (N_13163,N_12772,N_12891);
or U13164 (N_13164,N_12698,N_12868);
nand U13165 (N_13165,N_12787,N_12799);
nand U13166 (N_13166,N_12691,N_12760);
xnor U13167 (N_13167,N_12694,N_12732);
or U13168 (N_13168,N_12691,N_12723);
xnor U13169 (N_13169,N_12628,N_12800);
and U13170 (N_13170,N_12881,N_12600);
nor U13171 (N_13171,N_12854,N_12628);
and U13172 (N_13172,N_12793,N_12763);
or U13173 (N_13173,N_12635,N_12699);
or U13174 (N_13174,N_12814,N_12749);
or U13175 (N_13175,N_12716,N_12745);
nor U13176 (N_13176,N_12651,N_12797);
nand U13177 (N_13177,N_12648,N_12804);
xnor U13178 (N_13178,N_12820,N_12701);
nand U13179 (N_13179,N_12775,N_12809);
and U13180 (N_13180,N_12886,N_12622);
and U13181 (N_13181,N_12724,N_12882);
or U13182 (N_13182,N_12770,N_12713);
nand U13183 (N_13183,N_12895,N_12737);
and U13184 (N_13184,N_12843,N_12738);
or U13185 (N_13185,N_12713,N_12714);
nor U13186 (N_13186,N_12662,N_12620);
or U13187 (N_13187,N_12723,N_12690);
and U13188 (N_13188,N_12675,N_12819);
xor U13189 (N_13189,N_12724,N_12768);
or U13190 (N_13190,N_12651,N_12712);
nand U13191 (N_13191,N_12613,N_12643);
or U13192 (N_13192,N_12700,N_12857);
nand U13193 (N_13193,N_12805,N_12724);
nand U13194 (N_13194,N_12790,N_12700);
or U13195 (N_13195,N_12756,N_12846);
nand U13196 (N_13196,N_12724,N_12659);
nand U13197 (N_13197,N_12719,N_12798);
xor U13198 (N_13198,N_12751,N_12850);
nand U13199 (N_13199,N_12781,N_12816);
nand U13200 (N_13200,N_12930,N_12931);
xor U13201 (N_13201,N_13103,N_13143);
nand U13202 (N_13202,N_13183,N_13040);
and U13203 (N_13203,N_12991,N_13177);
nand U13204 (N_13204,N_13084,N_12921);
and U13205 (N_13205,N_12985,N_12975);
nand U13206 (N_13206,N_13115,N_13157);
xor U13207 (N_13207,N_13184,N_13146);
xor U13208 (N_13208,N_13179,N_12924);
and U13209 (N_13209,N_13130,N_12958);
xnor U13210 (N_13210,N_13189,N_13155);
and U13211 (N_13211,N_13015,N_13149);
nor U13212 (N_13212,N_13049,N_13065);
xor U13213 (N_13213,N_13132,N_13185);
nand U13214 (N_13214,N_13042,N_13166);
xor U13215 (N_13215,N_13029,N_13122);
or U13216 (N_13216,N_13058,N_12972);
nand U13217 (N_13217,N_13055,N_13195);
nand U13218 (N_13218,N_13148,N_13068);
nor U13219 (N_13219,N_13013,N_12951);
nand U13220 (N_13220,N_13072,N_13160);
nand U13221 (N_13221,N_13026,N_13192);
xnor U13222 (N_13222,N_12957,N_13045);
nand U13223 (N_13223,N_13048,N_13178);
or U13224 (N_13224,N_13004,N_12908);
or U13225 (N_13225,N_12911,N_13070);
nor U13226 (N_13226,N_12967,N_12956);
xor U13227 (N_13227,N_13001,N_12905);
xnor U13228 (N_13228,N_13125,N_13181);
or U13229 (N_13229,N_13098,N_13096);
or U13230 (N_13230,N_12909,N_13038);
nor U13231 (N_13231,N_12979,N_13071);
xnor U13232 (N_13232,N_13190,N_13082);
or U13233 (N_13233,N_13170,N_13147);
nand U13234 (N_13234,N_13020,N_12953);
xnor U13235 (N_13235,N_13019,N_12974);
xor U13236 (N_13236,N_13134,N_12982);
and U13237 (N_13237,N_13100,N_12938);
nand U13238 (N_13238,N_13069,N_13076);
nor U13239 (N_13239,N_13191,N_13150);
xnor U13240 (N_13240,N_12925,N_13074);
nand U13241 (N_13241,N_13078,N_12916);
or U13242 (N_13242,N_13174,N_12981);
nand U13243 (N_13243,N_12963,N_13129);
nor U13244 (N_13244,N_12961,N_12906);
or U13245 (N_13245,N_12936,N_12943);
nand U13246 (N_13246,N_13135,N_13139);
nand U13247 (N_13247,N_13163,N_13094);
nor U13248 (N_13248,N_13176,N_13054);
nor U13249 (N_13249,N_13154,N_12992);
and U13250 (N_13250,N_13117,N_12903);
or U13251 (N_13251,N_13093,N_13080);
nand U13252 (N_13252,N_13051,N_13012);
xnor U13253 (N_13253,N_13035,N_12940);
nor U13254 (N_13254,N_12937,N_13011);
and U13255 (N_13255,N_13025,N_13091);
and U13256 (N_13256,N_13112,N_13073);
or U13257 (N_13257,N_13046,N_13032);
nor U13258 (N_13258,N_12988,N_13034);
xor U13259 (N_13259,N_13107,N_13108);
xnor U13260 (N_13260,N_13126,N_13059);
and U13261 (N_13261,N_12954,N_13161);
xor U13262 (N_13262,N_12971,N_13153);
xnor U13263 (N_13263,N_13196,N_13077);
xor U13264 (N_13264,N_13050,N_12922);
nand U13265 (N_13265,N_12995,N_13111);
xor U13266 (N_13266,N_12977,N_13156);
nand U13267 (N_13267,N_13007,N_13079);
and U13268 (N_13268,N_12902,N_12976);
and U13269 (N_13269,N_12920,N_12942);
nand U13270 (N_13270,N_13124,N_13017);
or U13271 (N_13271,N_13182,N_13056);
nor U13272 (N_13272,N_13131,N_13052);
xnor U13273 (N_13273,N_13092,N_13120);
or U13274 (N_13274,N_13036,N_13016);
nand U13275 (N_13275,N_13173,N_12928);
nor U13276 (N_13276,N_13133,N_12907);
or U13277 (N_13277,N_13060,N_13066);
or U13278 (N_13278,N_12978,N_12919);
or U13279 (N_13279,N_12939,N_13137);
nor U13280 (N_13280,N_13141,N_13027);
and U13281 (N_13281,N_13087,N_12900);
nor U13282 (N_13282,N_13194,N_13062);
and U13283 (N_13283,N_13104,N_13047);
or U13284 (N_13284,N_12999,N_13198);
and U13285 (N_13285,N_12993,N_12948);
and U13286 (N_13286,N_13116,N_13167);
and U13287 (N_13287,N_13021,N_13023);
and U13288 (N_13288,N_13159,N_13109);
xor U13289 (N_13289,N_13097,N_13099);
nand U13290 (N_13290,N_13063,N_12941);
xnor U13291 (N_13291,N_12947,N_13088);
xnor U13292 (N_13292,N_13101,N_13164);
nand U13293 (N_13293,N_12952,N_13118);
and U13294 (N_13294,N_12998,N_12986);
nand U13295 (N_13295,N_13018,N_12915);
or U13296 (N_13296,N_12912,N_13142);
nor U13297 (N_13297,N_13193,N_13197);
xnor U13298 (N_13298,N_12926,N_12970);
nand U13299 (N_13299,N_13028,N_13138);
nand U13300 (N_13300,N_12964,N_12968);
nand U13301 (N_13301,N_13002,N_12934);
and U13302 (N_13302,N_13188,N_12918);
and U13303 (N_13303,N_13119,N_12984);
xnor U13304 (N_13304,N_13151,N_13010);
xnor U13305 (N_13305,N_12973,N_12965);
nand U13306 (N_13306,N_13168,N_12904);
nor U13307 (N_13307,N_12962,N_12932);
or U13308 (N_13308,N_13113,N_13030);
nand U13309 (N_13309,N_12990,N_12914);
or U13310 (N_13310,N_13086,N_13005);
or U13311 (N_13311,N_13144,N_13095);
and U13312 (N_13312,N_13140,N_12935);
nand U13313 (N_13313,N_13165,N_13162);
or U13314 (N_13314,N_12929,N_13136);
nand U13315 (N_13315,N_13199,N_12949);
or U13316 (N_13316,N_12901,N_13022);
nand U13317 (N_13317,N_13057,N_12980);
or U13318 (N_13318,N_12933,N_13031);
and U13319 (N_13319,N_12959,N_13053);
nand U13320 (N_13320,N_13039,N_13043);
and U13321 (N_13321,N_12966,N_12987);
or U13322 (N_13322,N_13169,N_12944);
or U13323 (N_13323,N_13105,N_13009);
or U13324 (N_13324,N_12927,N_13089);
and U13325 (N_13325,N_13158,N_13172);
nand U13326 (N_13326,N_13024,N_13008);
and U13327 (N_13327,N_13044,N_12960);
and U13328 (N_13328,N_13102,N_13041);
or U13329 (N_13329,N_13121,N_12917);
nor U13330 (N_13330,N_12996,N_12994);
xor U13331 (N_13331,N_13180,N_13145);
nor U13332 (N_13332,N_13003,N_12946);
nand U13333 (N_13333,N_13014,N_13000);
nand U13334 (N_13334,N_13090,N_12955);
nor U13335 (N_13335,N_12945,N_12989);
or U13336 (N_13336,N_13075,N_13114);
nand U13337 (N_13337,N_12923,N_13152);
nand U13338 (N_13338,N_13171,N_13123);
xor U13339 (N_13339,N_12910,N_13081);
nand U13340 (N_13340,N_13186,N_13067);
xor U13341 (N_13341,N_13085,N_12997);
and U13342 (N_13342,N_13033,N_13106);
nand U13343 (N_13343,N_13127,N_12983);
xnor U13344 (N_13344,N_13064,N_13175);
xnor U13345 (N_13345,N_13061,N_13037);
nor U13346 (N_13346,N_12913,N_12950);
xor U13347 (N_13347,N_13006,N_13128);
nor U13348 (N_13348,N_12969,N_13187);
nand U13349 (N_13349,N_13110,N_13083);
nor U13350 (N_13350,N_12994,N_12931);
nor U13351 (N_13351,N_12955,N_13088);
or U13352 (N_13352,N_12999,N_12913);
nand U13353 (N_13353,N_12939,N_13138);
and U13354 (N_13354,N_13171,N_13014);
xor U13355 (N_13355,N_13038,N_12975);
nand U13356 (N_13356,N_13078,N_12955);
or U13357 (N_13357,N_12922,N_13183);
nand U13358 (N_13358,N_13095,N_12997);
and U13359 (N_13359,N_13025,N_12958);
xor U13360 (N_13360,N_13056,N_13014);
nor U13361 (N_13361,N_13193,N_12975);
nor U13362 (N_13362,N_12965,N_12968);
or U13363 (N_13363,N_13091,N_13199);
xnor U13364 (N_13364,N_13054,N_12950);
nand U13365 (N_13365,N_13193,N_12952);
and U13366 (N_13366,N_13109,N_12908);
or U13367 (N_13367,N_13146,N_13156);
and U13368 (N_13368,N_12950,N_12924);
nor U13369 (N_13369,N_12919,N_13020);
or U13370 (N_13370,N_13083,N_13141);
or U13371 (N_13371,N_12916,N_12954);
nand U13372 (N_13372,N_13005,N_12929);
and U13373 (N_13373,N_12907,N_13119);
xor U13374 (N_13374,N_13040,N_13083);
xnor U13375 (N_13375,N_12973,N_13128);
and U13376 (N_13376,N_13088,N_13099);
nand U13377 (N_13377,N_12981,N_13088);
and U13378 (N_13378,N_13153,N_13188);
nand U13379 (N_13379,N_12984,N_13053);
and U13380 (N_13380,N_12944,N_13032);
and U13381 (N_13381,N_12985,N_13147);
nor U13382 (N_13382,N_13056,N_13076);
or U13383 (N_13383,N_13132,N_13083);
nand U13384 (N_13384,N_13000,N_13173);
nor U13385 (N_13385,N_12980,N_13197);
nor U13386 (N_13386,N_13021,N_12901);
or U13387 (N_13387,N_13115,N_13128);
nor U13388 (N_13388,N_12927,N_13064);
xnor U13389 (N_13389,N_13166,N_12966);
and U13390 (N_13390,N_13002,N_12976);
xor U13391 (N_13391,N_12928,N_13053);
xnor U13392 (N_13392,N_13193,N_13117);
and U13393 (N_13393,N_12942,N_13011);
xnor U13394 (N_13394,N_13182,N_12987);
and U13395 (N_13395,N_13089,N_13186);
nor U13396 (N_13396,N_13101,N_13126);
nor U13397 (N_13397,N_13000,N_13029);
and U13398 (N_13398,N_13076,N_13017);
nand U13399 (N_13399,N_13153,N_13021);
xnor U13400 (N_13400,N_13193,N_13006);
nand U13401 (N_13401,N_12969,N_12991);
nand U13402 (N_13402,N_12976,N_12908);
or U13403 (N_13403,N_12981,N_12930);
xnor U13404 (N_13404,N_13116,N_13141);
nand U13405 (N_13405,N_13038,N_13062);
nor U13406 (N_13406,N_13028,N_13024);
nand U13407 (N_13407,N_12987,N_13191);
and U13408 (N_13408,N_13185,N_13197);
or U13409 (N_13409,N_12911,N_13138);
nand U13410 (N_13410,N_13002,N_12942);
or U13411 (N_13411,N_12921,N_13111);
nor U13412 (N_13412,N_13134,N_12997);
nand U13413 (N_13413,N_13132,N_13194);
or U13414 (N_13414,N_13068,N_12931);
nand U13415 (N_13415,N_13100,N_13023);
nand U13416 (N_13416,N_12936,N_13078);
nor U13417 (N_13417,N_12998,N_12995);
or U13418 (N_13418,N_13125,N_13173);
nand U13419 (N_13419,N_13178,N_13148);
nand U13420 (N_13420,N_13185,N_13021);
or U13421 (N_13421,N_12958,N_12903);
xnor U13422 (N_13422,N_12963,N_12938);
nor U13423 (N_13423,N_13059,N_13025);
nor U13424 (N_13424,N_13076,N_13119);
or U13425 (N_13425,N_12916,N_12960);
xor U13426 (N_13426,N_13096,N_13056);
xor U13427 (N_13427,N_13062,N_13193);
nand U13428 (N_13428,N_12919,N_13157);
nor U13429 (N_13429,N_13005,N_12908);
nand U13430 (N_13430,N_12992,N_13066);
nor U13431 (N_13431,N_13005,N_13155);
or U13432 (N_13432,N_12966,N_12958);
or U13433 (N_13433,N_13169,N_13057);
and U13434 (N_13434,N_12999,N_13188);
xnor U13435 (N_13435,N_13196,N_13059);
nor U13436 (N_13436,N_13017,N_13090);
nand U13437 (N_13437,N_13001,N_13048);
xnor U13438 (N_13438,N_13088,N_13170);
xor U13439 (N_13439,N_12918,N_12932);
xor U13440 (N_13440,N_13032,N_13160);
nor U13441 (N_13441,N_13042,N_13116);
xor U13442 (N_13442,N_12963,N_12998);
and U13443 (N_13443,N_13118,N_13093);
nor U13444 (N_13444,N_13116,N_13099);
xnor U13445 (N_13445,N_13059,N_13155);
nand U13446 (N_13446,N_13025,N_12952);
or U13447 (N_13447,N_13150,N_12966);
nand U13448 (N_13448,N_13098,N_13155);
or U13449 (N_13449,N_13055,N_12984);
or U13450 (N_13450,N_13048,N_13111);
or U13451 (N_13451,N_12919,N_13119);
and U13452 (N_13452,N_13035,N_13108);
xnor U13453 (N_13453,N_13157,N_12971);
nor U13454 (N_13454,N_13168,N_13186);
nand U13455 (N_13455,N_12905,N_12914);
and U13456 (N_13456,N_12900,N_12962);
nor U13457 (N_13457,N_13032,N_13152);
nand U13458 (N_13458,N_13192,N_13067);
or U13459 (N_13459,N_12991,N_13185);
or U13460 (N_13460,N_12983,N_13150);
nand U13461 (N_13461,N_12994,N_12986);
nor U13462 (N_13462,N_13178,N_13110);
and U13463 (N_13463,N_12978,N_13072);
and U13464 (N_13464,N_13018,N_13172);
nand U13465 (N_13465,N_13014,N_13119);
xor U13466 (N_13466,N_12989,N_13085);
nor U13467 (N_13467,N_13158,N_13177);
nor U13468 (N_13468,N_13116,N_12960);
xor U13469 (N_13469,N_13023,N_13133);
xor U13470 (N_13470,N_13004,N_13038);
and U13471 (N_13471,N_13089,N_12929);
and U13472 (N_13472,N_13132,N_13003);
nor U13473 (N_13473,N_12923,N_13178);
and U13474 (N_13474,N_12917,N_12990);
or U13475 (N_13475,N_12942,N_13056);
nand U13476 (N_13476,N_13186,N_13120);
and U13477 (N_13477,N_13157,N_13159);
xor U13478 (N_13478,N_13165,N_12943);
nor U13479 (N_13479,N_13147,N_13123);
and U13480 (N_13480,N_13180,N_12980);
and U13481 (N_13481,N_13034,N_13099);
xor U13482 (N_13482,N_13105,N_13035);
nor U13483 (N_13483,N_12943,N_12955);
nand U13484 (N_13484,N_13099,N_12952);
and U13485 (N_13485,N_13138,N_13073);
nand U13486 (N_13486,N_13059,N_13027);
xnor U13487 (N_13487,N_12961,N_13062);
and U13488 (N_13488,N_13030,N_13009);
nor U13489 (N_13489,N_13197,N_13094);
and U13490 (N_13490,N_13147,N_13095);
nor U13491 (N_13491,N_12969,N_13042);
or U13492 (N_13492,N_12932,N_12953);
and U13493 (N_13493,N_13143,N_12966);
and U13494 (N_13494,N_13061,N_13134);
xor U13495 (N_13495,N_13092,N_13134);
and U13496 (N_13496,N_13057,N_13004);
or U13497 (N_13497,N_13063,N_13165);
and U13498 (N_13498,N_12916,N_12914);
nor U13499 (N_13499,N_13066,N_12956);
or U13500 (N_13500,N_13276,N_13334);
nand U13501 (N_13501,N_13275,N_13365);
nand U13502 (N_13502,N_13303,N_13309);
and U13503 (N_13503,N_13496,N_13469);
nor U13504 (N_13504,N_13206,N_13467);
and U13505 (N_13505,N_13456,N_13476);
nand U13506 (N_13506,N_13489,N_13434);
nor U13507 (N_13507,N_13201,N_13391);
nand U13508 (N_13508,N_13253,N_13335);
xor U13509 (N_13509,N_13293,N_13242);
or U13510 (N_13510,N_13422,N_13319);
nor U13511 (N_13511,N_13485,N_13423);
or U13512 (N_13512,N_13397,N_13401);
nor U13513 (N_13513,N_13298,N_13453);
and U13514 (N_13514,N_13271,N_13460);
nand U13515 (N_13515,N_13409,N_13412);
nand U13516 (N_13516,N_13333,N_13246);
or U13517 (N_13517,N_13224,N_13288);
nor U13518 (N_13518,N_13244,N_13277);
and U13519 (N_13519,N_13459,N_13348);
or U13520 (N_13520,N_13465,N_13220);
and U13521 (N_13521,N_13226,N_13321);
xor U13522 (N_13522,N_13233,N_13477);
and U13523 (N_13523,N_13274,N_13358);
or U13524 (N_13524,N_13214,N_13390);
and U13525 (N_13525,N_13320,N_13428);
xor U13526 (N_13526,N_13411,N_13399);
and U13527 (N_13527,N_13331,N_13302);
or U13528 (N_13528,N_13464,N_13458);
or U13529 (N_13529,N_13424,N_13261);
nand U13530 (N_13530,N_13382,N_13340);
and U13531 (N_13531,N_13338,N_13481);
nor U13532 (N_13532,N_13445,N_13497);
or U13533 (N_13533,N_13249,N_13408);
xnor U13534 (N_13534,N_13356,N_13430);
xnor U13535 (N_13535,N_13366,N_13228);
nor U13536 (N_13536,N_13222,N_13360);
nor U13537 (N_13537,N_13429,N_13347);
nor U13538 (N_13538,N_13414,N_13362);
xor U13539 (N_13539,N_13216,N_13452);
or U13540 (N_13540,N_13342,N_13322);
or U13541 (N_13541,N_13223,N_13357);
or U13542 (N_13542,N_13438,N_13234);
xnor U13543 (N_13543,N_13406,N_13323);
or U13544 (N_13544,N_13427,N_13203);
xnor U13545 (N_13545,N_13306,N_13370);
or U13546 (N_13546,N_13364,N_13241);
nand U13547 (N_13547,N_13376,N_13385);
nand U13548 (N_13548,N_13439,N_13260);
or U13549 (N_13549,N_13402,N_13368);
and U13550 (N_13550,N_13446,N_13492);
and U13551 (N_13551,N_13369,N_13432);
or U13552 (N_13552,N_13479,N_13450);
xor U13553 (N_13553,N_13257,N_13248);
xor U13554 (N_13554,N_13351,N_13405);
and U13555 (N_13555,N_13495,N_13332);
nor U13556 (N_13556,N_13404,N_13263);
or U13557 (N_13557,N_13482,N_13202);
nor U13558 (N_13558,N_13316,N_13239);
nand U13559 (N_13559,N_13442,N_13417);
xor U13560 (N_13560,N_13264,N_13484);
nor U13561 (N_13561,N_13250,N_13258);
nand U13562 (N_13562,N_13483,N_13418);
or U13563 (N_13563,N_13251,N_13381);
and U13564 (N_13564,N_13290,N_13294);
nor U13565 (N_13565,N_13426,N_13389);
nand U13566 (N_13566,N_13393,N_13387);
xnor U13567 (N_13567,N_13312,N_13487);
or U13568 (N_13568,N_13448,N_13462);
xnor U13569 (N_13569,N_13235,N_13359);
nand U13570 (N_13570,N_13451,N_13396);
or U13571 (N_13571,N_13295,N_13291);
and U13572 (N_13572,N_13441,N_13210);
or U13573 (N_13573,N_13419,N_13215);
xor U13574 (N_13574,N_13225,N_13243);
and U13575 (N_13575,N_13256,N_13212);
and U13576 (N_13576,N_13415,N_13337);
xor U13577 (N_13577,N_13470,N_13421);
nand U13578 (N_13578,N_13454,N_13493);
or U13579 (N_13579,N_13304,N_13352);
and U13580 (N_13580,N_13204,N_13310);
xor U13581 (N_13581,N_13392,N_13240);
or U13582 (N_13582,N_13284,N_13377);
xnor U13583 (N_13583,N_13217,N_13433);
nand U13584 (N_13584,N_13372,N_13272);
nor U13585 (N_13585,N_13339,N_13336);
nand U13586 (N_13586,N_13361,N_13207);
nor U13587 (N_13587,N_13229,N_13255);
nor U13588 (N_13588,N_13285,N_13488);
or U13589 (N_13589,N_13245,N_13300);
or U13590 (N_13590,N_13211,N_13231);
or U13591 (N_13591,N_13444,N_13394);
or U13592 (N_13592,N_13416,N_13420);
nand U13593 (N_13593,N_13273,N_13341);
and U13594 (N_13594,N_13286,N_13480);
and U13595 (N_13595,N_13498,N_13468);
nand U13596 (N_13596,N_13259,N_13435);
and U13597 (N_13597,N_13281,N_13270);
nand U13598 (N_13598,N_13324,N_13205);
nand U13599 (N_13599,N_13326,N_13478);
xnor U13600 (N_13600,N_13328,N_13330);
or U13601 (N_13601,N_13314,N_13374);
nand U13602 (N_13602,N_13471,N_13311);
and U13603 (N_13603,N_13209,N_13344);
nand U13604 (N_13604,N_13349,N_13236);
nand U13605 (N_13605,N_13279,N_13386);
xnor U13606 (N_13606,N_13254,N_13218);
xnor U13607 (N_13607,N_13289,N_13317);
and U13608 (N_13608,N_13486,N_13373);
nor U13609 (N_13609,N_13230,N_13280);
and U13610 (N_13610,N_13355,N_13473);
nor U13611 (N_13611,N_13327,N_13353);
nand U13612 (N_13612,N_13472,N_13375);
nor U13613 (N_13613,N_13227,N_13395);
nand U13614 (N_13614,N_13449,N_13343);
nor U13615 (N_13615,N_13221,N_13474);
nor U13616 (N_13616,N_13463,N_13305);
nand U13617 (N_13617,N_13268,N_13490);
and U13618 (N_13618,N_13313,N_13266);
or U13619 (N_13619,N_13265,N_13287);
or U13620 (N_13620,N_13237,N_13267);
or U13621 (N_13621,N_13350,N_13213);
or U13622 (N_13622,N_13208,N_13443);
nand U13623 (N_13623,N_13407,N_13346);
or U13624 (N_13624,N_13278,N_13301);
or U13625 (N_13625,N_13283,N_13499);
nor U13626 (N_13626,N_13384,N_13440);
or U13627 (N_13627,N_13345,N_13388);
or U13628 (N_13628,N_13282,N_13410);
xor U13629 (N_13629,N_13219,N_13378);
xnor U13630 (N_13630,N_13457,N_13238);
nand U13631 (N_13631,N_13308,N_13299);
or U13632 (N_13632,N_13367,N_13262);
nand U13633 (N_13633,N_13379,N_13296);
or U13634 (N_13634,N_13425,N_13292);
or U13635 (N_13635,N_13413,N_13232);
nand U13636 (N_13636,N_13475,N_13491);
or U13637 (N_13637,N_13466,N_13315);
xor U13638 (N_13638,N_13247,N_13455);
xnor U13639 (N_13639,N_13363,N_13269);
nand U13640 (N_13640,N_13200,N_13252);
xor U13641 (N_13641,N_13329,N_13494);
and U13642 (N_13642,N_13297,N_13403);
nor U13643 (N_13643,N_13447,N_13325);
nor U13644 (N_13644,N_13400,N_13461);
nor U13645 (N_13645,N_13380,N_13383);
nand U13646 (N_13646,N_13436,N_13318);
or U13647 (N_13647,N_13354,N_13437);
nor U13648 (N_13648,N_13398,N_13431);
or U13649 (N_13649,N_13371,N_13307);
or U13650 (N_13650,N_13390,N_13278);
xnor U13651 (N_13651,N_13263,N_13315);
and U13652 (N_13652,N_13309,N_13271);
and U13653 (N_13653,N_13244,N_13403);
and U13654 (N_13654,N_13349,N_13487);
xor U13655 (N_13655,N_13346,N_13378);
and U13656 (N_13656,N_13428,N_13323);
xnor U13657 (N_13657,N_13274,N_13477);
nand U13658 (N_13658,N_13242,N_13350);
or U13659 (N_13659,N_13483,N_13492);
and U13660 (N_13660,N_13323,N_13264);
xnor U13661 (N_13661,N_13263,N_13370);
nand U13662 (N_13662,N_13400,N_13476);
xnor U13663 (N_13663,N_13375,N_13201);
nor U13664 (N_13664,N_13347,N_13288);
and U13665 (N_13665,N_13430,N_13414);
nand U13666 (N_13666,N_13344,N_13221);
nand U13667 (N_13667,N_13496,N_13251);
xor U13668 (N_13668,N_13275,N_13455);
or U13669 (N_13669,N_13247,N_13239);
nand U13670 (N_13670,N_13432,N_13496);
nor U13671 (N_13671,N_13321,N_13446);
nand U13672 (N_13672,N_13476,N_13293);
or U13673 (N_13673,N_13428,N_13417);
or U13674 (N_13674,N_13235,N_13366);
and U13675 (N_13675,N_13388,N_13224);
nor U13676 (N_13676,N_13218,N_13357);
and U13677 (N_13677,N_13317,N_13439);
or U13678 (N_13678,N_13434,N_13398);
nand U13679 (N_13679,N_13333,N_13301);
nand U13680 (N_13680,N_13384,N_13377);
nand U13681 (N_13681,N_13219,N_13350);
nor U13682 (N_13682,N_13479,N_13492);
xor U13683 (N_13683,N_13337,N_13373);
xnor U13684 (N_13684,N_13460,N_13331);
nor U13685 (N_13685,N_13297,N_13233);
xnor U13686 (N_13686,N_13396,N_13288);
xor U13687 (N_13687,N_13328,N_13379);
or U13688 (N_13688,N_13469,N_13353);
and U13689 (N_13689,N_13319,N_13484);
nand U13690 (N_13690,N_13324,N_13328);
nor U13691 (N_13691,N_13382,N_13210);
nor U13692 (N_13692,N_13492,N_13381);
nand U13693 (N_13693,N_13441,N_13276);
and U13694 (N_13694,N_13302,N_13376);
and U13695 (N_13695,N_13268,N_13329);
or U13696 (N_13696,N_13288,N_13277);
nand U13697 (N_13697,N_13299,N_13486);
xor U13698 (N_13698,N_13444,N_13243);
or U13699 (N_13699,N_13362,N_13393);
and U13700 (N_13700,N_13418,N_13286);
and U13701 (N_13701,N_13436,N_13420);
or U13702 (N_13702,N_13498,N_13316);
nor U13703 (N_13703,N_13242,N_13496);
xnor U13704 (N_13704,N_13315,N_13267);
nor U13705 (N_13705,N_13426,N_13232);
or U13706 (N_13706,N_13283,N_13262);
and U13707 (N_13707,N_13378,N_13361);
and U13708 (N_13708,N_13483,N_13375);
xor U13709 (N_13709,N_13359,N_13285);
nand U13710 (N_13710,N_13404,N_13317);
or U13711 (N_13711,N_13456,N_13256);
nor U13712 (N_13712,N_13385,N_13275);
xor U13713 (N_13713,N_13251,N_13463);
nand U13714 (N_13714,N_13348,N_13238);
or U13715 (N_13715,N_13283,N_13265);
xor U13716 (N_13716,N_13486,N_13264);
nand U13717 (N_13717,N_13424,N_13363);
nand U13718 (N_13718,N_13341,N_13229);
xnor U13719 (N_13719,N_13201,N_13289);
nor U13720 (N_13720,N_13390,N_13482);
or U13721 (N_13721,N_13286,N_13430);
xor U13722 (N_13722,N_13451,N_13406);
nor U13723 (N_13723,N_13285,N_13425);
nand U13724 (N_13724,N_13348,N_13397);
xnor U13725 (N_13725,N_13310,N_13285);
nor U13726 (N_13726,N_13342,N_13390);
xnor U13727 (N_13727,N_13201,N_13404);
and U13728 (N_13728,N_13318,N_13433);
and U13729 (N_13729,N_13248,N_13363);
xnor U13730 (N_13730,N_13294,N_13247);
nand U13731 (N_13731,N_13461,N_13441);
nand U13732 (N_13732,N_13344,N_13287);
or U13733 (N_13733,N_13381,N_13442);
and U13734 (N_13734,N_13244,N_13253);
or U13735 (N_13735,N_13474,N_13230);
or U13736 (N_13736,N_13434,N_13380);
nor U13737 (N_13737,N_13330,N_13227);
nand U13738 (N_13738,N_13215,N_13387);
nand U13739 (N_13739,N_13255,N_13288);
nand U13740 (N_13740,N_13446,N_13441);
and U13741 (N_13741,N_13340,N_13433);
xor U13742 (N_13742,N_13202,N_13486);
xnor U13743 (N_13743,N_13204,N_13227);
nor U13744 (N_13744,N_13410,N_13376);
xor U13745 (N_13745,N_13496,N_13454);
or U13746 (N_13746,N_13480,N_13321);
nor U13747 (N_13747,N_13322,N_13368);
nand U13748 (N_13748,N_13279,N_13246);
and U13749 (N_13749,N_13392,N_13331);
and U13750 (N_13750,N_13383,N_13273);
and U13751 (N_13751,N_13409,N_13450);
and U13752 (N_13752,N_13264,N_13332);
nor U13753 (N_13753,N_13426,N_13290);
or U13754 (N_13754,N_13314,N_13462);
and U13755 (N_13755,N_13494,N_13259);
nor U13756 (N_13756,N_13431,N_13495);
and U13757 (N_13757,N_13349,N_13359);
or U13758 (N_13758,N_13445,N_13288);
xnor U13759 (N_13759,N_13226,N_13434);
or U13760 (N_13760,N_13447,N_13286);
nand U13761 (N_13761,N_13330,N_13331);
xor U13762 (N_13762,N_13410,N_13356);
nor U13763 (N_13763,N_13315,N_13479);
nand U13764 (N_13764,N_13296,N_13226);
xnor U13765 (N_13765,N_13389,N_13221);
nand U13766 (N_13766,N_13463,N_13277);
nand U13767 (N_13767,N_13413,N_13409);
and U13768 (N_13768,N_13423,N_13402);
nand U13769 (N_13769,N_13393,N_13499);
xnor U13770 (N_13770,N_13442,N_13412);
nor U13771 (N_13771,N_13498,N_13393);
or U13772 (N_13772,N_13220,N_13266);
or U13773 (N_13773,N_13289,N_13254);
xnor U13774 (N_13774,N_13377,N_13279);
nand U13775 (N_13775,N_13260,N_13358);
or U13776 (N_13776,N_13306,N_13405);
nand U13777 (N_13777,N_13293,N_13287);
or U13778 (N_13778,N_13270,N_13445);
nand U13779 (N_13779,N_13385,N_13240);
or U13780 (N_13780,N_13252,N_13407);
xnor U13781 (N_13781,N_13228,N_13374);
xor U13782 (N_13782,N_13217,N_13349);
and U13783 (N_13783,N_13273,N_13259);
nand U13784 (N_13784,N_13378,N_13474);
or U13785 (N_13785,N_13433,N_13329);
nand U13786 (N_13786,N_13354,N_13268);
nor U13787 (N_13787,N_13242,N_13219);
and U13788 (N_13788,N_13308,N_13345);
nor U13789 (N_13789,N_13346,N_13225);
and U13790 (N_13790,N_13294,N_13272);
nor U13791 (N_13791,N_13337,N_13248);
nand U13792 (N_13792,N_13305,N_13279);
or U13793 (N_13793,N_13387,N_13304);
xor U13794 (N_13794,N_13335,N_13460);
xnor U13795 (N_13795,N_13205,N_13469);
nand U13796 (N_13796,N_13316,N_13341);
nor U13797 (N_13797,N_13402,N_13269);
nand U13798 (N_13798,N_13441,N_13495);
or U13799 (N_13799,N_13468,N_13481);
nand U13800 (N_13800,N_13786,N_13641);
xor U13801 (N_13801,N_13567,N_13726);
nor U13802 (N_13802,N_13523,N_13662);
and U13803 (N_13803,N_13561,N_13748);
nand U13804 (N_13804,N_13642,N_13649);
and U13805 (N_13805,N_13608,N_13627);
xnor U13806 (N_13806,N_13672,N_13795);
xnor U13807 (N_13807,N_13724,N_13626);
nand U13808 (N_13808,N_13751,N_13777);
xor U13809 (N_13809,N_13666,N_13535);
xnor U13810 (N_13810,N_13643,N_13583);
xor U13811 (N_13811,N_13699,N_13656);
or U13812 (N_13812,N_13698,N_13543);
and U13813 (N_13813,N_13651,N_13782);
and U13814 (N_13814,N_13611,N_13779);
and U13815 (N_13815,N_13771,N_13585);
or U13816 (N_13816,N_13640,N_13791);
nand U13817 (N_13817,N_13580,N_13784);
xor U13818 (N_13818,N_13624,N_13680);
xnor U13819 (N_13819,N_13638,N_13575);
or U13820 (N_13820,N_13703,N_13647);
nor U13821 (N_13821,N_13673,N_13716);
xor U13822 (N_13822,N_13667,N_13740);
or U13823 (N_13823,N_13658,N_13617);
xnor U13824 (N_13824,N_13581,N_13516);
nor U13825 (N_13825,N_13669,N_13646);
nand U13826 (N_13826,N_13765,N_13548);
and U13827 (N_13827,N_13592,N_13606);
xnor U13828 (N_13828,N_13616,N_13780);
nor U13829 (N_13829,N_13732,N_13720);
or U13830 (N_13830,N_13700,N_13714);
xor U13831 (N_13831,N_13533,N_13584);
or U13832 (N_13832,N_13718,N_13729);
or U13833 (N_13833,N_13601,N_13573);
or U13834 (N_13834,N_13564,N_13562);
nor U13835 (N_13835,N_13572,N_13644);
and U13836 (N_13836,N_13798,N_13752);
nor U13837 (N_13837,N_13660,N_13773);
nand U13838 (N_13838,N_13538,N_13540);
or U13839 (N_13839,N_13534,N_13770);
nand U13840 (N_13840,N_13633,N_13736);
or U13841 (N_13841,N_13735,N_13509);
or U13842 (N_13842,N_13514,N_13503);
xor U13843 (N_13843,N_13655,N_13521);
nand U13844 (N_13844,N_13557,N_13554);
or U13845 (N_13845,N_13505,N_13518);
nor U13846 (N_13846,N_13719,N_13674);
nand U13847 (N_13847,N_13625,N_13750);
nor U13848 (N_13848,N_13539,N_13595);
nand U13849 (N_13849,N_13727,N_13659);
and U13850 (N_13850,N_13639,N_13525);
nand U13851 (N_13851,N_13688,N_13734);
nor U13852 (N_13852,N_13717,N_13621);
xnor U13853 (N_13853,N_13747,N_13565);
or U13854 (N_13854,N_13531,N_13527);
or U13855 (N_13855,N_13749,N_13733);
and U13856 (N_13856,N_13737,N_13728);
or U13857 (N_13857,N_13789,N_13781);
nor U13858 (N_13858,N_13663,N_13690);
nand U13859 (N_13859,N_13787,N_13578);
or U13860 (N_13860,N_13632,N_13774);
xnor U13861 (N_13861,N_13559,N_13522);
or U13862 (N_13862,N_13671,N_13731);
or U13863 (N_13863,N_13507,N_13610);
nor U13864 (N_13864,N_13511,N_13555);
or U13865 (N_13865,N_13574,N_13614);
nor U13866 (N_13866,N_13678,N_13652);
and U13867 (N_13867,N_13725,N_13618);
and U13868 (N_13868,N_13796,N_13504);
nor U13869 (N_13869,N_13593,N_13687);
and U13870 (N_13870,N_13605,N_13730);
xor U13871 (N_13871,N_13705,N_13545);
nand U13872 (N_13872,N_13530,N_13582);
or U13873 (N_13873,N_13694,N_13775);
nand U13874 (N_13874,N_13742,N_13586);
xor U13875 (N_13875,N_13609,N_13682);
nor U13876 (N_13876,N_13500,N_13541);
or U13877 (N_13877,N_13689,N_13739);
nor U13878 (N_13878,N_13710,N_13706);
nand U13879 (N_13879,N_13723,N_13677);
nand U13880 (N_13880,N_13772,N_13715);
and U13881 (N_13881,N_13570,N_13697);
nand U13882 (N_13882,N_13546,N_13692);
xor U13883 (N_13883,N_13515,N_13569);
nand U13884 (N_13884,N_13704,N_13607);
nand U13885 (N_13885,N_13708,N_13799);
or U13886 (N_13886,N_13746,N_13758);
nand U13887 (N_13887,N_13637,N_13743);
and U13888 (N_13888,N_13517,N_13686);
or U13889 (N_13889,N_13679,N_13602);
nor U13890 (N_13890,N_13579,N_13634);
and U13891 (N_13891,N_13664,N_13685);
xor U13892 (N_13892,N_13510,N_13577);
xor U13893 (N_13893,N_13604,N_13793);
xnor U13894 (N_13894,N_13630,N_13506);
nand U13895 (N_13895,N_13785,N_13760);
or U13896 (N_13896,N_13612,N_13513);
nand U13897 (N_13897,N_13587,N_13741);
or U13898 (N_13898,N_13670,N_13753);
nand U13899 (N_13899,N_13738,N_13576);
and U13900 (N_13900,N_13589,N_13566);
and U13901 (N_13901,N_13681,N_13754);
nor U13902 (N_13902,N_13790,N_13757);
nand U13903 (N_13903,N_13620,N_13502);
nor U13904 (N_13904,N_13598,N_13556);
nor U13905 (N_13905,N_13615,N_13544);
and U13906 (N_13906,N_13675,N_13721);
nand U13907 (N_13907,N_13501,N_13661);
or U13908 (N_13908,N_13600,N_13768);
nor U13909 (N_13909,N_13693,N_13769);
nor U13910 (N_13910,N_13532,N_13519);
xor U13911 (N_13911,N_13524,N_13650);
or U13912 (N_13912,N_13744,N_13713);
nand U13913 (N_13913,N_13696,N_13701);
xnor U13914 (N_13914,N_13657,N_13529);
and U13915 (N_13915,N_13684,N_13756);
xor U13916 (N_13916,N_13776,N_13702);
and U13917 (N_13917,N_13613,N_13635);
or U13918 (N_13918,N_13794,N_13745);
xor U13919 (N_13919,N_13591,N_13767);
xnor U13920 (N_13920,N_13512,N_13653);
xnor U13921 (N_13921,N_13542,N_13792);
or U13922 (N_13922,N_13526,N_13631);
and U13923 (N_13923,N_13588,N_13665);
nor U13924 (N_13924,N_13766,N_13551);
or U13925 (N_13925,N_13628,N_13648);
or U13926 (N_13926,N_13619,N_13560);
and U13927 (N_13927,N_13629,N_13508);
and U13928 (N_13928,N_13783,N_13528);
nor U13929 (N_13929,N_13563,N_13764);
nor U13930 (N_13930,N_13711,N_13558);
nor U13931 (N_13931,N_13603,N_13761);
or U13932 (N_13932,N_13778,N_13712);
xor U13933 (N_13933,N_13549,N_13683);
xnor U13934 (N_13934,N_13668,N_13691);
nand U13935 (N_13935,N_13536,N_13571);
nand U13936 (N_13936,N_13788,N_13645);
nand U13937 (N_13937,N_13707,N_13520);
nand U13938 (N_13938,N_13654,N_13599);
xor U13939 (N_13939,N_13759,N_13636);
xnor U13940 (N_13940,N_13590,N_13797);
xor U13941 (N_13941,N_13762,N_13622);
xor U13942 (N_13942,N_13553,N_13755);
or U13943 (N_13943,N_13597,N_13552);
xnor U13944 (N_13944,N_13568,N_13695);
nand U13945 (N_13945,N_13537,N_13676);
or U13946 (N_13946,N_13547,N_13722);
nand U13947 (N_13947,N_13596,N_13594);
nor U13948 (N_13948,N_13709,N_13763);
nand U13949 (N_13949,N_13550,N_13623);
nand U13950 (N_13950,N_13685,N_13502);
and U13951 (N_13951,N_13791,N_13785);
or U13952 (N_13952,N_13594,N_13532);
xnor U13953 (N_13953,N_13654,N_13722);
nand U13954 (N_13954,N_13659,N_13653);
or U13955 (N_13955,N_13771,N_13679);
nand U13956 (N_13956,N_13741,N_13638);
xor U13957 (N_13957,N_13571,N_13797);
and U13958 (N_13958,N_13646,N_13555);
or U13959 (N_13959,N_13530,N_13614);
or U13960 (N_13960,N_13514,N_13796);
xor U13961 (N_13961,N_13689,N_13778);
xor U13962 (N_13962,N_13668,N_13743);
nand U13963 (N_13963,N_13721,N_13541);
nor U13964 (N_13964,N_13790,N_13731);
nand U13965 (N_13965,N_13677,N_13694);
or U13966 (N_13966,N_13756,N_13699);
and U13967 (N_13967,N_13509,N_13611);
nand U13968 (N_13968,N_13557,N_13770);
xnor U13969 (N_13969,N_13662,N_13734);
nand U13970 (N_13970,N_13537,N_13701);
nand U13971 (N_13971,N_13735,N_13633);
nor U13972 (N_13972,N_13562,N_13533);
nor U13973 (N_13973,N_13606,N_13614);
or U13974 (N_13974,N_13663,N_13513);
nand U13975 (N_13975,N_13696,N_13763);
nor U13976 (N_13976,N_13583,N_13678);
and U13977 (N_13977,N_13603,N_13684);
nand U13978 (N_13978,N_13539,N_13749);
and U13979 (N_13979,N_13621,N_13558);
nor U13980 (N_13980,N_13733,N_13548);
xor U13981 (N_13981,N_13762,N_13579);
and U13982 (N_13982,N_13790,N_13524);
xnor U13983 (N_13983,N_13638,N_13729);
nand U13984 (N_13984,N_13547,N_13563);
and U13985 (N_13985,N_13623,N_13647);
nand U13986 (N_13986,N_13630,N_13649);
xnor U13987 (N_13987,N_13726,N_13615);
or U13988 (N_13988,N_13500,N_13744);
or U13989 (N_13989,N_13757,N_13528);
xnor U13990 (N_13990,N_13749,N_13635);
xnor U13991 (N_13991,N_13516,N_13528);
nand U13992 (N_13992,N_13578,N_13517);
nand U13993 (N_13993,N_13748,N_13727);
nand U13994 (N_13994,N_13752,N_13655);
nand U13995 (N_13995,N_13684,N_13631);
and U13996 (N_13996,N_13579,N_13626);
nand U13997 (N_13997,N_13518,N_13615);
or U13998 (N_13998,N_13693,N_13764);
and U13999 (N_13999,N_13761,N_13593);
nand U14000 (N_14000,N_13735,N_13598);
nor U14001 (N_14001,N_13748,N_13553);
or U14002 (N_14002,N_13515,N_13751);
nor U14003 (N_14003,N_13678,N_13682);
nand U14004 (N_14004,N_13586,N_13587);
xor U14005 (N_14005,N_13504,N_13728);
and U14006 (N_14006,N_13740,N_13678);
xnor U14007 (N_14007,N_13768,N_13736);
xnor U14008 (N_14008,N_13506,N_13667);
and U14009 (N_14009,N_13665,N_13550);
and U14010 (N_14010,N_13559,N_13761);
nor U14011 (N_14011,N_13742,N_13650);
xnor U14012 (N_14012,N_13562,N_13729);
and U14013 (N_14013,N_13677,N_13762);
and U14014 (N_14014,N_13691,N_13615);
nor U14015 (N_14015,N_13589,N_13525);
xor U14016 (N_14016,N_13566,N_13680);
nand U14017 (N_14017,N_13650,N_13576);
and U14018 (N_14018,N_13737,N_13773);
nor U14019 (N_14019,N_13728,N_13744);
xor U14020 (N_14020,N_13729,N_13628);
and U14021 (N_14021,N_13512,N_13626);
or U14022 (N_14022,N_13600,N_13558);
or U14023 (N_14023,N_13787,N_13547);
and U14024 (N_14024,N_13725,N_13502);
and U14025 (N_14025,N_13535,N_13586);
nor U14026 (N_14026,N_13665,N_13533);
nand U14027 (N_14027,N_13730,N_13713);
or U14028 (N_14028,N_13522,N_13682);
and U14029 (N_14029,N_13640,N_13754);
xnor U14030 (N_14030,N_13679,N_13580);
nor U14031 (N_14031,N_13548,N_13564);
xnor U14032 (N_14032,N_13662,N_13625);
nor U14033 (N_14033,N_13621,N_13502);
nand U14034 (N_14034,N_13554,N_13747);
nor U14035 (N_14035,N_13780,N_13617);
nand U14036 (N_14036,N_13790,N_13628);
nand U14037 (N_14037,N_13674,N_13736);
nand U14038 (N_14038,N_13689,N_13731);
nor U14039 (N_14039,N_13580,N_13742);
nand U14040 (N_14040,N_13700,N_13649);
nor U14041 (N_14041,N_13506,N_13793);
or U14042 (N_14042,N_13637,N_13578);
or U14043 (N_14043,N_13603,N_13654);
xnor U14044 (N_14044,N_13568,N_13790);
or U14045 (N_14045,N_13539,N_13574);
nor U14046 (N_14046,N_13656,N_13694);
or U14047 (N_14047,N_13741,N_13508);
nand U14048 (N_14048,N_13525,N_13697);
nor U14049 (N_14049,N_13642,N_13652);
and U14050 (N_14050,N_13659,N_13795);
and U14051 (N_14051,N_13613,N_13790);
nor U14052 (N_14052,N_13703,N_13637);
or U14053 (N_14053,N_13562,N_13617);
or U14054 (N_14054,N_13523,N_13665);
xnor U14055 (N_14055,N_13773,N_13644);
xor U14056 (N_14056,N_13758,N_13782);
or U14057 (N_14057,N_13505,N_13747);
nor U14058 (N_14058,N_13514,N_13751);
and U14059 (N_14059,N_13727,N_13565);
nor U14060 (N_14060,N_13723,N_13538);
xor U14061 (N_14061,N_13564,N_13587);
or U14062 (N_14062,N_13534,N_13574);
xor U14063 (N_14063,N_13649,N_13580);
nand U14064 (N_14064,N_13504,N_13586);
and U14065 (N_14065,N_13788,N_13577);
xnor U14066 (N_14066,N_13698,N_13581);
and U14067 (N_14067,N_13773,N_13702);
and U14068 (N_14068,N_13651,N_13545);
nor U14069 (N_14069,N_13682,N_13502);
nor U14070 (N_14070,N_13533,N_13668);
nand U14071 (N_14071,N_13527,N_13552);
xnor U14072 (N_14072,N_13709,N_13646);
xor U14073 (N_14073,N_13531,N_13749);
and U14074 (N_14074,N_13671,N_13783);
and U14075 (N_14075,N_13667,N_13744);
nand U14076 (N_14076,N_13600,N_13774);
nand U14077 (N_14077,N_13674,N_13596);
nor U14078 (N_14078,N_13731,N_13531);
nor U14079 (N_14079,N_13708,N_13621);
or U14080 (N_14080,N_13726,N_13559);
nor U14081 (N_14081,N_13738,N_13636);
nand U14082 (N_14082,N_13520,N_13531);
nand U14083 (N_14083,N_13716,N_13785);
nand U14084 (N_14084,N_13706,N_13762);
xnor U14085 (N_14085,N_13794,N_13605);
nand U14086 (N_14086,N_13659,N_13660);
or U14087 (N_14087,N_13559,N_13780);
or U14088 (N_14088,N_13578,N_13627);
and U14089 (N_14089,N_13555,N_13759);
nor U14090 (N_14090,N_13588,N_13621);
and U14091 (N_14091,N_13599,N_13662);
nor U14092 (N_14092,N_13643,N_13632);
nor U14093 (N_14093,N_13721,N_13680);
xnor U14094 (N_14094,N_13673,N_13747);
or U14095 (N_14095,N_13621,N_13684);
and U14096 (N_14096,N_13770,N_13796);
nand U14097 (N_14097,N_13669,N_13680);
and U14098 (N_14098,N_13559,N_13570);
or U14099 (N_14099,N_13514,N_13745);
and U14100 (N_14100,N_13824,N_13890);
and U14101 (N_14101,N_14063,N_13961);
xor U14102 (N_14102,N_13968,N_14067);
xor U14103 (N_14103,N_13997,N_13981);
and U14104 (N_14104,N_13901,N_13918);
nand U14105 (N_14105,N_13831,N_14056);
and U14106 (N_14106,N_14009,N_14049);
nor U14107 (N_14107,N_13904,N_14007);
xnor U14108 (N_14108,N_14059,N_14035);
or U14109 (N_14109,N_13946,N_14077);
nand U14110 (N_14110,N_13810,N_13875);
and U14111 (N_14111,N_14078,N_13995);
nand U14112 (N_14112,N_13923,N_14000);
nor U14113 (N_14113,N_13958,N_13801);
nand U14114 (N_14114,N_13922,N_13917);
nand U14115 (N_14115,N_14031,N_13838);
nor U14116 (N_14116,N_14083,N_14079);
and U14117 (N_14117,N_14019,N_13883);
nor U14118 (N_14118,N_14036,N_13899);
nand U14119 (N_14119,N_14095,N_13873);
nand U14120 (N_14120,N_14068,N_13879);
nor U14121 (N_14121,N_14062,N_13842);
and U14122 (N_14122,N_13955,N_14010);
nor U14123 (N_14123,N_13983,N_13942);
nand U14124 (N_14124,N_14005,N_14037);
nand U14125 (N_14125,N_13945,N_14070);
nor U14126 (N_14126,N_13884,N_13889);
or U14127 (N_14127,N_14042,N_13856);
xor U14128 (N_14128,N_13866,N_13975);
nor U14129 (N_14129,N_13972,N_14050);
xor U14130 (N_14130,N_13966,N_13967);
or U14131 (N_14131,N_13869,N_14020);
and U14132 (N_14132,N_14055,N_13881);
or U14133 (N_14133,N_13862,N_13926);
or U14134 (N_14134,N_13982,N_13986);
or U14135 (N_14135,N_13872,N_13988);
nor U14136 (N_14136,N_14091,N_14014);
xnor U14137 (N_14137,N_13885,N_14034);
nand U14138 (N_14138,N_13809,N_13932);
or U14139 (N_14139,N_14045,N_13974);
nor U14140 (N_14140,N_13978,N_14013);
or U14141 (N_14141,N_13839,N_13950);
xnor U14142 (N_14142,N_13925,N_13854);
xor U14143 (N_14143,N_13800,N_14002);
xor U14144 (N_14144,N_13808,N_14053);
and U14145 (N_14145,N_13934,N_13857);
nor U14146 (N_14146,N_13912,N_13980);
xor U14147 (N_14147,N_13812,N_13877);
nor U14148 (N_14148,N_14085,N_14087);
or U14149 (N_14149,N_13822,N_13908);
or U14150 (N_14150,N_13939,N_13999);
xor U14151 (N_14151,N_14076,N_13861);
xor U14152 (N_14152,N_13853,N_13909);
xnor U14153 (N_14153,N_14038,N_13832);
nor U14154 (N_14154,N_13868,N_13846);
nand U14155 (N_14155,N_14048,N_13803);
xnor U14156 (N_14156,N_14030,N_14046);
nand U14157 (N_14157,N_14061,N_13823);
xnor U14158 (N_14158,N_13991,N_13850);
xnor U14159 (N_14159,N_14021,N_14084);
xnor U14160 (N_14160,N_13948,N_13870);
or U14161 (N_14161,N_13977,N_13992);
nor U14162 (N_14162,N_14098,N_13928);
nand U14163 (N_14163,N_14075,N_14094);
or U14164 (N_14164,N_13859,N_14026);
and U14165 (N_14165,N_14012,N_13916);
or U14166 (N_14166,N_14065,N_14006);
nand U14167 (N_14167,N_13807,N_13970);
nand U14168 (N_14168,N_14028,N_13919);
and U14169 (N_14169,N_13813,N_13903);
nor U14170 (N_14170,N_13880,N_13829);
and U14171 (N_14171,N_13871,N_13902);
xnor U14172 (N_14172,N_13816,N_13990);
and U14173 (N_14173,N_13892,N_13897);
nor U14174 (N_14174,N_13976,N_13878);
and U14175 (N_14175,N_13840,N_13936);
or U14176 (N_14176,N_13896,N_14058);
nand U14177 (N_14177,N_13841,N_13895);
or U14178 (N_14178,N_13843,N_14088);
or U14179 (N_14179,N_14096,N_14040);
or U14180 (N_14180,N_14073,N_13849);
nand U14181 (N_14181,N_14080,N_13844);
or U14182 (N_14182,N_13915,N_14027);
nor U14183 (N_14183,N_13938,N_13876);
and U14184 (N_14184,N_13848,N_14082);
nor U14185 (N_14185,N_13893,N_14071);
or U14186 (N_14186,N_13957,N_13886);
and U14187 (N_14187,N_14086,N_13847);
and U14188 (N_14188,N_13937,N_13834);
nand U14189 (N_14189,N_13973,N_14022);
or U14190 (N_14190,N_13891,N_13971);
and U14191 (N_14191,N_14057,N_13907);
nor U14192 (N_14192,N_13956,N_13814);
nor U14193 (N_14193,N_14043,N_14081);
nand U14194 (N_14194,N_14093,N_13833);
xnor U14195 (N_14195,N_14089,N_13888);
xor U14196 (N_14196,N_14023,N_13913);
or U14197 (N_14197,N_13805,N_13969);
or U14198 (N_14198,N_13851,N_13987);
nand U14199 (N_14199,N_13930,N_14011);
or U14200 (N_14200,N_14024,N_13818);
nor U14201 (N_14201,N_13927,N_13954);
nand U14202 (N_14202,N_13949,N_13924);
nor U14203 (N_14203,N_14039,N_14015);
xnor U14204 (N_14204,N_14090,N_13882);
or U14205 (N_14205,N_13962,N_13830);
and U14206 (N_14206,N_13910,N_13998);
nand U14207 (N_14207,N_14033,N_13941);
and U14208 (N_14208,N_13952,N_13836);
and U14209 (N_14209,N_14029,N_14004);
nor U14210 (N_14210,N_13845,N_13874);
or U14211 (N_14211,N_13900,N_13819);
xnor U14212 (N_14212,N_13905,N_13828);
and U14213 (N_14213,N_13906,N_13989);
or U14214 (N_14214,N_13920,N_13953);
or U14215 (N_14215,N_13898,N_13935);
xnor U14216 (N_14216,N_14047,N_13944);
xor U14217 (N_14217,N_13804,N_13964);
xnor U14218 (N_14218,N_13960,N_13826);
nand U14219 (N_14219,N_13984,N_14074);
xor U14220 (N_14220,N_13993,N_14017);
nor U14221 (N_14221,N_14001,N_14032);
xor U14222 (N_14222,N_14064,N_13947);
and U14223 (N_14223,N_13806,N_13887);
or U14224 (N_14224,N_14092,N_13929);
and U14225 (N_14225,N_13867,N_13855);
xnor U14226 (N_14226,N_14003,N_13979);
xor U14227 (N_14227,N_14044,N_13860);
nor U14228 (N_14228,N_13940,N_14016);
and U14229 (N_14229,N_14099,N_13894);
and U14230 (N_14230,N_13820,N_13811);
nor U14231 (N_14231,N_13914,N_13921);
and U14232 (N_14232,N_14025,N_13911);
and U14233 (N_14233,N_13825,N_14041);
or U14234 (N_14234,N_14066,N_14097);
xnor U14235 (N_14235,N_14060,N_13963);
nand U14236 (N_14236,N_13865,N_13994);
xnor U14237 (N_14237,N_13821,N_13959);
or U14238 (N_14238,N_13864,N_14008);
nand U14239 (N_14239,N_13827,N_13802);
nor U14240 (N_14240,N_13817,N_13852);
and U14241 (N_14241,N_13837,N_13965);
or U14242 (N_14242,N_13815,N_13931);
and U14243 (N_14243,N_13951,N_13943);
nand U14244 (N_14244,N_14051,N_14018);
nor U14245 (N_14245,N_14072,N_14054);
nand U14246 (N_14246,N_13858,N_14069);
or U14247 (N_14247,N_14052,N_13985);
nand U14248 (N_14248,N_13863,N_13996);
nand U14249 (N_14249,N_13835,N_13933);
xnor U14250 (N_14250,N_13937,N_13836);
nand U14251 (N_14251,N_14042,N_14063);
nand U14252 (N_14252,N_14074,N_14050);
nand U14253 (N_14253,N_13881,N_14033);
nor U14254 (N_14254,N_13814,N_14038);
nor U14255 (N_14255,N_13808,N_13821);
nand U14256 (N_14256,N_13911,N_14066);
nor U14257 (N_14257,N_13953,N_13972);
nor U14258 (N_14258,N_13927,N_13812);
and U14259 (N_14259,N_13834,N_14072);
xor U14260 (N_14260,N_13866,N_14095);
and U14261 (N_14261,N_13878,N_14030);
and U14262 (N_14262,N_13912,N_13921);
xnor U14263 (N_14263,N_13854,N_13914);
and U14264 (N_14264,N_14081,N_14059);
and U14265 (N_14265,N_14001,N_14096);
nor U14266 (N_14266,N_13879,N_13891);
and U14267 (N_14267,N_13818,N_13870);
nor U14268 (N_14268,N_13997,N_14082);
nand U14269 (N_14269,N_13981,N_14044);
nor U14270 (N_14270,N_13981,N_13854);
nor U14271 (N_14271,N_13808,N_14078);
nand U14272 (N_14272,N_13843,N_13858);
or U14273 (N_14273,N_14012,N_13921);
nor U14274 (N_14274,N_13807,N_13883);
xnor U14275 (N_14275,N_13846,N_13956);
nand U14276 (N_14276,N_13903,N_13983);
and U14277 (N_14277,N_14071,N_14031);
nor U14278 (N_14278,N_13930,N_14053);
nor U14279 (N_14279,N_14014,N_13938);
nand U14280 (N_14280,N_13949,N_13953);
nand U14281 (N_14281,N_13901,N_13903);
or U14282 (N_14282,N_13845,N_14062);
or U14283 (N_14283,N_13884,N_14013);
and U14284 (N_14284,N_13875,N_14029);
and U14285 (N_14285,N_14092,N_13885);
nand U14286 (N_14286,N_14090,N_13825);
xor U14287 (N_14287,N_13843,N_13937);
xor U14288 (N_14288,N_13954,N_13978);
nor U14289 (N_14289,N_13814,N_14022);
nand U14290 (N_14290,N_13980,N_14018);
or U14291 (N_14291,N_14003,N_14065);
nand U14292 (N_14292,N_13826,N_14023);
nor U14293 (N_14293,N_14026,N_13862);
and U14294 (N_14294,N_14017,N_13906);
nor U14295 (N_14295,N_13838,N_14057);
nand U14296 (N_14296,N_14000,N_13954);
nor U14297 (N_14297,N_13985,N_13869);
nor U14298 (N_14298,N_13982,N_14047);
or U14299 (N_14299,N_14098,N_13902);
xor U14300 (N_14300,N_13950,N_13822);
and U14301 (N_14301,N_13912,N_13819);
nor U14302 (N_14302,N_13819,N_13836);
nor U14303 (N_14303,N_13939,N_13904);
xnor U14304 (N_14304,N_14076,N_14001);
or U14305 (N_14305,N_13879,N_14036);
nand U14306 (N_14306,N_13822,N_14017);
nor U14307 (N_14307,N_14013,N_13879);
nand U14308 (N_14308,N_13962,N_14019);
nor U14309 (N_14309,N_13945,N_13967);
or U14310 (N_14310,N_14093,N_13884);
or U14311 (N_14311,N_13974,N_13927);
xor U14312 (N_14312,N_14018,N_13999);
and U14313 (N_14313,N_14013,N_13845);
nor U14314 (N_14314,N_14067,N_13836);
xnor U14315 (N_14315,N_13905,N_13875);
xor U14316 (N_14316,N_13827,N_14065);
xnor U14317 (N_14317,N_13940,N_13825);
or U14318 (N_14318,N_13986,N_13885);
nor U14319 (N_14319,N_13863,N_13972);
and U14320 (N_14320,N_13989,N_14091);
nand U14321 (N_14321,N_14015,N_14029);
or U14322 (N_14322,N_13958,N_13950);
nand U14323 (N_14323,N_14046,N_13952);
and U14324 (N_14324,N_13982,N_13957);
or U14325 (N_14325,N_14030,N_13994);
xor U14326 (N_14326,N_14063,N_13880);
nor U14327 (N_14327,N_14092,N_13984);
nand U14328 (N_14328,N_14052,N_14096);
xor U14329 (N_14329,N_14055,N_14089);
nand U14330 (N_14330,N_13985,N_13862);
or U14331 (N_14331,N_14009,N_14075);
or U14332 (N_14332,N_13828,N_14044);
nor U14333 (N_14333,N_14079,N_14016);
nand U14334 (N_14334,N_13987,N_13852);
and U14335 (N_14335,N_14029,N_14031);
or U14336 (N_14336,N_14099,N_13838);
nand U14337 (N_14337,N_13867,N_13979);
nor U14338 (N_14338,N_14058,N_13942);
and U14339 (N_14339,N_13940,N_13842);
xnor U14340 (N_14340,N_14057,N_13953);
nor U14341 (N_14341,N_14037,N_13812);
nor U14342 (N_14342,N_13829,N_13883);
and U14343 (N_14343,N_13938,N_13899);
or U14344 (N_14344,N_13975,N_14007);
and U14345 (N_14345,N_13941,N_14086);
nand U14346 (N_14346,N_13987,N_13917);
nand U14347 (N_14347,N_13960,N_14043);
nand U14348 (N_14348,N_13902,N_14080);
xor U14349 (N_14349,N_13978,N_14000);
or U14350 (N_14350,N_14029,N_13955);
nor U14351 (N_14351,N_14026,N_13879);
and U14352 (N_14352,N_13886,N_13870);
nor U14353 (N_14353,N_13873,N_13803);
xnor U14354 (N_14354,N_13875,N_13944);
nand U14355 (N_14355,N_14010,N_14035);
nor U14356 (N_14356,N_14090,N_14029);
nand U14357 (N_14357,N_13871,N_13908);
and U14358 (N_14358,N_14014,N_13835);
or U14359 (N_14359,N_14087,N_13854);
nand U14360 (N_14360,N_14086,N_14077);
or U14361 (N_14361,N_13944,N_13806);
or U14362 (N_14362,N_13969,N_14094);
and U14363 (N_14363,N_14078,N_13806);
or U14364 (N_14364,N_14024,N_14091);
nand U14365 (N_14365,N_13917,N_13915);
or U14366 (N_14366,N_14087,N_13993);
and U14367 (N_14367,N_13917,N_13802);
nor U14368 (N_14368,N_13853,N_13881);
xor U14369 (N_14369,N_14094,N_14028);
nand U14370 (N_14370,N_14074,N_13950);
nand U14371 (N_14371,N_14014,N_13874);
or U14372 (N_14372,N_14097,N_13988);
xnor U14373 (N_14373,N_13941,N_13943);
nor U14374 (N_14374,N_14061,N_14084);
xnor U14375 (N_14375,N_13814,N_13982);
or U14376 (N_14376,N_13892,N_13871);
or U14377 (N_14377,N_13980,N_14074);
nand U14378 (N_14378,N_13906,N_14053);
and U14379 (N_14379,N_13857,N_13979);
and U14380 (N_14380,N_13962,N_13994);
or U14381 (N_14381,N_13815,N_13902);
nor U14382 (N_14382,N_14083,N_13893);
or U14383 (N_14383,N_14040,N_13907);
nor U14384 (N_14384,N_13880,N_13965);
xnor U14385 (N_14385,N_14069,N_14035);
xor U14386 (N_14386,N_13985,N_14028);
and U14387 (N_14387,N_13998,N_13914);
xor U14388 (N_14388,N_13854,N_13802);
nand U14389 (N_14389,N_13827,N_14066);
or U14390 (N_14390,N_13824,N_14092);
xor U14391 (N_14391,N_13901,N_14095);
nand U14392 (N_14392,N_13983,N_13907);
nand U14393 (N_14393,N_14071,N_13900);
xnor U14394 (N_14394,N_13814,N_13842);
nor U14395 (N_14395,N_13955,N_13984);
and U14396 (N_14396,N_14001,N_14074);
xnor U14397 (N_14397,N_13823,N_13979);
and U14398 (N_14398,N_13890,N_14030);
xor U14399 (N_14399,N_13814,N_13927);
nand U14400 (N_14400,N_14351,N_14294);
or U14401 (N_14401,N_14196,N_14356);
nand U14402 (N_14402,N_14397,N_14172);
nand U14403 (N_14403,N_14287,N_14216);
nor U14404 (N_14404,N_14158,N_14233);
and U14405 (N_14405,N_14240,N_14342);
nand U14406 (N_14406,N_14178,N_14286);
or U14407 (N_14407,N_14338,N_14210);
nand U14408 (N_14408,N_14268,N_14219);
and U14409 (N_14409,N_14252,N_14269);
and U14410 (N_14410,N_14247,N_14398);
nand U14411 (N_14411,N_14163,N_14116);
or U14412 (N_14412,N_14176,N_14171);
and U14413 (N_14413,N_14130,N_14293);
and U14414 (N_14414,N_14204,N_14224);
or U14415 (N_14415,N_14315,N_14109);
and U14416 (N_14416,N_14226,N_14237);
nand U14417 (N_14417,N_14359,N_14142);
and U14418 (N_14418,N_14190,N_14396);
xnor U14419 (N_14419,N_14319,N_14152);
nand U14420 (N_14420,N_14117,N_14144);
or U14421 (N_14421,N_14156,N_14201);
xnor U14422 (N_14422,N_14112,N_14312);
nor U14423 (N_14423,N_14120,N_14376);
nor U14424 (N_14424,N_14197,N_14255);
nor U14425 (N_14425,N_14275,N_14105);
or U14426 (N_14426,N_14303,N_14284);
nor U14427 (N_14427,N_14245,N_14289);
or U14428 (N_14428,N_14298,N_14336);
nor U14429 (N_14429,N_14122,N_14343);
xnor U14430 (N_14430,N_14367,N_14347);
nor U14431 (N_14431,N_14132,N_14332);
nand U14432 (N_14432,N_14324,N_14357);
or U14433 (N_14433,N_14148,N_14164);
or U14434 (N_14434,N_14346,N_14159);
and U14435 (N_14435,N_14341,N_14259);
and U14436 (N_14436,N_14111,N_14177);
nand U14437 (N_14437,N_14127,N_14136);
nor U14438 (N_14438,N_14299,N_14153);
xor U14439 (N_14439,N_14349,N_14189);
and U14440 (N_14440,N_14100,N_14350);
nand U14441 (N_14441,N_14313,N_14211);
nand U14442 (N_14442,N_14358,N_14166);
or U14443 (N_14443,N_14390,N_14339);
and U14444 (N_14444,N_14234,N_14364);
nor U14445 (N_14445,N_14184,N_14369);
nor U14446 (N_14446,N_14180,N_14282);
and U14447 (N_14447,N_14121,N_14183);
and U14448 (N_14448,N_14150,N_14311);
or U14449 (N_14449,N_14328,N_14126);
nand U14450 (N_14450,N_14119,N_14370);
nand U14451 (N_14451,N_14129,N_14212);
and U14452 (N_14452,N_14232,N_14308);
xnor U14453 (N_14453,N_14124,N_14361);
nand U14454 (N_14454,N_14273,N_14188);
and U14455 (N_14455,N_14271,N_14227);
nand U14456 (N_14456,N_14193,N_14187);
xor U14457 (N_14457,N_14387,N_14320);
and U14458 (N_14458,N_14221,N_14123);
nand U14459 (N_14459,N_14242,N_14223);
nand U14460 (N_14460,N_14160,N_14202);
or U14461 (N_14461,N_14246,N_14145);
xor U14462 (N_14462,N_14200,N_14258);
nor U14463 (N_14463,N_14326,N_14215);
or U14464 (N_14464,N_14229,N_14264);
xor U14465 (N_14465,N_14385,N_14309);
or U14466 (N_14466,N_14118,N_14251);
nand U14467 (N_14467,N_14292,N_14222);
nand U14468 (N_14468,N_14399,N_14261);
xnor U14469 (N_14469,N_14337,N_14296);
or U14470 (N_14470,N_14191,N_14388);
and U14471 (N_14471,N_14182,N_14174);
xnor U14472 (N_14472,N_14321,N_14128);
xor U14473 (N_14473,N_14248,N_14263);
nor U14474 (N_14474,N_14137,N_14161);
xor U14475 (N_14475,N_14114,N_14225);
or U14476 (N_14476,N_14348,N_14244);
xnor U14477 (N_14477,N_14394,N_14194);
or U14478 (N_14478,N_14318,N_14301);
and U14479 (N_14479,N_14362,N_14214);
nor U14480 (N_14480,N_14300,N_14250);
nor U14481 (N_14481,N_14218,N_14169);
and U14482 (N_14482,N_14181,N_14382);
and U14483 (N_14483,N_14203,N_14213);
nor U14484 (N_14484,N_14295,N_14154);
nor U14485 (N_14485,N_14220,N_14325);
or U14486 (N_14486,N_14393,N_14149);
nor U14487 (N_14487,N_14254,N_14360);
nand U14488 (N_14488,N_14272,N_14143);
nor U14489 (N_14489,N_14344,N_14283);
nor U14490 (N_14490,N_14340,N_14107);
or U14491 (N_14491,N_14354,N_14297);
xnor U14492 (N_14492,N_14131,N_14374);
or U14493 (N_14493,N_14125,N_14353);
or U14494 (N_14494,N_14199,N_14377);
and U14495 (N_14495,N_14322,N_14316);
or U14496 (N_14496,N_14334,N_14277);
xor U14497 (N_14497,N_14155,N_14290);
or U14498 (N_14498,N_14115,N_14106);
xor U14499 (N_14499,N_14345,N_14291);
nor U14500 (N_14500,N_14278,N_14375);
and U14501 (N_14501,N_14256,N_14192);
nor U14502 (N_14502,N_14262,N_14175);
nand U14503 (N_14503,N_14238,N_14355);
and U14504 (N_14504,N_14389,N_14392);
or U14505 (N_14505,N_14228,N_14134);
xor U14506 (N_14506,N_14281,N_14102);
nor U14507 (N_14507,N_14205,N_14386);
and U14508 (N_14508,N_14267,N_14280);
xnor U14509 (N_14509,N_14366,N_14276);
nand U14510 (N_14510,N_14260,N_14103);
and U14511 (N_14511,N_14288,N_14162);
or U14512 (N_14512,N_14179,N_14147);
nand U14513 (N_14513,N_14373,N_14383);
nand U14514 (N_14514,N_14380,N_14140);
or U14515 (N_14515,N_14323,N_14352);
and U14516 (N_14516,N_14395,N_14139);
nand U14517 (N_14517,N_14306,N_14329);
nor U14518 (N_14518,N_14141,N_14327);
xnor U14519 (N_14519,N_14113,N_14241);
nor U14520 (N_14520,N_14151,N_14257);
nor U14521 (N_14521,N_14372,N_14249);
nor U14522 (N_14522,N_14330,N_14208);
and U14523 (N_14523,N_14170,N_14379);
or U14524 (N_14524,N_14133,N_14335);
and U14525 (N_14525,N_14206,N_14381);
xnor U14526 (N_14526,N_14253,N_14239);
xnor U14527 (N_14527,N_14173,N_14371);
xnor U14528 (N_14528,N_14365,N_14231);
nand U14529 (N_14529,N_14270,N_14138);
or U14530 (N_14530,N_14368,N_14285);
nand U14531 (N_14531,N_14135,N_14331);
xor U14532 (N_14532,N_14217,N_14266);
and U14533 (N_14533,N_14108,N_14186);
xnor U14534 (N_14534,N_14101,N_14146);
nand U14535 (N_14535,N_14236,N_14384);
nand U14536 (N_14536,N_14167,N_14310);
nor U14537 (N_14537,N_14378,N_14307);
or U14538 (N_14538,N_14104,N_14302);
or U14539 (N_14539,N_14209,N_14157);
nand U14540 (N_14540,N_14165,N_14305);
nor U14541 (N_14541,N_14391,N_14304);
nand U14542 (N_14542,N_14243,N_14274);
nor U14543 (N_14543,N_14195,N_14230);
nor U14544 (N_14544,N_14279,N_14185);
or U14545 (N_14545,N_14235,N_14314);
or U14546 (N_14546,N_14363,N_14198);
or U14547 (N_14547,N_14207,N_14265);
and U14548 (N_14548,N_14333,N_14317);
and U14549 (N_14549,N_14110,N_14168);
or U14550 (N_14550,N_14228,N_14243);
and U14551 (N_14551,N_14288,N_14289);
nor U14552 (N_14552,N_14370,N_14392);
or U14553 (N_14553,N_14381,N_14120);
nand U14554 (N_14554,N_14367,N_14329);
and U14555 (N_14555,N_14109,N_14193);
nand U14556 (N_14556,N_14281,N_14217);
nand U14557 (N_14557,N_14148,N_14182);
and U14558 (N_14558,N_14372,N_14383);
or U14559 (N_14559,N_14144,N_14308);
nand U14560 (N_14560,N_14179,N_14126);
and U14561 (N_14561,N_14321,N_14122);
and U14562 (N_14562,N_14332,N_14165);
nand U14563 (N_14563,N_14197,N_14389);
or U14564 (N_14564,N_14348,N_14267);
or U14565 (N_14565,N_14143,N_14399);
xor U14566 (N_14566,N_14227,N_14222);
nand U14567 (N_14567,N_14114,N_14246);
xor U14568 (N_14568,N_14392,N_14227);
or U14569 (N_14569,N_14272,N_14298);
or U14570 (N_14570,N_14235,N_14239);
xor U14571 (N_14571,N_14303,N_14348);
nor U14572 (N_14572,N_14345,N_14367);
and U14573 (N_14573,N_14107,N_14334);
or U14574 (N_14574,N_14163,N_14215);
or U14575 (N_14575,N_14388,N_14134);
nor U14576 (N_14576,N_14139,N_14207);
nand U14577 (N_14577,N_14151,N_14247);
or U14578 (N_14578,N_14295,N_14213);
and U14579 (N_14579,N_14139,N_14217);
xnor U14580 (N_14580,N_14371,N_14249);
and U14581 (N_14581,N_14270,N_14133);
nand U14582 (N_14582,N_14215,N_14181);
or U14583 (N_14583,N_14182,N_14124);
nand U14584 (N_14584,N_14133,N_14169);
nand U14585 (N_14585,N_14198,N_14395);
nor U14586 (N_14586,N_14230,N_14207);
nand U14587 (N_14587,N_14241,N_14383);
or U14588 (N_14588,N_14273,N_14379);
xnor U14589 (N_14589,N_14370,N_14207);
xnor U14590 (N_14590,N_14290,N_14378);
xnor U14591 (N_14591,N_14200,N_14320);
nor U14592 (N_14592,N_14396,N_14104);
xnor U14593 (N_14593,N_14366,N_14244);
nand U14594 (N_14594,N_14113,N_14121);
nand U14595 (N_14595,N_14168,N_14366);
and U14596 (N_14596,N_14132,N_14321);
nor U14597 (N_14597,N_14222,N_14106);
nand U14598 (N_14598,N_14373,N_14147);
nand U14599 (N_14599,N_14159,N_14146);
or U14600 (N_14600,N_14186,N_14192);
xnor U14601 (N_14601,N_14113,N_14348);
nor U14602 (N_14602,N_14177,N_14170);
nor U14603 (N_14603,N_14226,N_14201);
xnor U14604 (N_14604,N_14219,N_14223);
or U14605 (N_14605,N_14210,N_14369);
or U14606 (N_14606,N_14125,N_14241);
nor U14607 (N_14607,N_14188,N_14314);
xnor U14608 (N_14608,N_14170,N_14387);
and U14609 (N_14609,N_14377,N_14217);
nor U14610 (N_14610,N_14177,N_14160);
xor U14611 (N_14611,N_14194,N_14238);
nor U14612 (N_14612,N_14394,N_14296);
and U14613 (N_14613,N_14344,N_14119);
nor U14614 (N_14614,N_14362,N_14104);
nor U14615 (N_14615,N_14197,N_14109);
nor U14616 (N_14616,N_14237,N_14110);
xnor U14617 (N_14617,N_14227,N_14183);
xor U14618 (N_14618,N_14100,N_14140);
nand U14619 (N_14619,N_14355,N_14302);
xor U14620 (N_14620,N_14131,N_14327);
nor U14621 (N_14621,N_14125,N_14370);
nor U14622 (N_14622,N_14347,N_14300);
or U14623 (N_14623,N_14162,N_14115);
nand U14624 (N_14624,N_14170,N_14115);
xnor U14625 (N_14625,N_14359,N_14177);
and U14626 (N_14626,N_14210,N_14131);
nand U14627 (N_14627,N_14171,N_14223);
xor U14628 (N_14628,N_14383,N_14284);
and U14629 (N_14629,N_14363,N_14275);
nor U14630 (N_14630,N_14234,N_14317);
nor U14631 (N_14631,N_14315,N_14285);
xnor U14632 (N_14632,N_14389,N_14330);
xor U14633 (N_14633,N_14326,N_14124);
or U14634 (N_14634,N_14161,N_14217);
xnor U14635 (N_14635,N_14170,N_14131);
nand U14636 (N_14636,N_14398,N_14315);
xnor U14637 (N_14637,N_14339,N_14157);
xor U14638 (N_14638,N_14267,N_14354);
and U14639 (N_14639,N_14238,N_14362);
nand U14640 (N_14640,N_14167,N_14135);
nor U14641 (N_14641,N_14240,N_14216);
or U14642 (N_14642,N_14243,N_14371);
or U14643 (N_14643,N_14345,N_14196);
and U14644 (N_14644,N_14297,N_14185);
xor U14645 (N_14645,N_14104,N_14115);
or U14646 (N_14646,N_14216,N_14236);
nand U14647 (N_14647,N_14174,N_14351);
nor U14648 (N_14648,N_14260,N_14206);
xor U14649 (N_14649,N_14336,N_14207);
or U14650 (N_14650,N_14343,N_14215);
and U14651 (N_14651,N_14375,N_14370);
or U14652 (N_14652,N_14146,N_14207);
nand U14653 (N_14653,N_14277,N_14244);
nor U14654 (N_14654,N_14171,N_14278);
or U14655 (N_14655,N_14388,N_14210);
nand U14656 (N_14656,N_14308,N_14207);
or U14657 (N_14657,N_14240,N_14288);
xnor U14658 (N_14658,N_14146,N_14278);
or U14659 (N_14659,N_14363,N_14115);
or U14660 (N_14660,N_14235,N_14241);
xor U14661 (N_14661,N_14397,N_14226);
nor U14662 (N_14662,N_14136,N_14285);
or U14663 (N_14663,N_14361,N_14247);
nor U14664 (N_14664,N_14161,N_14116);
nand U14665 (N_14665,N_14154,N_14352);
nor U14666 (N_14666,N_14194,N_14323);
and U14667 (N_14667,N_14363,N_14226);
xor U14668 (N_14668,N_14224,N_14125);
and U14669 (N_14669,N_14132,N_14181);
nand U14670 (N_14670,N_14272,N_14151);
xnor U14671 (N_14671,N_14209,N_14399);
and U14672 (N_14672,N_14249,N_14233);
or U14673 (N_14673,N_14359,N_14377);
and U14674 (N_14674,N_14281,N_14104);
nor U14675 (N_14675,N_14287,N_14249);
or U14676 (N_14676,N_14347,N_14369);
nand U14677 (N_14677,N_14299,N_14300);
xor U14678 (N_14678,N_14154,N_14132);
nand U14679 (N_14679,N_14286,N_14146);
nor U14680 (N_14680,N_14272,N_14293);
nor U14681 (N_14681,N_14193,N_14308);
nand U14682 (N_14682,N_14338,N_14103);
nor U14683 (N_14683,N_14185,N_14218);
nor U14684 (N_14684,N_14199,N_14343);
and U14685 (N_14685,N_14373,N_14227);
and U14686 (N_14686,N_14182,N_14147);
or U14687 (N_14687,N_14196,N_14280);
and U14688 (N_14688,N_14131,N_14182);
nor U14689 (N_14689,N_14214,N_14224);
xnor U14690 (N_14690,N_14105,N_14212);
or U14691 (N_14691,N_14106,N_14185);
and U14692 (N_14692,N_14196,N_14222);
xor U14693 (N_14693,N_14323,N_14387);
nand U14694 (N_14694,N_14150,N_14270);
nor U14695 (N_14695,N_14142,N_14156);
nand U14696 (N_14696,N_14136,N_14370);
and U14697 (N_14697,N_14156,N_14141);
nor U14698 (N_14698,N_14391,N_14206);
nor U14699 (N_14699,N_14157,N_14368);
or U14700 (N_14700,N_14501,N_14564);
xor U14701 (N_14701,N_14491,N_14676);
and U14702 (N_14702,N_14499,N_14656);
or U14703 (N_14703,N_14620,N_14563);
nor U14704 (N_14704,N_14553,N_14698);
nand U14705 (N_14705,N_14452,N_14612);
or U14706 (N_14706,N_14603,N_14632);
and U14707 (N_14707,N_14684,N_14496);
nor U14708 (N_14708,N_14506,N_14631);
xnor U14709 (N_14709,N_14677,N_14595);
and U14710 (N_14710,N_14586,N_14481);
nand U14711 (N_14711,N_14627,N_14574);
nor U14712 (N_14712,N_14653,N_14414);
nand U14713 (N_14713,N_14470,N_14458);
and U14714 (N_14714,N_14527,N_14615);
and U14715 (N_14715,N_14664,N_14607);
xnor U14716 (N_14716,N_14687,N_14512);
nor U14717 (N_14717,N_14541,N_14482);
xor U14718 (N_14718,N_14635,N_14445);
xnor U14719 (N_14719,N_14558,N_14579);
and U14720 (N_14720,N_14544,N_14652);
or U14721 (N_14721,N_14614,N_14469);
and U14722 (N_14722,N_14438,N_14565);
or U14723 (N_14723,N_14431,N_14619);
xnor U14724 (N_14724,N_14435,N_14427);
nor U14725 (N_14725,N_14401,N_14457);
xnor U14726 (N_14726,N_14673,N_14562);
xnor U14727 (N_14727,N_14412,N_14679);
nand U14728 (N_14728,N_14543,N_14492);
or U14729 (N_14729,N_14559,N_14411);
nor U14730 (N_14730,N_14505,N_14683);
nor U14731 (N_14731,N_14573,N_14460);
and U14732 (N_14732,N_14616,N_14450);
nand U14733 (N_14733,N_14568,N_14517);
nor U14734 (N_14734,N_14473,N_14474);
xnor U14735 (N_14735,N_14675,N_14650);
nand U14736 (N_14736,N_14613,N_14464);
xor U14737 (N_14737,N_14655,N_14525);
nand U14738 (N_14738,N_14649,N_14548);
xnor U14739 (N_14739,N_14608,N_14488);
nand U14740 (N_14740,N_14549,N_14534);
xnor U14741 (N_14741,N_14526,N_14425);
or U14742 (N_14742,N_14540,N_14671);
or U14743 (N_14743,N_14493,N_14536);
and U14744 (N_14744,N_14467,N_14640);
nand U14745 (N_14745,N_14530,N_14639);
nand U14746 (N_14746,N_14476,N_14442);
nor U14747 (N_14747,N_14682,N_14692);
and U14748 (N_14748,N_14528,N_14518);
nand U14749 (N_14749,N_14509,N_14602);
and U14750 (N_14750,N_14599,N_14666);
and U14751 (N_14751,N_14490,N_14532);
xor U14752 (N_14752,N_14628,N_14513);
or U14753 (N_14753,N_14459,N_14629);
xor U14754 (N_14754,N_14555,N_14456);
nor U14755 (N_14755,N_14550,N_14537);
xor U14756 (N_14756,N_14584,N_14441);
or U14757 (N_14757,N_14522,N_14663);
or U14758 (N_14758,N_14471,N_14487);
nand U14759 (N_14759,N_14669,N_14417);
or U14760 (N_14760,N_14606,N_14577);
and U14761 (N_14761,N_14500,N_14668);
xnor U14762 (N_14762,N_14510,N_14508);
xor U14763 (N_14763,N_14626,N_14609);
xor U14764 (N_14764,N_14623,N_14693);
xor U14765 (N_14765,N_14685,N_14524);
xnor U14766 (N_14766,N_14611,N_14430);
xor U14767 (N_14767,N_14497,N_14633);
xnor U14768 (N_14768,N_14697,N_14580);
nand U14769 (N_14769,N_14659,N_14423);
xnor U14770 (N_14770,N_14409,N_14691);
or U14771 (N_14771,N_14651,N_14521);
and U14772 (N_14772,N_14600,N_14572);
nor U14773 (N_14773,N_14503,N_14604);
xnor U14774 (N_14774,N_14403,N_14408);
or U14775 (N_14775,N_14433,N_14437);
nand U14776 (N_14776,N_14432,N_14566);
or U14777 (N_14777,N_14489,N_14554);
and U14778 (N_14778,N_14420,N_14453);
and U14779 (N_14779,N_14516,N_14617);
and U14780 (N_14780,N_14535,N_14475);
or U14781 (N_14781,N_14618,N_14542);
or U14782 (N_14782,N_14581,N_14598);
xnor U14783 (N_14783,N_14443,N_14406);
nand U14784 (N_14784,N_14688,N_14462);
xor U14785 (N_14785,N_14557,N_14434);
nand U14786 (N_14786,N_14419,N_14696);
xnor U14787 (N_14787,N_14647,N_14502);
nor U14788 (N_14788,N_14576,N_14660);
nand U14789 (N_14789,N_14680,N_14416);
or U14790 (N_14790,N_14404,N_14661);
or U14791 (N_14791,N_14690,N_14674);
or U14792 (N_14792,N_14422,N_14531);
xor U14793 (N_14793,N_14480,N_14477);
nor U14794 (N_14794,N_14556,N_14465);
xor U14795 (N_14795,N_14429,N_14498);
xor U14796 (N_14796,N_14587,N_14644);
and U14797 (N_14797,N_14630,N_14446);
nand U14798 (N_14798,N_14514,N_14689);
xor U14799 (N_14799,N_14461,N_14519);
nor U14800 (N_14800,N_14421,N_14410);
or U14801 (N_14801,N_14494,N_14699);
or U14802 (N_14802,N_14643,N_14415);
or U14803 (N_14803,N_14484,N_14538);
or U14804 (N_14804,N_14436,N_14529);
and U14805 (N_14805,N_14625,N_14463);
nand U14806 (N_14806,N_14523,N_14657);
xnor U14807 (N_14807,N_14455,N_14520);
and U14808 (N_14808,N_14428,N_14585);
nand U14809 (N_14809,N_14575,N_14636);
nor U14810 (N_14810,N_14624,N_14546);
xor U14811 (N_14811,N_14597,N_14400);
nor U14812 (N_14812,N_14515,N_14426);
and U14813 (N_14813,N_14567,N_14439);
nor U14814 (N_14814,N_14582,N_14686);
nand U14815 (N_14815,N_14472,N_14670);
nor U14816 (N_14816,N_14665,N_14592);
nor U14817 (N_14817,N_14589,N_14444);
xor U14818 (N_14818,N_14466,N_14694);
xor U14819 (N_14819,N_14681,N_14507);
nor U14820 (N_14820,N_14583,N_14662);
and U14821 (N_14821,N_14539,N_14596);
or U14822 (N_14822,N_14561,N_14407);
xnor U14823 (N_14823,N_14601,N_14610);
xnor U14824 (N_14824,N_14571,N_14638);
nor U14825 (N_14825,N_14552,N_14578);
nor U14826 (N_14826,N_14448,N_14413);
or U14827 (N_14827,N_14641,N_14551);
nor U14828 (N_14828,N_14504,N_14593);
and U14829 (N_14829,N_14695,N_14547);
and U14830 (N_14830,N_14495,N_14440);
xnor U14831 (N_14831,N_14590,N_14658);
xor U14832 (N_14832,N_14560,N_14468);
or U14833 (N_14833,N_14454,N_14621);
or U14834 (N_14834,N_14634,N_14591);
nor U14835 (N_14835,N_14451,N_14605);
or U14836 (N_14836,N_14479,N_14672);
nand U14837 (N_14837,N_14402,N_14646);
and U14838 (N_14838,N_14570,N_14424);
xnor U14839 (N_14839,N_14486,N_14645);
nor U14840 (N_14840,N_14447,N_14405);
xnor U14841 (N_14841,N_14637,N_14485);
and U14842 (N_14842,N_14622,N_14667);
or U14843 (N_14843,N_14545,N_14533);
and U14844 (N_14844,N_14588,N_14642);
nor U14845 (N_14845,N_14449,N_14678);
xnor U14846 (N_14846,N_14511,N_14418);
or U14847 (N_14847,N_14654,N_14569);
and U14848 (N_14848,N_14483,N_14478);
or U14849 (N_14849,N_14648,N_14594);
xnor U14850 (N_14850,N_14625,N_14599);
or U14851 (N_14851,N_14407,N_14696);
or U14852 (N_14852,N_14423,N_14550);
nor U14853 (N_14853,N_14606,N_14576);
or U14854 (N_14854,N_14678,N_14693);
nor U14855 (N_14855,N_14642,N_14696);
or U14856 (N_14856,N_14653,N_14636);
nor U14857 (N_14857,N_14687,N_14696);
and U14858 (N_14858,N_14694,N_14607);
nor U14859 (N_14859,N_14521,N_14699);
or U14860 (N_14860,N_14674,N_14410);
or U14861 (N_14861,N_14659,N_14586);
or U14862 (N_14862,N_14479,N_14441);
and U14863 (N_14863,N_14576,N_14691);
or U14864 (N_14864,N_14533,N_14486);
and U14865 (N_14865,N_14574,N_14561);
or U14866 (N_14866,N_14625,N_14533);
xor U14867 (N_14867,N_14663,N_14656);
or U14868 (N_14868,N_14629,N_14662);
nor U14869 (N_14869,N_14452,N_14445);
or U14870 (N_14870,N_14617,N_14559);
and U14871 (N_14871,N_14447,N_14459);
and U14872 (N_14872,N_14542,N_14540);
and U14873 (N_14873,N_14576,N_14541);
xor U14874 (N_14874,N_14436,N_14522);
nor U14875 (N_14875,N_14461,N_14433);
and U14876 (N_14876,N_14586,N_14401);
xor U14877 (N_14877,N_14639,N_14602);
nand U14878 (N_14878,N_14465,N_14615);
and U14879 (N_14879,N_14646,N_14435);
xor U14880 (N_14880,N_14423,N_14507);
nor U14881 (N_14881,N_14437,N_14563);
or U14882 (N_14882,N_14674,N_14449);
nor U14883 (N_14883,N_14566,N_14400);
nand U14884 (N_14884,N_14596,N_14476);
xor U14885 (N_14885,N_14622,N_14639);
nand U14886 (N_14886,N_14408,N_14582);
nand U14887 (N_14887,N_14512,N_14432);
nor U14888 (N_14888,N_14653,N_14489);
xnor U14889 (N_14889,N_14625,N_14600);
nor U14890 (N_14890,N_14612,N_14630);
and U14891 (N_14891,N_14426,N_14453);
nor U14892 (N_14892,N_14635,N_14409);
nand U14893 (N_14893,N_14680,N_14474);
nor U14894 (N_14894,N_14519,N_14612);
nor U14895 (N_14895,N_14566,N_14689);
nor U14896 (N_14896,N_14676,N_14525);
nand U14897 (N_14897,N_14646,N_14541);
xor U14898 (N_14898,N_14676,N_14457);
nor U14899 (N_14899,N_14514,N_14541);
nand U14900 (N_14900,N_14525,N_14621);
xor U14901 (N_14901,N_14451,N_14650);
xor U14902 (N_14902,N_14489,N_14565);
nor U14903 (N_14903,N_14691,N_14686);
and U14904 (N_14904,N_14446,N_14409);
or U14905 (N_14905,N_14425,N_14459);
nand U14906 (N_14906,N_14573,N_14574);
nor U14907 (N_14907,N_14483,N_14692);
and U14908 (N_14908,N_14551,N_14438);
xor U14909 (N_14909,N_14401,N_14669);
and U14910 (N_14910,N_14668,N_14612);
or U14911 (N_14911,N_14472,N_14620);
xnor U14912 (N_14912,N_14588,N_14638);
and U14913 (N_14913,N_14699,N_14420);
nand U14914 (N_14914,N_14656,N_14483);
nand U14915 (N_14915,N_14452,N_14427);
nand U14916 (N_14916,N_14611,N_14532);
and U14917 (N_14917,N_14419,N_14635);
nor U14918 (N_14918,N_14508,N_14580);
nand U14919 (N_14919,N_14613,N_14588);
or U14920 (N_14920,N_14457,N_14535);
or U14921 (N_14921,N_14494,N_14594);
or U14922 (N_14922,N_14649,N_14659);
or U14923 (N_14923,N_14406,N_14622);
nand U14924 (N_14924,N_14466,N_14523);
or U14925 (N_14925,N_14645,N_14571);
or U14926 (N_14926,N_14467,N_14517);
nor U14927 (N_14927,N_14650,N_14512);
and U14928 (N_14928,N_14595,N_14404);
and U14929 (N_14929,N_14656,N_14581);
or U14930 (N_14930,N_14400,N_14598);
nand U14931 (N_14931,N_14476,N_14480);
and U14932 (N_14932,N_14592,N_14485);
xnor U14933 (N_14933,N_14542,N_14415);
or U14934 (N_14934,N_14512,N_14670);
and U14935 (N_14935,N_14602,N_14456);
and U14936 (N_14936,N_14510,N_14496);
nor U14937 (N_14937,N_14428,N_14432);
and U14938 (N_14938,N_14549,N_14686);
or U14939 (N_14939,N_14588,N_14489);
and U14940 (N_14940,N_14442,N_14574);
nand U14941 (N_14941,N_14489,N_14486);
xor U14942 (N_14942,N_14463,N_14427);
nor U14943 (N_14943,N_14650,N_14464);
nand U14944 (N_14944,N_14600,N_14583);
nand U14945 (N_14945,N_14609,N_14455);
nand U14946 (N_14946,N_14601,N_14547);
or U14947 (N_14947,N_14620,N_14635);
or U14948 (N_14948,N_14407,N_14629);
nand U14949 (N_14949,N_14570,N_14457);
xnor U14950 (N_14950,N_14660,N_14532);
nand U14951 (N_14951,N_14650,N_14672);
and U14952 (N_14952,N_14438,N_14667);
xor U14953 (N_14953,N_14440,N_14505);
xor U14954 (N_14954,N_14547,N_14548);
xor U14955 (N_14955,N_14638,N_14468);
and U14956 (N_14956,N_14660,N_14464);
nor U14957 (N_14957,N_14528,N_14647);
or U14958 (N_14958,N_14441,N_14495);
or U14959 (N_14959,N_14408,N_14531);
or U14960 (N_14960,N_14637,N_14634);
nor U14961 (N_14961,N_14524,N_14665);
nor U14962 (N_14962,N_14637,N_14603);
nor U14963 (N_14963,N_14638,N_14486);
xor U14964 (N_14964,N_14635,N_14444);
and U14965 (N_14965,N_14433,N_14434);
xor U14966 (N_14966,N_14454,N_14569);
or U14967 (N_14967,N_14455,N_14521);
and U14968 (N_14968,N_14617,N_14571);
and U14969 (N_14969,N_14463,N_14499);
nand U14970 (N_14970,N_14651,N_14560);
and U14971 (N_14971,N_14498,N_14490);
or U14972 (N_14972,N_14446,N_14416);
xnor U14973 (N_14973,N_14495,N_14403);
and U14974 (N_14974,N_14654,N_14606);
xor U14975 (N_14975,N_14668,N_14660);
or U14976 (N_14976,N_14621,N_14683);
xnor U14977 (N_14977,N_14479,N_14631);
xnor U14978 (N_14978,N_14487,N_14502);
nand U14979 (N_14979,N_14650,N_14578);
xor U14980 (N_14980,N_14489,N_14595);
or U14981 (N_14981,N_14650,N_14667);
nand U14982 (N_14982,N_14478,N_14623);
or U14983 (N_14983,N_14406,N_14459);
xor U14984 (N_14984,N_14667,N_14553);
xnor U14985 (N_14985,N_14611,N_14428);
or U14986 (N_14986,N_14604,N_14400);
or U14987 (N_14987,N_14548,N_14567);
xnor U14988 (N_14988,N_14448,N_14415);
xor U14989 (N_14989,N_14515,N_14574);
nand U14990 (N_14990,N_14622,N_14551);
xor U14991 (N_14991,N_14519,N_14628);
nand U14992 (N_14992,N_14534,N_14541);
or U14993 (N_14993,N_14531,N_14692);
nand U14994 (N_14994,N_14413,N_14531);
and U14995 (N_14995,N_14603,N_14494);
nor U14996 (N_14996,N_14413,N_14544);
or U14997 (N_14997,N_14605,N_14588);
nor U14998 (N_14998,N_14418,N_14655);
nand U14999 (N_14999,N_14553,N_14427);
xnor U15000 (N_15000,N_14978,N_14796);
nor U15001 (N_15001,N_14757,N_14774);
nor U15002 (N_15002,N_14760,N_14961);
nand U15003 (N_15003,N_14967,N_14939);
or U15004 (N_15004,N_14711,N_14972);
and U15005 (N_15005,N_14914,N_14903);
nor U15006 (N_15006,N_14884,N_14783);
nand U15007 (N_15007,N_14859,N_14845);
nand U15008 (N_15008,N_14919,N_14714);
xor U15009 (N_15009,N_14964,N_14854);
and U15010 (N_15010,N_14894,N_14981);
or U15011 (N_15011,N_14720,N_14813);
nor U15012 (N_15012,N_14990,N_14723);
and U15013 (N_15013,N_14997,N_14901);
xnor U15014 (N_15014,N_14940,N_14878);
nor U15015 (N_15015,N_14945,N_14984);
or U15016 (N_15016,N_14860,N_14891);
or U15017 (N_15017,N_14730,N_14863);
xnor U15018 (N_15018,N_14971,N_14921);
nand U15019 (N_15019,N_14965,N_14942);
or U15020 (N_15020,N_14920,N_14795);
or U15021 (N_15021,N_14758,N_14794);
and U15022 (N_15022,N_14946,N_14886);
xnor U15023 (N_15023,N_14855,N_14804);
nor U15024 (N_15024,N_14974,N_14800);
nor U15025 (N_15025,N_14721,N_14750);
or U15026 (N_15026,N_14725,N_14709);
and U15027 (N_15027,N_14824,N_14814);
and U15028 (N_15028,N_14954,N_14772);
and U15029 (N_15029,N_14833,N_14789);
and U15030 (N_15030,N_14858,N_14742);
nor U15031 (N_15031,N_14775,N_14768);
nand U15032 (N_15032,N_14846,N_14717);
nand U15033 (N_15033,N_14927,N_14707);
and U15034 (N_15034,N_14861,N_14900);
nand U15035 (N_15035,N_14989,N_14994);
or U15036 (N_15036,N_14787,N_14827);
nor U15037 (N_15037,N_14744,N_14767);
and U15038 (N_15038,N_14749,N_14870);
nor U15039 (N_15039,N_14985,N_14890);
nor U15040 (N_15040,N_14713,N_14839);
nor U15041 (N_15041,N_14732,N_14881);
nand U15042 (N_15042,N_14752,N_14712);
and U15043 (N_15043,N_14933,N_14841);
nand U15044 (N_15044,N_14733,N_14851);
or U15045 (N_15045,N_14948,N_14931);
nand U15046 (N_15046,N_14778,N_14710);
or U15047 (N_15047,N_14703,N_14977);
or U15048 (N_15048,N_14829,N_14923);
or U15049 (N_15049,N_14777,N_14843);
or U15050 (N_15050,N_14850,N_14876);
nand U15051 (N_15051,N_14797,N_14748);
or U15052 (N_15052,N_14791,N_14719);
nand U15053 (N_15053,N_14957,N_14810);
xnor U15054 (N_15054,N_14943,N_14837);
nor U15055 (N_15055,N_14806,N_14947);
xor U15056 (N_15056,N_14716,N_14792);
nand U15057 (N_15057,N_14998,N_14992);
xnor U15058 (N_15058,N_14706,N_14782);
xor U15059 (N_15059,N_14738,N_14916);
xor U15060 (N_15060,N_14722,N_14746);
or U15061 (N_15061,N_14727,N_14838);
and U15062 (N_15062,N_14816,N_14770);
and U15063 (N_15063,N_14702,N_14786);
nand U15064 (N_15064,N_14831,N_14802);
nand U15065 (N_15065,N_14852,N_14999);
and U15066 (N_15066,N_14963,N_14905);
or U15067 (N_15067,N_14924,N_14734);
xor U15068 (N_15068,N_14736,N_14879);
or U15069 (N_15069,N_14949,N_14812);
nor U15070 (N_15070,N_14938,N_14729);
nand U15071 (N_15071,N_14877,N_14960);
and U15072 (N_15072,N_14743,N_14823);
nand U15073 (N_15073,N_14873,N_14980);
nand U15074 (N_15074,N_14906,N_14762);
or U15075 (N_15075,N_14780,N_14962);
nor U15076 (N_15076,N_14737,N_14883);
and U15077 (N_15077,N_14895,N_14987);
and U15078 (N_15078,N_14842,N_14844);
and U15079 (N_15079,N_14897,N_14889);
xnor U15080 (N_15080,N_14917,N_14968);
or U15081 (N_15081,N_14887,N_14740);
xnor U15082 (N_15082,N_14807,N_14821);
nand U15083 (N_15083,N_14896,N_14773);
and U15084 (N_15084,N_14867,N_14937);
xor U15085 (N_15085,N_14898,N_14769);
or U15086 (N_15086,N_14708,N_14956);
nor U15087 (N_15087,N_14996,N_14975);
and U15088 (N_15088,N_14761,N_14818);
nand U15089 (N_15089,N_14988,N_14907);
and U15090 (N_15090,N_14893,N_14882);
or U15091 (N_15091,N_14902,N_14934);
and U15092 (N_15092,N_14857,N_14763);
xor U15093 (N_15093,N_14941,N_14790);
nand U15094 (N_15094,N_14853,N_14741);
or U15095 (N_15095,N_14771,N_14728);
nor U15096 (N_15096,N_14995,N_14701);
nand U15097 (N_15097,N_14929,N_14830);
nor U15098 (N_15098,N_14776,N_14825);
xor U15099 (N_15099,N_14826,N_14815);
and U15100 (N_15100,N_14820,N_14908);
and U15101 (N_15101,N_14745,N_14718);
xnor U15102 (N_15102,N_14869,N_14910);
or U15103 (N_15103,N_14866,N_14784);
or U15104 (N_15104,N_14847,N_14819);
or U15105 (N_15105,N_14849,N_14788);
and U15106 (N_15106,N_14950,N_14928);
nor U15107 (N_15107,N_14836,N_14817);
nor U15108 (N_15108,N_14918,N_14872);
or U15109 (N_15109,N_14724,N_14922);
nor U15110 (N_15110,N_14756,N_14739);
nor U15111 (N_15111,N_14912,N_14805);
nor U15112 (N_15112,N_14944,N_14705);
nand U15113 (N_15113,N_14700,N_14735);
and U15114 (N_15114,N_14835,N_14856);
xor U15115 (N_15115,N_14899,N_14798);
nand U15116 (N_15116,N_14726,N_14754);
nor U15117 (N_15117,N_14865,N_14911);
nand U15118 (N_15118,N_14885,N_14888);
and U15119 (N_15119,N_14880,N_14765);
nand U15120 (N_15120,N_14973,N_14753);
nand U15121 (N_15121,N_14755,N_14970);
nand U15122 (N_15122,N_14785,N_14966);
nand U15123 (N_15123,N_14874,N_14986);
or U15124 (N_15124,N_14932,N_14982);
xor U15125 (N_15125,N_14811,N_14759);
and U15126 (N_15126,N_14864,N_14715);
or U15127 (N_15127,N_14801,N_14822);
xnor U15128 (N_15128,N_14840,N_14828);
or U15129 (N_15129,N_14935,N_14834);
or U15130 (N_15130,N_14868,N_14904);
or U15131 (N_15131,N_14976,N_14930);
or U15132 (N_15132,N_14871,N_14991);
nand U15133 (N_15133,N_14799,N_14993);
or U15134 (N_15134,N_14793,N_14731);
xor U15135 (N_15135,N_14747,N_14958);
nor U15136 (N_15136,N_14779,N_14925);
or U15137 (N_15137,N_14926,N_14909);
or U15138 (N_15138,N_14862,N_14832);
and U15139 (N_15139,N_14766,N_14951);
nor U15140 (N_15140,N_14875,N_14781);
nor U15141 (N_15141,N_14803,N_14969);
and U15142 (N_15142,N_14848,N_14764);
or U15143 (N_15143,N_14913,N_14704);
nand U15144 (N_15144,N_14751,N_14953);
xnor U15145 (N_15145,N_14979,N_14955);
xnor U15146 (N_15146,N_14809,N_14915);
and U15147 (N_15147,N_14892,N_14936);
nand U15148 (N_15148,N_14808,N_14959);
nand U15149 (N_15149,N_14983,N_14952);
nor U15150 (N_15150,N_14730,N_14707);
xnor U15151 (N_15151,N_14851,N_14832);
xor U15152 (N_15152,N_14840,N_14726);
nand U15153 (N_15153,N_14870,N_14835);
or U15154 (N_15154,N_14933,N_14758);
xnor U15155 (N_15155,N_14878,N_14931);
nor U15156 (N_15156,N_14872,N_14738);
xnor U15157 (N_15157,N_14748,N_14882);
nor U15158 (N_15158,N_14928,N_14942);
nor U15159 (N_15159,N_14951,N_14744);
or U15160 (N_15160,N_14966,N_14914);
nand U15161 (N_15161,N_14834,N_14773);
xnor U15162 (N_15162,N_14850,N_14784);
nor U15163 (N_15163,N_14804,N_14880);
nor U15164 (N_15164,N_14825,N_14887);
xor U15165 (N_15165,N_14878,N_14972);
nand U15166 (N_15166,N_14825,N_14924);
nor U15167 (N_15167,N_14833,N_14759);
xnor U15168 (N_15168,N_14926,N_14779);
or U15169 (N_15169,N_14715,N_14904);
or U15170 (N_15170,N_14771,N_14835);
and U15171 (N_15171,N_14967,N_14943);
or U15172 (N_15172,N_14911,N_14701);
and U15173 (N_15173,N_14718,N_14774);
xnor U15174 (N_15174,N_14799,N_14704);
xor U15175 (N_15175,N_14934,N_14781);
nor U15176 (N_15176,N_14909,N_14815);
and U15177 (N_15177,N_14722,N_14805);
and U15178 (N_15178,N_14869,N_14962);
nor U15179 (N_15179,N_14974,N_14787);
nand U15180 (N_15180,N_14919,N_14916);
xor U15181 (N_15181,N_14858,N_14777);
nor U15182 (N_15182,N_14879,N_14726);
nand U15183 (N_15183,N_14722,N_14758);
and U15184 (N_15184,N_14810,N_14825);
and U15185 (N_15185,N_14860,N_14867);
nand U15186 (N_15186,N_14793,N_14996);
and U15187 (N_15187,N_14856,N_14875);
nor U15188 (N_15188,N_14780,N_14950);
nand U15189 (N_15189,N_14846,N_14993);
or U15190 (N_15190,N_14908,N_14702);
and U15191 (N_15191,N_14728,N_14881);
and U15192 (N_15192,N_14968,N_14843);
nand U15193 (N_15193,N_14929,N_14815);
and U15194 (N_15194,N_14741,N_14987);
or U15195 (N_15195,N_14917,N_14978);
xor U15196 (N_15196,N_14958,N_14780);
nor U15197 (N_15197,N_14831,N_14855);
nand U15198 (N_15198,N_14826,N_14773);
and U15199 (N_15199,N_14760,N_14894);
or U15200 (N_15200,N_14810,N_14968);
nand U15201 (N_15201,N_14999,N_14939);
xor U15202 (N_15202,N_14767,N_14926);
nand U15203 (N_15203,N_14930,N_14724);
or U15204 (N_15204,N_14725,N_14723);
and U15205 (N_15205,N_14798,N_14705);
nand U15206 (N_15206,N_14975,N_14799);
nor U15207 (N_15207,N_14741,N_14826);
nand U15208 (N_15208,N_14991,N_14881);
nor U15209 (N_15209,N_14768,N_14895);
nor U15210 (N_15210,N_14741,N_14701);
nand U15211 (N_15211,N_14722,N_14711);
xor U15212 (N_15212,N_14922,N_14853);
nor U15213 (N_15213,N_14871,N_14994);
or U15214 (N_15214,N_14953,N_14902);
nand U15215 (N_15215,N_14827,N_14991);
and U15216 (N_15216,N_14847,N_14867);
and U15217 (N_15217,N_14872,N_14991);
xnor U15218 (N_15218,N_14880,N_14864);
or U15219 (N_15219,N_14810,N_14871);
nand U15220 (N_15220,N_14728,N_14801);
nand U15221 (N_15221,N_14722,N_14840);
nor U15222 (N_15222,N_14719,N_14881);
and U15223 (N_15223,N_14741,N_14828);
or U15224 (N_15224,N_14774,N_14841);
nand U15225 (N_15225,N_14806,N_14996);
nor U15226 (N_15226,N_14700,N_14788);
xnor U15227 (N_15227,N_14737,N_14824);
nor U15228 (N_15228,N_14707,N_14760);
or U15229 (N_15229,N_14737,N_14788);
and U15230 (N_15230,N_14821,N_14767);
nand U15231 (N_15231,N_14702,N_14931);
nand U15232 (N_15232,N_14912,N_14753);
nand U15233 (N_15233,N_14903,N_14896);
or U15234 (N_15234,N_14761,N_14779);
xor U15235 (N_15235,N_14838,N_14809);
nand U15236 (N_15236,N_14766,N_14812);
nand U15237 (N_15237,N_14742,N_14836);
or U15238 (N_15238,N_14933,N_14824);
nor U15239 (N_15239,N_14783,N_14832);
nand U15240 (N_15240,N_14794,N_14842);
nand U15241 (N_15241,N_14761,N_14923);
nor U15242 (N_15242,N_14806,N_14918);
nand U15243 (N_15243,N_14743,N_14908);
or U15244 (N_15244,N_14978,N_14878);
and U15245 (N_15245,N_14734,N_14968);
nand U15246 (N_15246,N_14858,N_14814);
and U15247 (N_15247,N_14838,N_14915);
or U15248 (N_15248,N_14745,N_14972);
nand U15249 (N_15249,N_14820,N_14841);
or U15250 (N_15250,N_14865,N_14785);
or U15251 (N_15251,N_14778,N_14883);
and U15252 (N_15252,N_14815,N_14714);
or U15253 (N_15253,N_14704,N_14888);
or U15254 (N_15254,N_14886,N_14811);
and U15255 (N_15255,N_14779,N_14721);
and U15256 (N_15256,N_14794,N_14844);
nand U15257 (N_15257,N_14842,N_14886);
and U15258 (N_15258,N_14821,N_14931);
xor U15259 (N_15259,N_14987,N_14831);
xor U15260 (N_15260,N_14990,N_14800);
xnor U15261 (N_15261,N_14791,N_14937);
or U15262 (N_15262,N_14843,N_14976);
or U15263 (N_15263,N_14750,N_14745);
nand U15264 (N_15264,N_14886,N_14725);
nand U15265 (N_15265,N_14961,N_14853);
or U15266 (N_15266,N_14904,N_14755);
nor U15267 (N_15267,N_14718,N_14777);
or U15268 (N_15268,N_14919,N_14800);
nand U15269 (N_15269,N_14881,N_14856);
and U15270 (N_15270,N_14751,N_14888);
and U15271 (N_15271,N_14797,N_14911);
nand U15272 (N_15272,N_14754,N_14811);
nand U15273 (N_15273,N_14979,N_14789);
or U15274 (N_15274,N_14846,N_14719);
and U15275 (N_15275,N_14764,N_14773);
and U15276 (N_15276,N_14892,N_14924);
nor U15277 (N_15277,N_14795,N_14720);
nand U15278 (N_15278,N_14738,N_14942);
or U15279 (N_15279,N_14982,N_14899);
nor U15280 (N_15280,N_14822,N_14744);
xor U15281 (N_15281,N_14826,N_14963);
xnor U15282 (N_15282,N_14779,N_14942);
or U15283 (N_15283,N_14906,N_14857);
and U15284 (N_15284,N_14975,N_14752);
nand U15285 (N_15285,N_14864,N_14828);
or U15286 (N_15286,N_14716,N_14980);
nor U15287 (N_15287,N_14754,N_14815);
and U15288 (N_15288,N_14758,N_14889);
nor U15289 (N_15289,N_14818,N_14840);
and U15290 (N_15290,N_14912,N_14809);
nand U15291 (N_15291,N_14784,N_14852);
nand U15292 (N_15292,N_14728,N_14719);
xnor U15293 (N_15293,N_14994,N_14967);
and U15294 (N_15294,N_14803,N_14950);
xor U15295 (N_15295,N_14913,N_14887);
nor U15296 (N_15296,N_14872,N_14816);
nand U15297 (N_15297,N_14820,N_14828);
nand U15298 (N_15298,N_14897,N_14856);
xnor U15299 (N_15299,N_14909,N_14743);
nor U15300 (N_15300,N_15159,N_15104);
or U15301 (N_15301,N_15042,N_15208);
nand U15302 (N_15302,N_15010,N_15021);
or U15303 (N_15303,N_15262,N_15275);
xnor U15304 (N_15304,N_15024,N_15255);
xor U15305 (N_15305,N_15111,N_15153);
xor U15306 (N_15306,N_15271,N_15165);
or U15307 (N_15307,N_15047,N_15158);
nor U15308 (N_15308,N_15294,N_15059);
xor U15309 (N_15309,N_15265,N_15070);
or U15310 (N_15310,N_15261,N_15210);
or U15311 (N_15311,N_15121,N_15001);
xnor U15312 (N_15312,N_15013,N_15061);
nor U15313 (N_15313,N_15072,N_15202);
and U15314 (N_15314,N_15119,N_15172);
or U15315 (N_15315,N_15114,N_15205);
and U15316 (N_15316,N_15068,N_15009);
xor U15317 (N_15317,N_15243,N_15170);
xnor U15318 (N_15318,N_15297,N_15122);
or U15319 (N_15319,N_15178,N_15045);
nand U15320 (N_15320,N_15143,N_15272);
and U15321 (N_15321,N_15195,N_15293);
xnor U15322 (N_15322,N_15112,N_15081);
nor U15323 (N_15323,N_15270,N_15175);
nor U15324 (N_15324,N_15152,N_15179);
nor U15325 (N_15325,N_15100,N_15128);
xnor U15326 (N_15326,N_15204,N_15134);
xor U15327 (N_15327,N_15129,N_15237);
nor U15328 (N_15328,N_15177,N_15066);
nand U15329 (N_15329,N_15238,N_15180);
and U15330 (N_15330,N_15290,N_15133);
and U15331 (N_15331,N_15199,N_15196);
and U15332 (N_15332,N_15215,N_15228);
nand U15333 (N_15333,N_15156,N_15110);
or U15334 (N_15334,N_15011,N_15249);
nor U15335 (N_15335,N_15240,N_15281);
or U15336 (N_15336,N_15246,N_15039);
xnor U15337 (N_15337,N_15162,N_15226);
nor U15338 (N_15338,N_15169,N_15284);
xnor U15339 (N_15339,N_15218,N_15221);
or U15340 (N_15340,N_15233,N_15223);
and U15341 (N_15341,N_15142,N_15231);
and U15342 (N_15342,N_15025,N_15012);
xnor U15343 (N_15343,N_15147,N_15168);
xor U15344 (N_15344,N_15136,N_15023);
xnor U15345 (N_15345,N_15015,N_15279);
nand U15346 (N_15346,N_15028,N_15097);
nor U15347 (N_15347,N_15087,N_15299);
nor U15348 (N_15348,N_15101,N_15131);
or U15349 (N_15349,N_15161,N_15194);
nand U15350 (N_15350,N_15115,N_15092);
or U15351 (N_15351,N_15171,N_15258);
nand U15352 (N_15352,N_15190,N_15004);
xnor U15353 (N_15353,N_15099,N_15053);
nand U15354 (N_15354,N_15079,N_15086);
or U15355 (N_15355,N_15184,N_15005);
or U15356 (N_15356,N_15096,N_15257);
or U15357 (N_15357,N_15127,N_15252);
nor U15358 (N_15358,N_15049,N_15106);
and U15359 (N_15359,N_15135,N_15227);
xor U15360 (N_15360,N_15055,N_15295);
and U15361 (N_15361,N_15264,N_15230);
xor U15362 (N_15362,N_15076,N_15046);
or U15363 (N_15363,N_15080,N_15285);
nor U15364 (N_15364,N_15298,N_15244);
and U15365 (N_15365,N_15183,N_15085);
nand U15366 (N_15366,N_15187,N_15274);
or U15367 (N_15367,N_15051,N_15224);
nand U15368 (N_15368,N_15269,N_15071);
nand U15369 (N_15369,N_15222,N_15268);
xor U15370 (N_15370,N_15232,N_15213);
or U15371 (N_15371,N_15200,N_15229);
xnor U15372 (N_15372,N_15173,N_15182);
nand U15373 (N_15373,N_15007,N_15148);
xor U15374 (N_15374,N_15043,N_15266);
and U15375 (N_15375,N_15250,N_15094);
and U15376 (N_15376,N_15002,N_15186);
and U15377 (N_15377,N_15149,N_15283);
or U15378 (N_15378,N_15235,N_15019);
or U15379 (N_15379,N_15286,N_15146);
nand U15380 (N_15380,N_15212,N_15123);
or U15381 (N_15381,N_15247,N_15069);
and U15382 (N_15382,N_15132,N_15256);
xnor U15383 (N_15383,N_15107,N_15103);
nand U15384 (N_15384,N_15054,N_15063);
xnor U15385 (N_15385,N_15277,N_15280);
and U15386 (N_15386,N_15098,N_15207);
nor U15387 (N_15387,N_15095,N_15031);
or U15388 (N_15388,N_15248,N_15181);
or U15389 (N_15389,N_15130,N_15044);
or U15390 (N_15390,N_15254,N_15203);
xnor U15391 (N_15391,N_15034,N_15120);
nand U15392 (N_15392,N_15078,N_15139);
xor U15393 (N_15393,N_15056,N_15263);
nand U15394 (N_15394,N_15201,N_15260);
or U15395 (N_15395,N_15174,N_15189);
or U15396 (N_15396,N_15113,N_15057);
nand U15397 (N_15397,N_15155,N_15000);
or U15398 (N_15398,N_15060,N_15050);
and U15399 (N_15399,N_15220,N_15030);
or U15400 (N_15400,N_15282,N_15091);
or U15401 (N_15401,N_15058,N_15154);
nor U15402 (N_15402,N_15003,N_15029);
nor U15403 (N_15403,N_15150,N_15242);
or U15404 (N_15404,N_15141,N_15117);
and U15405 (N_15405,N_15188,N_15018);
nor U15406 (N_15406,N_15288,N_15273);
nand U15407 (N_15407,N_15077,N_15291);
and U15408 (N_15408,N_15105,N_15126);
or U15409 (N_15409,N_15234,N_15206);
and U15410 (N_15410,N_15214,N_15074);
and U15411 (N_15411,N_15016,N_15160);
and U15412 (N_15412,N_15287,N_15035);
xor U15413 (N_15413,N_15278,N_15245);
nand U15414 (N_15414,N_15089,N_15032);
or U15415 (N_15415,N_15289,N_15192);
nand U15416 (N_15416,N_15197,N_15062);
nand U15417 (N_15417,N_15027,N_15191);
nand U15418 (N_15418,N_15125,N_15108);
or U15419 (N_15419,N_15109,N_15006);
nand U15420 (N_15420,N_15041,N_15088);
and U15421 (N_15421,N_15137,N_15167);
nand U15422 (N_15422,N_15151,N_15073);
xnor U15423 (N_15423,N_15022,N_15083);
nor U15424 (N_15424,N_15211,N_15185);
or U15425 (N_15425,N_15033,N_15064);
nand U15426 (N_15426,N_15198,N_15038);
or U15427 (N_15427,N_15251,N_15140);
xor U15428 (N_15428,N_15048,N_15276);
nand U15429 (N_15429,N_15144,N_15163);
nor U15430 (N_15430,N_15267,N_15036);
xnor U15431 (N_15431,N_15216,N_15236);
nor U15432 (N_15432,N_15067,N_15219);
nor U15433 (N_15433,N_15116,N_15020);
xor U15434 (N_15434,N_15193,N_15292);
or U15435 (N_15435,N_15145,N_15017);
nand U15436 (N_15436,N_15093,N_15040);
nand U15437 (N_15437,N_15118,N_15075);
or U15438 (N_15438,N_15026,N_15138);
and U15439 (N_15439,N_15164,N_15239);
nor U15440 (N_15440,N_15102,N_15259);
nor U15441 (N_15441,N_15008,N_15090);
xnor U15442 (N_15442,N_15241,N_15166);
or U15443 (N_15443,N_15176,N_15296);
or U15444 (N_15444,N_15084,N_15253);
nand U15445 (N_15445,N_15157,N_15065);
and U15446 (N_15446,N_15014,N_15209);
and U15447 (N_15447,N_15225,N_15217);
or U15448 (N_15448,N_15124,N_15052);
xnor U15449 (N_15449,N_15037,N_15082);
nand U15450 (N_15450,N_15186,N_15140);
xnor U15451 (N_15451,N_15271,N_15298);
and U15452 (N_15452,N_15061,N_15166);
xnor U15453 (N_15453,N_15067,N_15185);
xnor U15454 (N_15454,N_15038,N_15204);
or U15455 (N_15455,N_15103,N_15040);
nand U15456 (N_15456,N_15102,N_15219);
nand U15457 (N_15457,N_15284,N_15187);
nand U15458 (N_15458,N_15175,N_15081);
xor U15459 (N_15459,N_15299,N_15195);
nand U15460 (N_15460,N_15246,N_15275);
xnor U15461 (N_15461,N_15238,N_15046);
xnor U15462 (N_15462,N_15050,N_15076);
xor U15463 (N_15463,N_15256,N_15025);
nand U15464 (N_15464,N_15230,N_15242);
and U15465 (N_15465,N_15281,N_15062);
nand U15466 (N_15466,N_15051,N_15024);
and U15467 (N_15467,N_15141,N_15070);
or U15468 (N_15468,N_15209,N_15069);
or U15469 (N_15469,N_15022,N_15288);
and U15470 (N_15470,N_15084,N_15121);
nor U15471 (N_15471,N_15247,N_15197);
nand U15472 (N_15472,N_15154,N_15172);
nand U15473 (N_15473,N_15120,N_15290);
and U15474 (N_15474,N_15256,N_15238);
or U15475 (N_15475,N_15096,N_15040);
and U15476 (N_15476,N_15273,N_15099);
nor U15477 (N_15477,N_15002,N_15142);
nor U15478 (N_15478,N_15123,N_15073);
or U15479 (N_15479,N_15030,N_15058);
xor U15480 (N_15480,N_15219,N_15132);
nor U15481 (N_15481,N_15020,N_15286);
xnor U15482 (N_15482,N_15070,N_15060);
or U15483 (N_15483,N_15245,N_15062);
xor U15484 (N_15484,N_15285,N_15066);
and U15485 (N_15485,N_15005,N_15189);
and U15486 (N_15486,N_15127,N_15044);
nand U15487 (N_15487,N_15271,N_15205);
or U15488 (N_15488,N_15240,N_15053);
or U15489 (N_15489,N_15224,N_15018);
and U15490 (N_15490,N_15086,N_15041);
and U15491 (N_15491,N_15022,N_15172);
xor U15492 (N_15492,N_15084,N_15235);
nor U15493 (N_15493,N_15083,N_15118);
xor U15494 (N_15494,N_15144,N_15056);
nand U15495 (N_15495,N_15005,N_15253);
xor U15496 (N_15496,N_15086,N_15280);
xnor U15497 (N_15497,N_15041,N_15171);
xnor U15498 (N_15498,N_15129,N_15096);
and U15499 (N_15499,N_15279,N_15240);
or U15500 (N_15500,N_15094,N_15153);
and U15501 (N_15501,N_15022,N_15294);
nor U15502 (N_15502,N_15176,N_15139);
xor U15503 (N_15503,N_15186,N_15249);
nor U15504 (N_15504,N_15222,N_15204);
or U15505 (N_15505,N_15203,N_15147);
and U15506 (N_15506,N_15189,N_15072);
or U15507 (N_15507,N_15209,N_15078);
or U15508 (N_15508,N_15138,N_15011);
and U15509 (N_15509,N_15242,N_15029);
xor U15510 (N_15510,N_15263,N_15282);
nor U15511 (N_15511,N_15211,N_15066);
nor U15512 (N_15512,N_15215,N_15051);
nand U15513 (N_15513,N_15106,N_15054);
nor U15514 (N_15514,N_15298,N_15290);
or U15515 (N_15515,N_15043,N_15282);
xor U15516 (N_15516,N_15240,N_15272);
nand U15517 (N_15517,N_15047,N_15102);
nand U15518 (N_15518,N_15054,N_15059);
nor U15519 (N_15519,N_15042,N_15204);
xor U15520 (N_15520,N_15041,N_15289);
xor U15521 (N_15521,N_15168,N_15037);
xor U15522 (N_15522,N_15232,N_15270);
xor U15523 (N_15523,N_15249,N_15234);
xor U15524 (N_15524,N_15011,N_15107);
and U15525 (N_15525,N_15106,N_15088);
and U15526 (N_15526,N_15007,N_15085);
xor U15527 (N_15527,N_15089,N_15148);
nand U15528 (N_15528,N_15197,N_15209);
nor U15529 (N_15529,N_15114,N_15080);
xnor U15530 (N_15530,N_15171,N_15137);
or U15531 (N_15531,N_15283,N_15213);
xor U15532 (N_15532,N_15015,N_15155);
nor U15533 (N_15533,N_15060,N_15097);
and U15534 (N_15534,N_15223,N_15145);
nand U15535 (N_15535,N_15170,N_15299);
nand U15536 (N_15536,N_15032,N_15118);
nor U15537 (N_15537,N_15098,N_15206);
nor U15538 (N_15538,N_15106,N_15251);
xnor U15539 (N_15539,N_15147,N_15103);
or U15540 (N_15540,N_15262,N_15022);
and U15541 (N_15541,N_15125,N_15268);
nand U15542 (N_15542,N_15044,N_15271);
or U15543 (N_15543,N_15127,N_15188);
or U15544 (N_15544,N_15264,N_15218);
or U15545 (N_15545,N_15146,N_15061);
and U15546 (N_15546,N_15271,N_15031);
and U15547 (N_15547,N_15139,N_15005);
nor U15548 (N_15548,N_15273,N_15211);
nor U15549 (N_15549,N_15151,N_15290);
or U15550 (N_15550,N_15017,N_15284);
nand U15551 (N_15551,N_15273,N_15029);
xor U15552 (N_15552,N_15109,N_15023);
xor U15553 (N_15553,N_15047,N_15120);
nor U15554 (N_15554,N_15021,N_15158);
xnor U15555 (N_15555,N_15084,N_15231);
or U15556 (N_15556,N_15071,N_15230);
and U15557 (N_15557,N_15284,N_15228);
nand U15558 (N_15558,N_15157,N_15032);
or U15559 (N_15559,N_15134,N_15241);
or U15560 (N_15560,N_15026,N_15031);
and U15561 (N_15561,N_15185,N_15212);
and U15562 (N_15562,N_15183,N_15087);
nor U15563 (N_15563,N_15018,N_15141);
or U15564 (N_15564,N_15121,N_15168);
nand U15565 (N_15565,N_15212,N_15016);
xnor U15566 (N_15566,N_15229,N_15268);
or U15567 (N_15567,N_15144,N_15001);
or U15568 (N_15568,N_15073,N_15260);
xor U15569 (N_15569,N_15200,N_15018);
and U15570 (N_15570,N_15049,N_15281);
xnor U15571 (N_15571,N_15108,N_15269);
nor U15572 (N_15572,N_15288,N_15286);
and U15573 (N_15573,N_15084,N_15029);
nand U15574 (N_15574,N_15157,N_15189);
nand U15575 (N_15575,N_15222,N_15255);
or U15576 (N_15576,N_15218,N_15204);
and U15577 (N_15577,N_15170,N_15079);
and U15578 (N_15578,N_15196,N_15183);
nand U15579 (N_15579,N_15076,N_15113);
or U15580 (N_15580,N_15128,N_15174);
and U15581 (N_15581,N_15243,N_15218);
or U15582 (N_15582,N_15058,N_15294);
or U15583 (N_15583,N_15230,N_15153);
and U15584 (N_15584,N_15209,N_15185);
and U15585 (N_15585,N_15007,N_15153);
nand U15586 (N_15586,N_15147,N_15166);
or U15587 (N_15587,N_15270,N_15220);
xnor U15588 (N_15588,N_15196,N_15288);
and U15589 (N_15589,N_15184,N_15074);
xnor U15590 (N_15590,N_15093,N_15205);
xnor U15591 (N_15591,N_15241,N_15032);
and U15592 (N_15592,N_15205,N_15291);
nand U15593 (N_15593,N_15218,N_15119);
and U15594 (N_15594,N_15113,N_15077);
or U15595 (N_15595,N_15249,N_15251);
and U15596 (N_15596,N_15251,N_15017);
nand U15597 (N_15597,N_15111,N_15049);
nor U15598 (N_15598,N_15293,N_15211);
and U15599 (N_15599,N_15003,N_15086);
and U15600 (N_15600,N_15505,N_15577);
and U15601 (N_15601,N_15550,N_15318);
nor U15602 (N_15602,N_15383,N_15503);
nand U15603 (N_15603,N_15467,N_15418);
xnor U15604 (N_15604,N_15320,N_15327);
xor U15605 (N_15605,N_15426,N_15410);
or U15606 (N_15606,N_15516,N_15317);
or U15607 (N_15607,N_15420,N_15463);
nor U15608 (N_15608,N_15399,N_15509);
xor U15609 (N_15609,N_15345,N_15543);
nor U15610 (N_15610,N_15485,N_15560);
nor U15611 (N_15611,N_15579,N_15433);
xnor U15612 (N_15612,N_15434,N_15329);
or U15613 (N_15613,N_15557,N_15519);
or U15614 (N_15614,N_15362,N_15357);
or U15615 (N_15615,N_15444,N_15595);
nand U15616 (N_15616,N_15382,N_15551);
nor U15617 (N_15617,N_15562,N_15436);
xnor U15618 (N_15618,N_15568,N_15451);
nand U15619 (N_15619,N_15561,N_15571);
nor U15620 (N_15620,N_15342,N_15337);
or U15621 (N_15621,N_15507,N_15376);
or U15622 (N_15622,N_15487,N_15529);
nand U15623 (N_15623,N_15498,N_15552);
or U15624 (N_15624,N_15502,N_15555);
nor U15625 (N_15625,N_15431,N_15581);
xor U15626 (N_15626,N_15428,N_15532);
and U15627 (N_15627,N_15578,N_15334);
and U15628 (N_15628,N_15300,N_15338);
xor U15629 (N_15629,N_15441,N_15398);
nand U15630 (N_15630,N_15378,N_15301);
xor U15631 (N_15631,N_15363,N_15512);
nand U15632 (N_15632,N_15305,N_15554);
or U15633 (N_15633,N_15586,N_15304);
or U15634 (N_15634,N_15477,N_15452);
xnor U15635 (N_15635,N_15306,N_15352);
nor U15636 (N_15636,N_15351,N_15440);
nor U15637 (N_15637,N_15397,N_15443);
or U15638 (N_15638,N_15567,N_15589);
nor U15639 (N_15639,N_15437,N_15439);
or U15640 (N_15640,N_15457,N_15384);
xor U15641 (N_15641,N_15423,N_15530);
nor U15642 (N_15642,N_15360,N_15447);
xnor U15643 (N_15643,N_15474,N_15573);
xnor U15644 (N_15644,N_15421,N_15330);
or U15645 (N_15645,N_15597,N_15387);
nand U15646 (N_15646,N_15558,N_15394);
and U15647 (N_15647,N_15566,N_15303);
xnor U15648 (N_15648,N_15564,N_15479);
nand U15649 (N_15649,N_15324,N_15525);
or U15650 (N_15650,N_15599,N_15489);
xor U15651 (N_15651,N_15582,N_15537);
and U15652 (N_15652,N_15535,N_15454);
xor U15653 (N_15653,N_15548,N_15596);
nor U15654 (N_15654,N_15417,N_15392);
and U15655 (N_15655,N_15598,N_15367);
nand U15656 (N_15656,N_15580,N_15432);
nor U15657 (N_15657,N_15464,N_15359);
nand U15658 (N_15658,N_15312,N_15326);
nor U15659 (N_15659,N_15335,N_15563);
xor U15660 (N_15660,N_15372,N_15478);
xnor U15661 (N_15661,N_15390,N_15511);
nor U15662 (N_15662,N_15336,N_15325);
xor U15663 (N_15663,N_15400,N_15381);
xor U15664 (N_15664,N_15349,N_15435);
and U15665 (N_15665,N_15361,N_15476);
or U15666 (N_15666,N_15339,N_15544);
or U15667 (N_15667,N_15526,N_15412);
or U15668 (N_15668,N_15499,N_15379);
xnor U15669 (N_15669,N_15486,N_15380);
nand U15670 (N_15670,N_15565,N_15373);
nand U15671 (N_15671,N_15471,N_15388);
and U15672 (N_15672,N_15425,N_15402);
nand U15673 (N_15673,N_15468,N_15522);
or U15674 (N_15674,N_15493,N_15510);
xnor U15675 (N_15675,N_15411,N_15587);
or U15676 (N_15676,N_15539,N_15308);
nand U15677 (N_15677,N_15442,N_15460);
nor U15678 (N_15678,N_15430,N_15403);
nor U15679 (N_15679,N_15371,N_15302);
or U15680 (N_15680,N_15496,N_15414);
or U15681 (N_15681,N_15538,N_15483);
and U15682 (N_15682,N_15356,N_15500);
and U15683 (N_15683,N_15574,N_15584);
and U15684 (N_15684,N_15350,N_15309);
nand U15685 (N_15685,N_15521,N_15540);
xor U15686 (N_15686,N_15527,N_15341);
or U15687 (N_15687,N_15575,N_15466);
and U15688 (N_15688,N_15514,N_15316);
xor U15689 (N_15689,N_15546,N_15310);
nor U15690 (N_15690,N_15368,N_15406);
and U15691 (N_15691,N_15408,N_15438);
nand U15692 (N_15692,N_15470,N_15307);
xor U15693 (N_15693,N_15409,N_15386);
nand U15694 (N_15694,N_15333,N_15506);
xnor U15695 (N_15695,N_15355,N_15491);
nor U15696 (N_15696,N_15413,N_15427);
xor U15697 (N_15697,N_15585,N_15559);
or U15698 (N_15698,N_15453,N_15482);
and U15699 (N_15699,N_15448,N_15570);
xor U15700 (N_15700,N_15343,N_15508);
nand U15701 (N_15701,N_15545,N_15315);
nand U15702 (N_15702,N_15473,N_15344);
xor U15703 (N_15703,N_15524,N_15340);
nand U15704 (N_15704,N_15370,N_15364);
and U15705 (N_15705,N_15484,N_15536);
and U15706 (N_15706,N_15407,N_15475);
nor U15707 (N_15707,N_15328,N_15501);
and U15708 (N_15708,N_15553,N_15576);
xnor U15709 (N_15709,N_15593,N_15462);
and U15710 (N_15710,N_15534,N_15523);
or U15711 (N_15711,N_15401,N_15405);
nor U15712 (N_15712,N_15445,N_15449);
or U15713 (N_15713,N_15323,N_15396);
xor U15714 (N_15714,N_15458,N_15450);
nor U15715 (N_15715,N_15313,N_15490);
xor U15716 (N_15716,N_15569,N_15549);
nor U15717 (N_15717,N_15369,N_15415);
and U15718 (N_15718,N_15377,N_15346);
and U15719 (N_15719,N_15347,N_15547);
xor U15720 (N_15720,N_15492,N_15533);
or U15721 (N_15721,N_15389,N_15469);
or U15722 (N_15722,N_15531,N_15354);
nand U15723 (N_15723,N_15416,N_15395);
nor U15724 (N_15724,N_15424,N_15375);
xor U15725 (N_15725,N_15495,N_15374);
or U15726 (N_15726,N_15517,N_15348);
xnor U15727 (N_15727,N_15455,N_15591);
xor U15728 (N_15728,N_15515,N_15385);
and U15729 (N_15729,N_15314,N_15332);
nor U15730 (N_15730,N_15542,N_15541);
or U15731 (N_15731,N_15365,N_15321);
nor U15732 (N_15732,N_15419,N_15461);
nor U15733 (N_15733,N_15528,N_15572);
nand U15734 (N_15734,N_15404,N_15422);
and U15735 (N_15735,N_15429,N_15472);
nand U15736 (N_15736,N_15592,N_15480);
nor U15737 (N_15737,N_15513,N_15504);
xnor U15738 (N_15738,N_15590,N_15594);
nor U15739 (N_15739,N_15358,N_15459);
or U15740 (N_15740,N_15556,N_15583);
and U15741 (N_15741,N_15520,N_15481);
or U15742 (N_15742,N_15588,N_15465);
or U15743 (N_15743,N_15391,N_15488);
xnor U15744 (N_15744,N_15319,N_15353);
nand U15745 (N_15745,N_15322,N_15331);
nor U15746 (N_15746,N_15518,N_15393);
nor U15747 (N_15747,N_15366,N_15311);
nand U15748 (N_15748,N_15456,N_15494);
xor U15749 (N_15749,N_15497,N_15446);
nand U15750 (N_15750,N_15365,N_15425);
or U15751 (N_15751,N_15401,N_15581);
nand U15752 (N_15752,N_15383,N_15409);
or U15753 (N_15753,N_15469,N_15382);
xor U15754 (N_15754,N_15352,N_15409);
and U15755 (N_15755,N_15566,N_15509);
and U15756 (N_15756,N_15489,N_15483);
xnor U15757 (N_15757,N_15385,N_15329);
nand U15758 (N_15758,N_15400,N_15597);
nand U15759 (N_15759,N_15469,N_15555);
and U15760 (N_15760,N_15337,N_15456);
and U15761 (N_15761,N_15359,N_15450);
or U15762 (N_15762,N_15484,N_15497);
xor U15763 (N_15763,N_15476,N_15581);
xor U15764 (N_15764,N_15503,N_15366);
and U15765 (N_15765,N_15579,N_15532);
nor U15766 (N_15766,N_15554,N_15536);
nor U15767 (N_15767,N_15506,N_15404);
nand U15768 (N_15768,N_15430,N_15342);
or U15769 (N_15769,N_15317,N_15302);
xor U15770 (N_15770,N_15370,N_15300);
or U15771 (N_15771,N_15443,N_15453);
or U15772 (N_15772,N_15581,N_15481);
nand U15773 (N_15773,N_15316,N_15501);
nor U15774 (N_15774,N_15407,N_15419);
and U15775 (N_15775,N_15377,N_15477);
and U15776 (N_15776,N_15332,N_15596);
nand U15777 (N_15777,N_15496,N_15592);
xor U15778 (N_15778,N_15570,N_15455);
xnor U15779 (N_15779,N_15477,N_15578);
nand U15780 (N_15780,N_15469,N_15328);
nor U15781 (N_15781,N_15476,N_15515);
xnor U15782 (N_15782,N_15597,N_15402);
nor U15783 (N_15783,N_15342,N_15550);
nand U15784 (N_15784,N_15548,N_15448);
nand U15785 (N_15785,N_15535,N_15384);
and U15786 (N_15786,N_15527,N_15363);
or U15787 (N_15787,N_15461,N_15381);
nor U15788 (N_15788,N_15411,N_15392);
and U15789 (N_15789,N_15430,N_15518);
or U15790 (N_15790,N_15597,N_15401);
nor U15791 (N_15791,N_15441,N_15498);
nor U15792 (N_15792,N_15417,N_15373);
and U15793 (N_15793,N_15541,N_15589);
or U15794 (N_15794,N_15396,N_15320);
nor U15795 (N_15795,N_15563,N_15366);
xor U15796 (N_15796,N_15353,N_15538);
nor U15797 (N_15797,N_15339,N_15300);
or U15798 (N_15798,N_15351,N_15487);
nand U15799 (N_15799,N_15564,N_15498);
nor U15800 (N_15800,N_15398,N_15461);
or U15801 (N_15801,N_15456,N_15305);
nand U15802 (N_15802,N_15561,N_15300);
and U15803 (N_15803,N_15487,N_15567);
nand U15804 (N_15804,N_15584,N_15336);
nand U15805 (N_15805,N_15365,N_15482);
and U15806 (N_15806,N_15341,N_15392);
xor U15807 (N_15807,N_15460,N_15547);
nand U15808 (N_15808,N_15425,N_15465);
or U15809 (N_15809,N_15467,N_15503);
and U15810 (N_15810,N_15503,N_15320);
xor U15811 (N_15811,N_15315,N_15399);
and U15812 (N_15812,N_15447,N_15484);
nand U15813 (N_15813,N_15361,N_15598);
nand U15814 (N_15814,N_15539,N_15570);
xnor U15815 (N_15815,N_15364,N_15359);
and U15816 (N_15816,N_15552,N_15492);
and U15817 (N_15817,N_15309,N_15593);
nand U15818 (N_15818,N_15505,N_15370);
or U15819 (N_15819,N_15383,N_15378);
or U15820 (N_15820,N_15545,N_15433);
or U15821 (N_15821,N_15366,N_15543);
nor U15822 (N_15822,N_15456,N_15325);
nor U15823 (N_15823,N_15541,N_15510);
xor U15824 (N_15824,N_15499,N_15562);
nand U15825 (N_15825,N_15557,N_15475);
xnor U15826 (N_15826,N_15330,N_15466);
xnor U15827 (N_15827,N_15412,N_15356);
or U15828 (N_15828,N_15524,N_15410);
or U15829 (N_15829,N_15404,N_15448);
nor U15830 (N_15830,N_15322,N_15509);
nand U15831 (N_15831,N_15325,N_15333);
or U15832 (N_15832,N_15528,N_15437);
nand U15833 (N_15833,N_15303,N_15534);
or U15834 (N_15834,N_15490,N_15465);
nand U15835 (N_15835,N_15596,N_15587);
nand U15836 (N_15836,N_15498,N_15573);
and U15837 (N_15837,N_15525,N_15379);
xnor U15838 (N_15838,N_15451,N_15564);
nand U15839 (N_15839,N_15330,N_15590);
nor U15840 (N_15840,N_15565,N_15462);
nand U15841 (N_15841,N_15434,N_15512);
nor U15842 (N_15842,N_15415,N_15472);
nor U15843 (N_15843,N_15593,N_15356);
or U15844 (N_15844,N_15431,N_15427);
nand U15845 (N_15845,N_15527,N_15445);
xor U15846 (N_15846,N_15428,N_15308);
xor U15847 (N_15847,N_15564,N_15446);
nand U15848 (N_15848,N_15466,N_15350);
or U15849 (N_15849,N_15329,N_15345);
nor U15850 (N_15850,N_15519,N_15414);
nor U15851 (N_15851,N_15572,N_15575);
or U15852 (N_15852,N_15539,N_15406);
xnor U15853 (N_15853,N_15521,N_15434);
nand U15854 (N_15854,N_15527,N_15344);
xnor U15855 (N_15855,N_15308,N_15337);
or U15856 (N_15856,N_15392,N_15400);
or U15857 (N_15857,N_15573,N_15585);
or U15858 (N_15858,N_15413,N_15355);
xnor U15859 (N_15859,N_15462,N_15380);
or U15860 (N_15860,N_15428,N_15479);
nor U15861 (N_15861,N_15387,N_15443);
xnor U15862 (N_15862,N_15353,N_15372);
xor U15863 (N_15863,N_15582,N_15511);
nor U15864 (N_15864,N_15442,N_15585);
or U15865 (N_15865,N_15500,N_15492);
xnor U15866 (N_15866,N_15464,N_15472);
nor U15867 (N_15867,N_15578,N_15419);
nor U15868 (N_15868,N_15432,N_15389);
xnor U15869 (N_15869,N_15595,N_15397);
nand U15870 (N_15870,N_15467,N_15431);
nor U15871 (N_15871,N_15371,N_15458);
nand U15872 (N_15872,N_15361,N_15438);
nor U15873 (N_15873,N_15453,N_15373);
nor U15874 (N_15874,N_15312,N_15354);
or U15875 (N_15875,N_15469,N_15326);
and U15876 (N_15876,N_15324,N_15467);
and U15877 (N_15877,N_15478,N_15355);
or U15878 (N_15878,N_15552,N_15345);
nor U15879 (N_15879,N_15442,N_15493);
nor U15880 (N_15880,N_15321,N_15547);
nand U15881 (N_15881,N_15388,N_15412);
nor U15882 (N_15882,N_15435,N_15571);
or U15883 (N_15883,N_15427,N_15419);
nor U15884 (N_15884,N_15457,N_15351);
xnor U15885 (N_15885,N_15535,N_15526);
nand U15886 (N_15886,N_15526,N_15347);
xnor U15887 (N_15887,N_15447,N_15488);
and U15888 (N_15888,N_15384,N_15450);
nor U15889 (N_15889,N_15551,N_15538);
nor U15890 (N_15890,N_15421,N_15349);
or U15891 (N_15891,N_15304,N_15569);
nand U15892 (N_15892,N_15592,N_15562);
or U15893 (N_15893,N_15529,N_15408);
nand U15894 (N_15894,N_15386,N_15358);
nor U15895 (N_15895,N_15542,N_15467);
or U15896 (N_15896,N_15518,N_15392);
nand U15897 (N_15897,N_15378,N_15564);
xnor U15898 (N_15898,N_15557,N_15553);
nor U15899 (N_15899,N_15449,N_15342);
or U15900 (N_15900,N_15822,N_15882);
xor U15901 (N_15901,N_15744,N_15793);
or U15902 (N_15902,N_15717,N_15879);
nor U15903 (N_15903,N_15656,N_15835);
or U15904 (N_15904,N_15718,N_15840);
nand U15905 (N_15905,N_15674,N_15629);
and U15906 (N_15906,N_15687,N_15620);
or U15907 (N_15907,N_15646,N_15821);
nand U15908 (N_15908,N_15626,N_15621);
nand U15909 (N_15909,N_15788,N_15731);
and U15910 (N_15910,N_15894,N_15673);
or U15911 (N_15911,N_15860,N_15809);
xnor U15912 (N_15912,N_15874,N_15801);
and U15913 (N_15913,N_15833,N_15769);
nor U15914 (N_15914,N_15751,N_15796);
xnor U15915 (N_15915,N_15741,N_15783);
and U15916 (N_15916,N_15750,N_15863);
or U15917 (N_15917,N_15649,N_15828);
or U15918 (N_15918,N_15755,N_15842);
nor U15919 (N_15919,N_15647,N_15701);
xnor U15920 (N_15920,N_15612,N_15864);
or U15921 (N_15921,N_15766,N_15634);
xnor U15922 (N_15922,N_15730,N_15618);
xnor U15923 (N_15923,N_15825,N_15876);
xor U15924 (N_15924,N_15797,N_15732);
nand U15925 (N_15925,N_15684,N_15816);
xor U15926 (N_15926,N_15676,N_15726);
nor U15927 (N_15927,N_15712,N_15688);
xnor U15928 (N_15928,N_15720,N_15625);
and U15929 (N_15929,N_15651,N_15811);
xnor U15930 (N_15930,N_15705,N_15770);
nor U15931 (N_15931,N_15680,N_15675);
xor U15932 (N_15932,N_15606,N_15703);
and U15933 (N_15933,N_15791,N_15645);
nand U15934 (N_15934,N_15633,N_15807);
xnor U15935 (N_15935,N_15891,N_15780);
nor U15936 (N_15936,N_15692,N_15658);
or U15937 (N_15937,N_15857,N_15848);
and U15938 (N_15938,N_15873,N_15771);
nor U15939 (N_15939,N_15608,N_15870);
and U15940 (N_15940,N_15686,N_15823);
xor U15941 (N_15941,N_15733,N_15839);
nor U15942 (N_15942,N_15767,N_15867);
nand U15943 (N_15943,N_15852,N_15679);
nor U15944 (N_15944,N_15641,N_15710);
or U15945 (N_15945,N_15762,N_15846);
nor U15946 (N_15946,N_15670,N_15868);
nor U15947 (N_15947,N_15704,N_15885);
nand U15948 (N_15948,N_15654,N_15697);
or U15949 (N_15949,N_15896,N_15856);
xnor U15950 (N_15950,N_15752,N_15764);
and U15951 (N_15951,N_15691,N_15756);
nor U15952 (N_15952,N_15624,N_15818);
nor U15953 (N_15953,N_15844,N_15812);
or U15954 (N_15954,N_15655,N_15820);
and U15955 (N_15955,N_15662,N_15849);
xor U15956 (N_15956,N_15808,N_15802);
nor U15957 (N_15957,N_15859,N_15630);
and U15958 (N_15958,N_15814,N_15806);
and U15959 (N_15959,N_15636,N_15895);
nor U15960 (N_15960,N_15681,N_15711);
and U15961 (N_15961,N_15660,N_15843);
or U15962 (N_15962,N_15619,N_15714);
nand U15963 (N_15963,N_15795,N_15798);
nor U15964 (N_15964,N_15616,N_15897);
and U15965 (N_15965,N_15878,N_15836);
xnor U15966 (N_15966,N_15683,N_15607);
xor U15967 (N_15967,N_15889,N_15761);
and U15968 (N_15968,N_15890,N_15749);
xnor U15969 (N_15969,N_15648,N_15785);
and U15970 (N_15970,N_15815,N_15622);
xnor U15971 (N_15971,N_15694,N_15871);
nand U15972 (N_15972,N_15700,N_15610);
xnor U15973 (N_15973,N_15774,N_15736);
nand U15974 (N_15974,N_15725,N_15777);
xor U15975 (N_15975,N_15810,N_15778);
nand U15976 (N_15976,N_15862,N_15790);
nand U15977 (N_15977,N_15743,N_15838);
or U15978 (N_15978,N_15775,N_15602);
nor U15979 (N_15979,N_15695,N_15643);
or U15980 (N_15980,N_15742,N_15600);
xor U15981 (N_15981,N_15824,N_15872);
xor U15982 (N_15982,N_15804,N_15841);
nand U15983 (N_15983,N_15851,N_15758);
nand U15984 (N_15984,N_15800,N_15668);
nand U15985 (N_15985,N_15779,N_15696);
and U15986 (N_15986,N_15690,N_15702);
nor U15987 (N_15987,N_15792,N_15665);
xor U15988 (N_15988,N_15786,N_15784);
and U15989 (N_15989,N_15826,N_15617);
or U15990 (N_15990,N_15830,N_15754);
nand U15991 (N_15991,N_15898,N_15604);
nand U15992 (N_15992,N_15671,N_15729);
or U15993 (N_15993,N_15854,N_15734);
nor U15994 (N_15994,N_15635,N_15613);
nand U15995 (N_15995,N_15776,N_15640);
and U15996 (N_15996,N_15739,N_15735);
and U15997 (N_15997,N_15603,N_15866);
nor U15998 (N_15998,N_15716,N_15677);
xor U15999 (N_15999,N_15713,N_15899);
nor U16000 (N_16000,N_15757,N_15638);
nand U16001 (N_16001,N_15781,N_15672);
xor U16002 (N_16002,N_15787,N_15637);
and U16003 (N_16003,N_15759,N_15650);
nor U16004 (N_16004,N_15853,N_15623);
and U16005 (N_16005,N_15737,N_15858);
and U16006 (N_16006,N_15642,N_15869);
and U16007 (N_16007,N_15829,N_15805);
nand U16008 (N_16008,N_15847,N_15760);
nor U16009 (N_16009,N_15601,N_15609);
nor U16010 (N_16010,N_15614,N_15819);
xor U16011 (N_16011,N_15765,N_15753);
xnor U16012 (N_16012,N_15855,N_15659);
and U16013 (N_16013,N_15667,N_15627);
nand U16014 (N_16014,N_15605,N_15831);
or U16015 (N_16015,N_15880,N_15693);
nor U16016 (N_16016,N_15768,N_15698);
nor U16017 (N_16017,N_15707,N_15763);
and U16018 (N_16018,N_15669,N_15794);
nor U16019 (N_16019,N_15631,N_15772);
or U16020 (N_16020,N_15682,N_15664);
xor U16021 (N_16021,N_15887,N_15813);
and U16022 (N_16022,N_15657,N_15745);
or U16023 (N_16023,N_15803,N_15721);
xnor U16024 (N_16024,N_15834,N_15748);
and U16025 (N_16025,N_15773,N_15850);
nand U16026 (N_16026,N_15661,N_15865);
and U16027 (N_16027,N_15837,N_15747);
xor U16028 (N_16028,N_15789,N_15881);
and U16029 (N_16029,N_15875,N_15722);
nor U16030 (N_16030,N_15827,N_15832);
xor U16031 (N_16031,N_15861,N_15877);
nor U16032 (N_16032,N_15615,N_15706);
xor U16033 (N_16033,N_15740,N_15893);
and U16034 (N_16034,N_15799,N_15845);
or U16035 (N_16035,N_15782,N_15892);
nor U16036 (N_16036,N_15746,N_15663);
and U16037 (N_16037,N_15724,N_15709);
and U16038 (N_16038,N_15817,N_15728);
or U16039 (N_16039,N_15653,N_15639);
and U16040 (N_16040,N_15719,N_15644);
nor U16041 (N_16041,N_15886,N_15628);
and U16042 (N_16042,N_15708,N_15883);
nor U16043 (N_16043,N_15689,N_15884);
or U16044 (N_16044,N_15678,N_15888);
and U16045 (N_16045,N_15666,N_15632);
and U16046 (N_16046,N_15723,N_15738);
and U16047 (N_16047,N_15727,N_15699);
and U16048 (N_16048,N_15715,N_15652);
or U16049 (N_16049,N_15611,N_15685);
nand U16050 (N_16050,N_15756,N_15847);
nand U16051 (N_16051,N_15693,N_15718);
and U16052 (N_16052,N_15659,N_15766);
or U16053 (N_16053,N_15799,N_15843);
or U16054 (N_16054,N_15673,N_15885);
or U16055 (N_16055,N_15802,N_15842);
nand U16056 (N_16056,N_15713,N_15610);
nand U16057 (N_16057,N_15667,N_15858);
nor U16058 (N_16058,N_15767,N_15893);
or U16059 (N_16059,N_15745,N_15604);
xnor U16060 (N_16060,N_15898,N_15737);
or U16061 (N_16061,N_15654,N_15690);
nand U16062 (N_16062,N_15669,N_15731);
nor U16063 (N_16063,N_15663,N_15648);
or U16064 (N_16064,N_15653,N_15802);
nor U16065 (N_16065,N_15704,N_15810);
or U16066 (N_16066,N_15895,N_15772);
nor U16067 (N_16067,N_15838,N_15721);
or U16068 (N_16068,N_15623,N_15688);
and U16069 (N_16069,N_15803,N_15696);
xnor U16070 (N_16070,N_15753,N_15818);
or U16071 (N_16071,N_15824,N_15749);
xor U16072 (N_16072,N_15734,N_15657);
or U16073 (N_16073,N_15788,N_15730);
or U16074 (N_16074,N_15708,N_15866);
nor U16075 (N_16075,N_15706,N_15720);
nand U16076 (N_16076,N_15714,N_15697);
or U16077 (N_16077,N_15639,N_15728);
nor U16078 (N_16078,N_15759,N_15853);
or U16079 (N_16079,N_15768,N_15872);
nor U16080 (N_16080,N_15767,N_15894);
and U16081 (N_16081,N_15728,N_15758);
nor U16082 (N_16082,N_15703,N_15741);
nor U16083 (N_16083,N_15806,N_15828);
nor U16084 (N_16084,N_15696,N_15850);
and U16085 (N_16085,N_15765,N_15790);
nor U16086 (N_16086,N_15734,N_15767);
and U16087 (N_16087,N_15721,N_15695);
or U16088 (N_16088,N_15751,N_15696);
and U16089 (N_16089,N_15643,N_15698);
nand U16090 (N_16090,N_15709,N_15754);
or U16091 (N_16091,N_15788,N_15858);
nand U16092 (N_16092,N_15644,N_15703);
and U16093 (N_16093,N_15783,N_15845);
nand U16094 (N_16094,N_15804,N_15616);
or U16095 (N_16095,N_15899,N_15604);
xnor U16096 (N_16096,N_15614,N_15664);
nand U16097 (N_16097,N_15655,N_15756);
and U16098 (N_16098,N_15898,N_15665);
nand U16099 (N_16099,N_15673,N_15706);
and U16100 (N_16100,N_15729,N_15625);
and U16101 (N_16101,N_15860,N_15879);
nand U16102 (N_16102,N_15839,N_15727);
nor U16103 (N_16103,N_15848,N_15877);
nand U16104 (N_16104,N_15853,N_15833);
nor U16105 (N_16105,N_15626,N_15635);
nor U16106 (N_16106,N_15805,N_15671);
or U16107 (N_16107,N_15688,N_15718);
and U16108 (N_16108,N_15826,N_15723);
nor U16109 (N_16109,N_15615,N_15870);
nand U16110 (N_16110,N_15789,N_15715);
nand U16111 (N_16111,N_15776,N_15881);
nor U16112 (N_16112,N_15806,N_15719);
xnor U16113 (N_16113,N_15608,N_15627);
nor U16114 (N_16114,N_15792,N_15854);
or U16115 (N_16115,N_15753,N_15662);
nand U16116 (N_16116,N_15824,N_15826);
nand U16117 (N_16117,N_15663,N_15748);
nand U16118 (N_16118,N_15887,N_15649);
and U16119 (N_16119,N_15703,N_15757);
xor U16120 (N_16120,N_15705,N_15888);
xnor U16121 (N_16121,N_15816,N_15694);
xnor U16122 (N_16122,N_15623,N_15780);
and U16123 (N_16123,N_15887,N_15716);
nand U16124 (N_16124,N_15602,N_15809);
xor U16125 (N_16125,N_15606,N_15845);
or U16126 (N_16126,N_15860,N_15847);
nand U16127 (N_16127,N_15671,N_15820);
nand U16128 (N_16128,N_15764,N_15824);
nand U16129 (N_16129,N_15779,N_15882);
or U16130 (N_16130,N_15690,N_15804);
and U16131 (N_16131,N_15624,N_15659);
or U16132 (N_16132,N_15785,N_15896);
nand U16133 (N_16133,N_15631,N_15851);
and U16134 (N_16134,N_15622,N_15702);
nand U16135 (N_16135,N_15697,N_15883);
xor U16136 (N_16136,N_15888,N_15681);
xor U16137 (N_16137,N_15677,N_15814);
nor U16138 (N_16138,N_15661,N_15822);
xor U16139 (N_16139,N_15750,N_15748);
or U16140 (N_16140,N_15670,N_15623);
xnor U16141 (N_16141,N_15701,N_15756);
nand U16142 (N_16142,N_15617,N_15817);
nor U16143 (N_16143,N_15885,N_15612);
nor U16144 (N_16144,N_15819,N_15634);
xnor U16145 (N_16145,N_15807,N_15752);
xnor U16146 (N_16146,N_15730,N_15734);
or U16147 (N_16147,N_15623,N_15777);
nand U16148 (N_16148,N_15638,N_15864);
xor U16149 (N_16149,N_15705,N_15617);
or U16150 (N_16150,N_15813,N_15841);
nand U16151 (N_16151,N_15816,N_15851);
nand U16152 (N_16152,N_15896,N_15669);
nor U16153 (N_16153,N_15750,N_15869);
nand U16154 (N_16154,N_15678,N_15695);
nor U16155 (N_16155,N_15778,N_15704);
nor U16156 (N_16156,N_15778,N_15740);
nand U16157 (N_16157,N_15758,N_15642);
or U16158 (N_16158,N_15879,N_15736);
xor U16159 (N_16159,N_15816,N_15847);
or U16160 (N_16160,N_15809,N_15647);
and U16161 (N_16161,N_15859,N_15834);
nor U16162 (N_16162,N_15731,N_15769);
xnor U16163 (N_16163,N_15611,N_15661);
xor U16164 (N_16164,N_15632,N_15672);
or U16165 (N_16165,N_15834,N_15815);
nand U16166 (N_16166,N_15719,N_15700);
nor U16167 (N_16167,N_15651,N_15867);
nand U16168 (N_16168,N_15686,N_15601);
xor U16169 (N_16169,N_15796,N_15795);
or U16170 (N_16170,N_15875,N_15612);
xor U16171 (N_16171,N_15678,N_15749);
xor U16172 (N_16172,N_15736,N_15637);
nor U16173 (N_16173,N_15833,N_15781);
xor U16174 (N_16174,N_15876,N_15814);
nand U16175 (N_16175,N_15628,N_15803);
nand U16176 (N_16176,N_15678,N_15739);
nor U16177 (N_16177,N_15872,N_15776);
and U16178 (N_16178,N_15812,N_15625);
nor U16179 (N_16179,N_15887,N_15605);
xor U16180 (N_16180,N_15854,N_15682);
nand U16181 (N_16181,N_15713,N_15618);
or U16182 (N_16182,N_15702,N_15639);
xnor U16183 (N_16183,N_15873,N_15868);
nand U16184 (N_16184,N_15850,N_15751);
nor U16185 (N_16185,N_15793,N_15663);
nand U16186 (N_16186,N_15765,N_15613);
nor U16187 (N_16187,N_15732,N_15826);
or U16188 (N_16188,N_15759,N_15747);
nor U16189 (N_16189,N_15669,N_15796);
nand U16190 (N_16190,N_15776,N_15825);
and U16191 (N_16191,N_15651,N_15686);
xnor U16192 (N_16192,N_15719,N_15751);
nand U16193 (N_16193,N_15857,N_15827);
xor U16194 (N_16194,N_15623,N_15790);
nor U16195 (N_16195,N_15858,N_15652);
and U16196 (N_16196,N_15644,N_15608);
or U16197 (N_16197,N_15742,N_15694);
or U16198 (N_16198,N_15658,N_15718);
nor U16199 (N_16199,N_15672,N_15746);
xnor U16200 (N_16200,N_16005,N_16061);
and U16201 (N_16201,N_15924,N_15986);
xnor U16202 (N_16202,N_15979,N_16152);
xor U16203 (N_16203,N_16171,N_16058);
nor U16204 (N_16204,N_15908,N_16069);
nand U16205 (N_16205,N_16191,N_16143);
nor U16206 (N_16206,N_15915,N_16119);
nand U16207 (N_16207,N_15993,N_15948);
and U16208 (N_16208,N_16177,N_16111);
xnor U16209 (N_16209,N_16195,N_15933);
nor U16210 (N_16210,N_15928,N_15999);
and U16211 (N_16211,N_16006,N_16052);
and U16212 (N_16212,N_16010,N_16108);
xnor U16213 (N_16213,N_16097,N_16187);
and U16214 (N_16214,N_16055,N_16031);
nand U16215 (N_16215,N_16003,N_15920);
nor U16216 (N_16216,N_16109,N_16157);
xor U16217 (N_16217,N_15909,N_16062);
xor U16218 (N_16218,N_16159,N_16064);
nor U16219 (N_16219,N_16140,N_16011);
or U16220 (N_16220,N_16093,N_15944);
nand U16221 (N_16221,N_16167,N_16092);
nor U16222 (N_16222,N_15932,N_16023);
or U16223 (N_16223,N_16176,N_16007);
nor U16224 (N_16224,N_15929,N_16013);
and U16225 (N_16225,N_16183,N_16138);
and U16226 (N_16226,N_16017,N_15907);
xor U16227 (N_16227,N_16089,N_16053);
xor U16228 (N_16228,N_16146,N_16197);
xor U16229 (N_16229,N_16118,N_16084);
nand U16230 (N_16230,N_15974,N_16001);
or U16231 (N_16231,N_16036,N_15900);
nor U16232 (N_16232,N_16170,N_16156);
nor U16233 (N_16233,N_16014,N_16051);
xor U16234 (N_16234,N_16116,N_16033);
and U16235 (N_16235,N_15966,N_16066);
and U16236 (N_16236,N_16040,N_15936);
and U16237 (N_16237,N_16161,N_16027);
nor U16238 (N_16238,N_16004,N_16144);
and U16239 (N_16239,N_16002,N_15923);
or U16240 (N_16240,N_16076,N_16151);
and U16241 (N_16241,N_16039,N_16080);
xor U16242 (N_16242,N_15984,N_15977);
xnor U16243 (N_16243,N_15946,N_15981);
xnor U16244 (N_16244,N_15978,N_16101);
xnor U16245 (N_16245,N_16065,N_15918);
xor U16246 (N_16246,N_16032,N_16196);
nor U16247 (N_16247,N_16135,N_16120);
xor U16248 (N_16248,N_16112,N_16188);
and U16249 (N_16249,N_15997,N_15921);
nand U16250 (N_16250,N_15955,N_16085);
xnor U16251 (N_16251,N_16075,N_16150);
and U16252 (N_16252,N_15988,N_16077);
and U16253 (N_16253,N_15991,N_15911);
or U16254 (N_16254,N_16181,N_15992);
or U16255 (N_16255,N_15970,N_16153);
xnor U16256 (N_16256,N_16030,N_15973);
or U16257 (N_16257,N_16175,N_16100);
and U16258 (N_16258,N_16132,N_16133);
or U16259 (N_16259,N_16198,N_16098);
nand U16260 (N_16260,N_16178,N_16121);
or U16261 (N_16261,N_16193,N_16019);
xnor U16262 (N_16262,N_16130,N_15931);
nand U16263 (N_16263,N_16071,N_16042);
xnor U16264 (N_16264,N_15951,N_16173);
and U16265 (N_16265,N_16012,N_16049);
or U16266 (N_16266,N_16045,N_16035);
and U16267 (N_16267,N_15935,N_16041);
nand U16268 (N_16268,N_16018,N_16048);
xor U16269 (N_16269,N_15938,N_16127);
xor U16270 (N_16270,N_15960,N_16190);
xnor U16271 (N_16271,N_16148,N_16182);
xor U16272 (N_16272,N_15971,N_15963);
and U16273 (N_16273,N_15904,N_16192);
nor U16274 (N_16274,N_16091,N_16180);
xnor U16275 (N_16275,N_15913,N_16113);
xnor U16276 (N_16276,N_16028,N_16057);
nand U16277 (N_16277,N_16154,N_16060);
xor U16278 (N_16278,N_16141,N_16184);
nor U16279 (N_16279,N_15925,N_15906);
xnor U16280 (N_16280,N_15954,N_16126);
nor U16281 (N_16281,N_15937,N_16043);
xor U16282 (N_16282,N_15917,N_16068);
nor U16283 (N_16283,N_15957,N_16082);
and U16284 (N_16284,N_15902,N_15952);
xor U16285 (N_16285,N_16034,N_16199);
or U16286 (N_16286,N_15901,N_15961);
and U16287 (N_16287,N_16106,N_16088);
xnor U16288 (N_16288,N_15922,N_16072);
nand U16289 (N_16289,N_16074,N_16166);
xor U16290 (N_16290,N_16087,N_16086);
or U16291 (N_16291,N_16185,N_15934);
and U16292 (N_16292,N_16169,N_15975);
xor U16293 (N_16293,N_15916,N_15903);
or U16294 (N_16294,N_16090,N_15995);
xor U16295 (N_16295,N_16162,N_15976);
nor U16296 (N_16296,N_16024,N_16059);
nand U16297 (N_16297,N_15956,N_16047);
nand U16298 (N_16298,N_16164,N_15926);
and U16299 (N_16299,N_16103,N_16131);
xnor U16300 (N_16300,N_16020,N_15927);
nand U16301 (N_16301,N_16015,N_16070);
or U16302 (N_16302,N_16147,N_16021);
xor U16303 (N_16303,N_15940,N_15950);
nand U16304 (N_16304,N_15980,N_15914);
nor U16305 (N_16305,N_15959,N_16142);
nor U16306 (N_16306,N_15947,N_15964);
nor U16307 (N_16307,N_15941,N_16009);
nor U16308 (N_16308,N_16029,N_16163);
or U16309 (N_16309,N_16063,N_15905);
or U16310 (N_16310,N_16044,N_16160);
xnor U16311 (N_16311,N_15953,N_15942);
or U16312 (N_16312,N_16155,N_15945);
nor U16313 (N_16313,N_16025,N_16114);
or U16314 (N_16314,N_16158,N_16179);
and U16315 (N_16315,N_15919,N_15990);
xor U16316 (N_16316,N_16000,N_15939);
xnor U16317 (N_16317,N_16168,N_15987);
xnor U16318 (N_16318,N_15930,N_16139);
or U16319 (N_16319,N_16189,N_16096);
or U16320 (N_16320,N_16137,N_16078);
or U16321 (N_16321,N_16136,N_15912);
xnor U16322 (N_16322,N_16067,N_15994);
or U16323 (N_16323,N_16099,N_16038);
or U16324 (N_16324,N_16115,N_15982);
or U16325 (N_16325,N_16008,N_16124);
or U16326 (N_16326,N_16110,N_15958);
nand U16327 (N_16327,N_16149,N_15969);
or U16328 (N_16328,N_15983,N_16128);
and U16329 (N_16329,N_16050,N_15962);
xnor U16330 (N_16330,N_16134,N_16056);
nand U16331 (N_16331,N_16073,N_15985);
nand U16332 (N_16332,N_16194,N_16125);
or U16333 (N_16333,N_16026,N_15996);
nor U16334 (N_16334,N_16022,N_16172);
or U16335 (N_16335,N_15967,N_15965);
or U16336 (N_16336,N_16095,N_15972);
and U16337 (N_16337,N_16104,N_16037);
and U16338 (N_16338,N_15998,N_15943);
nand U16339 (N_16339,N_15968,N_16054);
nand U16340 (N_16340,N_15949,N_16079);
nor U16341 (N_16341,N_16117,N_16107);
nand U16342 (N_16342,N_16174,N_16123);
or U16343 (N_16343,N_16145,N_15910);
and U16344 (N_16344,N_16129,N_16016);
xor U16345 (N_16345,N_16186,N_16105);
xnor U16346 (N_16346,N_16083,N_16046);
nand U16347 (N_16347,N_16081,N_16122);
xnor U16348 (N_16348,N_16094,N_16102);
nand U16349 (N_16349,N_15989,N_16165);
nand U16350 (N_16350,N_15984,N_15976);
and U16351 (N_16351,N_16160,N_16185);
or U16352 (N_16352,N_16172,N_16056);
nand U16353 (N_16353,N_15971,N_15996);
xnor U16354 (N_16354,N_15932,N_16038);
xnor U16355 (N_16355,N_16069,N_15977);
xnor U16356 (N_16356,N_15901,N_16069);
or U16357 (N_16357,N_15931,N_16197);
xor U16358 (N_16358,N_16137,N_16071);
nand U16359 (N_16359,N_15944,N_16016);
and U16360 (N_16360,N_15917,N_15935);
nand U16361 (N_16361,N_16100,N_15973);
xor U16362 (N_16362,N_15947,N_16063);
nand U16363 (N_16363,N_15957,N_15901);
or U16364 (N_16364,N_16164,N_16138);
nor U16365 (N_16365,N_15987,N_16189);
and U16366 (N_16366,N_15931,N_15971);
nand U16367 (N_16367,N_15962,N_15946);
xnor U16368 (N_16368,N_16188,N_16154);
nor U16369 (N_16369,N_16032,N_16047);
or U16370 (N_16370,N_16001,N_15928);
nand U16371 (N_16371,N_16132,N_15922);
or U16372 (N_16372,N_16133,N_16059);
xnor U16373 (N_16373,N_16069,N_16143);
and U16374 (N_16374,N_16040,N_16190);
or U16375 (N_16375,N_16090,N_15959);
nor U16376 (N_16376,N_16015,N_15932);
xnor U16377 (N_16377,N_15976,N_15967);
nor U16378 (N_16378,N_16100,N_15984);
nand U16379 (N_16379,N_16052,N_16051);
xnor U16380 (N_16380,N_16119,N_15932);
nand U16381 (N_16381,N_16195,N_15967);
and U16382 (N_16382,N_15919,N_16113);
nand U16383 (N_16383,N_16139,N_15968);
nand U16384 (N_16384,N_15994,N_16060);
or U16385 (N_16385,N_16061,N_15978);
xor U16386 (N_16386,N_15934,N_16036);
nor U16387 (N_16387,N_15973,N_16094);
xor U16388 (N_16388,N_15914,N_16017);
xnor U16389 (N_16389,N_16176,N_16114);
or U16390 (N_16390,N_16120,N_15908);
nor U16391 (N_16391,N_15969,N_15980);
xnor U16392 (N_16392,N_16098,N_16130);
xor U16393 (N_16393,N_15963,N_16159);
or U16394 (N_16394,N_16092,N_16038);
and U16395 (N_16395,N_16008,N_16058);
nor U16396 (N_16396,N_16085,N_16105);
xor U16397 (N_16397,N_15964,N_16159);
nor U16398 (N_16398,N_16193,N_15927);
nor U16399 (N_16399,N_15978,N_16163);
xnor U16400 (N_16400,N_16057,N_16077);
nand U16401 (N_16401,N_16139,N_15909);
nand U16402 (N_16402,N_15963,N_15945);
and U16403 (N_16403,N_16197,N_16124);
or U16404 (N_16404,N_16140,N_16108);
xor U16405 (N_16405,N_16054,N_15992);
or U16406 (N_16406,N_16120,N_16045);
xor U16407 (N_16407,N_16199,N_16054);
or U16408 (N_16408,N_15960,N_16130);
and U16409 (N_16409,N_16175,N_15909);
nand U16410 (N_16410,N_15945,N_16001);
nor U16411 (N_16411,N_16062,N_16092);
or U16412 (N_16412,N_16129,N_15956);
nand U16413 (N_16413,N_16099,N_16132);
and U16414 (N_16414,N_16192,N_15999);
xnor U16415 (N_16415,N_16055,N_16117);
and U16416 (N_16416,N_16181,N_15902);
xor U16417 (N_16417,N_16031,N_15975);
or U16418 (N_16418,N_15955,N_16125);
and U16419 (N_16419,N_15914,N_15925);
nand U16420 (N_16420,N_16036,N_16024);
or U16421 (N_16421,N_16088,N_16067);
xor U16422 (N_16422,N_15933,N_16101);
nor U16423 (N_16423,N_16021,N_15955);
nand U16424 (N_16424,N_15956,N_16161);
and U16425 (N_16425,N_15999,N_16107);
nor U16426 (N_16426,N_16174,N_15994);
xnor U16427 (N_16427,N_16189,N_16037);
or U16428 (N_16428,N_15910,N_15962);
and U16429 (N_16429,N_15987,N_16015);
or U16430 (N_16430,N_16095,N_16021);
or U16431 (N_16431,N_16109,N_15922);
or U16432 (N_16432,N_16056,N_15924);
nand U16433 (N_16433,N_16153,N_16113);
xnor U16434 (N_16434,N_15999,N_16053);
and U16435 (N_16435,N_16017,N_16011);
nor U16436 (N_16436,N_16014,N_16105);
nand U16437 (N_16437,N_16031,N_16140);
or U16438 (N_16438,N_16064,N_15965);
or U16439 (N_16439,N_15971,N_16117);
and U16440 (N_16440,N_15992,N_16153);
or U16441 (N_16441,N_16066,N_16076);
or U16442 (N_16442,N_16054,N_16104);
xor U16443 (N_16443,N_16189,N_15974);
or U16444 (N_16444,N_16155,N_15927);
nand U16445 (N_16445,N_16037,N_16038);
nor U16446 (N_16446,N_16187,N_15937);
xnor U16447 (N_16447,N_16086,N_15942);
nor U16448 (N_16448,N_16130,N_16061);
nand U16449 (N_16449,N_16077,N_16182);
and U16450 (N_16450,N_16046,N_16030);
nor U16451 (N_16451,N_15989,N_16145);
nand U16452 (N_16452,N_16175,N_16052);
or U16453 (N_16453,N_16181,N_15981);
xnor U16454 (N_16454,N_16095,N_16027);
nor U16455 (N_16455,N_16161,N_15972);
xnor U16456 (N_16456,N_16018,N_16044);
or U16457 (N_16457,N_16186,N_16092);
xnor U16458 (N_16458,N_16181,N_16192);
and U16459 (N_16459,N_16045,N_16110);
xor U16460 (N_16460,N_16074,N_16185);
nor U16461 (N_16461,N_16101,N_16147);
nor U16462 (N_16462,N_16001,N_16018);
nor U16463 (N_16463,N_16017,N_15937);
or U16464 (N_16464,N_16106,N_15922);
xnor U16465 (N_16465,N_16166,N_16050);
nor U16466 (N_16466,N_16169,N_15970);
nor U16467 (N_16467,N_16020,N_16053);
xor U16468 (N_16468,N_15938,N_16169);
or U16469 (N_16469,N_16004,N_15984);
xnor U16470 (N_16470,N_15939,N_15971);
nor U16471 (N_16471,N_16079,N_16143);
nor U16472 (N_16472,N_15924,N_16085);
nor U16473 (N_16473,N_16192,N_16114);
xnor U16474 (N_16474,N_16150,N_15904);
xnor U16475 (N_16475,N_16114,N_16000);
and U16476 (N_16476,N_16110,N_16109);
nor U16477 (N_16477,N_15971,N_15978);
or U16478 (N_16478,N_16167,N_16081);
xnor U16479 (N_16479,N_16073,N_15991);
or U16480 (N_16480,N_16151,N_15972);
nand U16481 (N_16481,N_16025,N_16023);
xor U16482 (N_16482,N_16039,N_16122);
xnor U16483 (N_16483,N_16044,N_16015);
nand U16484 (N_16484,N_16152,N_15951);
or U16485 (N_16485,N_15911,N_16049);
nor U16486 (N_16486,N_16171,N_16116);
nand U16487 (N_16487,N_16063,N_15959);
nand U16488 (N_16488,N_16150,N_16187);
or U16489 (N_16489,N_15960,N_16114);
xnor U16490 (N_16490,N_16154,N_15943);
xor U16491 (N_16491,N_15934,N_15994);
xor U16492 (N_16492,N_15988,N_15977);
nor U16493 (N_16493,N_16156,N_16108);
nor U16494 (N_16494,N_16056,N_15900);
or U16495 (N_16495,N_15917,N_15949);
nand U16496 (N_16496,N_16126,N_15929);
nand U16497 (N_16497,N_15941,N_15996);
or U16498 (N_16498,N_16148,N_16188);
nand U16499 (N_16499,N_16115,N_15925);
or U16500 (N_16500,N_16330,N_16249);
or U16501 (N_16501,N_16488,N_16266);
nor U16502 (N_16502,N_16309,N_16333);
nand U16503 (N_16503,N_16247,N_16365);
and U16504 (N_16504,N_16460,N_16338);
and U16505 (N_16505,N_16355,N_16214);
nor U16506 (N_16506,N_16381,N_16363);
nor U16507 (N_16507,N_16229,N_16302);
and U16508 (N_16508,N_16386,N_16335);
and U16509 (N_16509,N_16236,N_16449);
nand U16510 (N_16510,N_16375,N_16201);
and U16511 (N_16511,N_16495,N_16459);
nand U16512 (N_16512,N_16453,N_16348);
nand U16513 (N_16513,N_16341,N_16206);
nor U16514 (N_16514,N_16462,N_16350);
and U16515 (N_16515,N_16432,N_16346);
nand U16516 (N_16516,N_16376,N_16245);
or U16517 (N_16517,N_16398,N_16224);
and U16518 (N_16518,N_16310,N_16467);
or U16519 (N_16519,N_16256,N_16405);
or U16520 (N_16520,N_16480,N_16400);
xor U16521 (N_16521,N_16440,N_16307);
and U16522 (N_16522,N_16272,N_16220);
xor U16523 (N_16523,N_16336,N_16288);
and U16524 (N_16524,N_16326,N_16429);
xnor U16525 (N_16525,N_16286,N_16457);
xor U16526 (N_16526,N_16478,N_16441);
nor U16527 (N_16527,N_16215,N_16418);
xor U16528 (N_16528,N_16489,N_16209);
xor U16529 (N_16529,N_16444,N_16268);
or U16530 (N_16530,N_16347,N_16411);
nand U16531 (N_16531,N_16474,N_16316);
nand U16532 (N_16532,N_16237,N_16402);
nor U16533 (N_16533,N_16379,N_16234);
xnor U16534 (N_16534,N_16223,N_16371);
nand U16535 (N_16535,N_16282,N_16303);
and U16536 (N_16536,N_16290,N_16322);
or U16537 (N_16537,N_16461,N_16428);
xnor U16538 (N_16538,N_16472,N_16273);
xor U16539 (N_16539,N_16469,N_16468);
or U16540 (N_16540,N_16210,N_16203);
nor U16541 (N_16541,N_16208,N_16393);
nor U16542 (N_16542,N_16439,N_16354);
nor U16543 (N_16543,N_16325,N_16494);
nand U16544 (N_16544,N_16216,N_16483);
nor U16545 (N_16545,N_16366,N_16205);
nor U16546 (N_16546,N_16443,N_16442);
nand U16547 (N_16547,N_16451,N_16403);
and U16548 (N_16548,N_16491,N_16383);
nand U16549 (N_16549,N_16239,N_16300);
and U16550 (N_16550,N_16254,N_16235);
or U16551 (N_16551,N_16259,N_16269);
or U16552 (N_16552,N_16496,N_16485);
nand U16553 (N_16553,N_16238,N_16240);
nor U16554 (N_16554,N_16301,N_16499);
or U16555 (N_16555,N_16267,N_16378);
or U16556 (N_16556,N_16465,N_16455);
nor U16557 (N_16557,N_16434,N_16388);
nor U16558 (N_16558,N_16463,N_16261);
nand U16559 (N_16559,N_16364,N_16498);
or U16560 (N_16560,N_16321,N_16360);
xor U16561 (N_16561,N_16446,N_16370);
and U16562 (N_16562,N_16222,N_16407);
xor U16563 (N_16563,N_16298,N_16251);
nor U16564 (N_16564,N_16263,N_16389);
xnor U16565 (N_16565,N_16357,N_16327);
nor U16566 (N_16566,N_16277,N_16242);
xor U16567 (N_16567,N_16437,N_16426);
and U16568 (N_16568,N_16404,N_16436);
or U16569 (N_16569,N_16257,N_16226);
xnor U16570 (N_16570,N_16274,N_16427);
and U16571 (N_16571,N_16231,N_16415);
nor U16572 (N_16572,N_16250,N_16482);
and U16573 (N_16573,N_16417,N_16470);
xor U16574 (N_16574,N_16296,N_16204);
nand U16575 (N_16575,N_16359,N_16394);
nand U16576 (N_16576,N_16358,N_16456);
or U16577 (N_16577,N_16291,N_16447);
xnor U16578 (N_16578,N_16227,N_16289);
nor U16579 (N_16579,N_16414,N_16217);
nor U16580 (N_16580,N_16362,N_16372);
nor U16581 (N_16581,N_16243,N_16305);
or U16582 (N_16582,N_16284,N_16320);
and U16583 (N_16583,N_16323,N_16314);
xnor U16584 (N_16584,N_16421,N_16324);
and U16585 (N_16585,N_16343,N_16410);
xnor U16586 (N_16586,N_16315,N_16270);
nand U16587 (N_16587,N_16329,N_16318);
xor U16588 (N_16588,N_16413,N_16262);
or U16589 (N_16589,N_16487,N_16252);
xor U16590 (N_16590,N_16477,N_16382);
and U16591 (N_16591,N_16344,N_16401);
xnor U16592 (N_16592,N_16409,N_16232);
nand U16593 (N_16593,N_16479,N_16304);
and U16594 (N_16594,N_16430,N_16484);
xor U16595 (N_16595,N_16458,N_16221);
nor U16596 (N_16596,N_16431,N_16416);
nor U16597 (N_16597,N_16287,N_16253);
nand U16598 (N_16598,N_16278,N_16373);
nand U16599 (N_16599,N_16280,N_16374);
nor U16600 (N_16600,N_16433,N_16406);
and U16601 (N_16601,N_16248,N_16241);
nand U16602 (N_16602,N_16339,N_16337);
nand U16603 (N_16603,N_16353,N_16424);
nor U16604 (N_16604,N_16448,N_16481);
nor U16605 (N_16605,N_16319,N_16306);
xor U16606 (N_16606,N_16212,N_16297);
nor U16607 (N_16607,N_16377,N_16308);
nor U16608 (N_16608,N_16317,N_16356);
xnor U16609 (N_16609,N_16369,N_16295);
or U16610 (N_16610,N_16328,N_16255);
nand U16611 (N_16611,N_16387,N_16420);
and U16612 (N_16612,N_16258,N_16396);
nor U16613 (N_16613,N_16391,N_16233);
or U16614 (N_16614,N_16361,N_16368);
and U16615 (N_16615,N_16349,N_16345);
nand U16616 (N_16616,N_16207,N_16332);
and U16617 (N_16617,N_16464,N_16312);
and U16618 (N_16618,N_16211,N_16497);
nand U16619 (N_16619,N_16492,N_16294);
or U16620 (N_16620,N_16450,N_16473);
or U16621 (N_16621,N_16385,N_16380);
xnor U16622 (N_16622,N_16202,N_16311);
and U16623 (N_16623,N_16471,N_16419);
nor U16624 (N_16624,N_16265,N_16225);
nor U16625 (N_16625,N_16244,N_16367);
nor U16626 (N_16626,N_16340,N_16200);
xor U16627 (N_16627,N_16331,N_16399);
xnor U16628 (N_16628,N_16218,N_16342);
nand U16629 (N_16629,N_16351,N_16435);
and U16630 (N_16630,N_16293,N_16397);
and U16631 (N_16631,N_16384,N_16422);
xor U16632 (N_16632,N_16228,N_16438);
or U16633 (N_16633,N_16476,N_16445);
nand U16634 (N_16634,N_16392,N_16466);
nand U16635 (N_16635,N_16283,N_16454);
and U16636 (N_16636,N_16271,N_16281);
xor U16637 (N_16637,N_16352,N_16219);
nand U16638 (N_16638,N_16486,N_16475);
xnor U16639 (N_16639,N_16279,N_16246);
or U16640 (N_16640,N_16425,N_16423);
nand U16641 (N_16641,N_16276,N_16260);
and U16642 (N_16642,N_16408,N_16285);
or U16643 (N_16643,N_16313,N_16493);
and U16644 (N_16644,N_16412,N_16230);
or U16645 (N_16645,N_16334,N_16490);
and U16646 (N_16646,N_16390,N_16299);
xor U16647 (N_16647,N_16264,N_16292);
xor U16648 (N_16648,N_16275,N_16452);
nor U16649 (N_16649,N_16213,N_16395);
and U16650 (N_16650,N_16222,N_16282);
nor U16651 (N_16651,N_16301,N_16418);
xnor U16652 (N_16652,N_16247,N_16405);
nand U16653 (N_16653,N_16384,N_16286);
nor U16654 (N_16654,N_16466,N_16469);
and U16655 (N_16655,N_16435,N_16279);
and U16656 (N_16656,N_16457,N_16495);
and U16657 (N_16657,N_16250,N_16420);
xor U16658 (N_16658,N_16355,N_16232);
or U16659 (N_16659,N_16463,N_16241);
nor U16660 (N_16660,N_16304,N_16395);
and U16661 (N_16661,N_16373,N_16308);
and U16662 (N_16662,N_16290,N_16317);
xor U16663 (N_16663,N_16366,N_16376);
nor U16664 (N_16664,N_16483,N_16492);
xor U16665 (N_16665,N_16462,N_16429);
xnor U16666 (N_16666,N_16371,N_16314);
or U16667 (N_16667,N_16392,N_16279);
or U16668 (N_16668,N_16314,N_16266);
nor U16669 (N_16669,N_16393,N_16427);
nor U16670 (N_16670,N_16211,N_16220);
or U16671 (N_16671,N_16435,N_16228);
xor U16672 (N_16672,N_16483,N_16489);
nand U16673 (N_16673,N_16396,N_16219);
or U16674 (N_16674,N_16476,N_16485);
or U16675 (N_16675,N_16272,N_16242);
xor U16676 (N_16676,N_16381,N_16265);
xor U16677 (N_16677,N_16402,N_16475);
or U16678 (N_16678,N_16221,N_16434);
and U16679 (N_16679,N_16344,N_16280);
nand U16680 (N_16680,N_16488,N_16373);
nand U16681 (N_16681,N_16206,N_16413);
and U16682 (N_16682,N_16298,N_16476);
or U16683 (N_16683,N_16229,N_16363);
or U16684 (N_16684,N_16283,N_16469);
and U16685 (N_16685,N_16234,N_16423);
or U16686 (N_16686,N_16410,N_16413);
or U16687 (N_16687,N_16246,N_16380);
and U16688 (N_16688,N_16276,N_16374);
and U16689 (N_16689,N_16327,N_16353);
nand U16690 (N_16690,N_16489,N_16219);
nor U16691 (N_16691,N_16406,N_16403);
and U16692 (N_16692,N_16488,N_16290);
nand U16693 (N_16693,N_16361,N_16348);
xor U16694 (N_16694,N_16317,N_16414);
xor U16695 (N_16695,N_16226,N_16378);
nand U16696 (N_16696,N_16428,N_16245);
or U16697 (N_16697,N_16302,N_16231);
nand U16698 (N_16698,N_16491,N_16282);
and U16699 (N_16699,N_16369,N_16386);
and U16700 (N_16700,N_16395,N_16437);
nand U16701 (N_16701,N_16301,N_16266);
nand U16702 (N_16702,N_16396,N_16304);
nand U16703 (N_16703,N_16243,N_16364);
nor U16704 (N_16704,N_16337,N_16363);
xnor U16705 (N_16705,N_16468,N_16381);
nor U16706 (N_16706,N_16489,N_16343);
and U16707 (N_16707,N_16407,N_16237);
xor U16708 (N_16708,N_16270,N_16253);
and U16709 (N_16709,N_16237,N_16254);
or U16710 (N_16710,N_16297,N_16441);
xnor U16711 (N_16711,N_16242,N_16443);
nor U16712 (N_16712,N_16480,N_16342);
nand U16713 (N_16713,N_16335,N_16305);
nand U16714 (N_16714,N_16468,N_16208);
and U16715 (N_16715,N_16233,N_16269);
xor U16716 (N_16716,N_16368,N_16313);
xnor U16717 (N_16717,N_16216,N_16380);
and U16718 (N_16718,N_16314,N_16251);
and U16719 (N_16719,N_16477,N_16465);
nor U16720 (N_16720,N_16264,N_16451);
nand U16721 (N_16721,N_16259,N_16433);
nor U16722 (N_16722,N_16452,N_16304);
or U16723 (N_16723,N_16469,N_16445);
and U16724 (N_16724,N_16494,N_16477);
nand U16725 (N_16725,N_16451,N_16477);
xor U16726 (N_16726,N_16303,N_16245);
xor U16727 (N_16727,N_16289,N_16343);
and U16728 (N_16728,N_16237,N_16247);
nand U16729 (N_16729,N_16492,N_16319);
and U16730 (N_16730,N_16440,N_16400);
or U16731 (N_16731,N_16469,N_16435);
nor U16732 (N_16732,N_16482,N_16440);
nand U16733 (N_16733,N_16285,N_16324);
and U16734 (N_16734,N_16401,N_16305);
nor U16735 (N_16735,N_16403,N_16302);
nand U16736 (N_16736,N_16255,N_16410);
and U16737 (N_16737,N_16356,N_16499);
nor U16738 (N_16738,N_16381,N_16404);
and U16739 (N_16739,N_16312,N_16377);
xnor U16740 (N_16740,N_16404,N_16482);
nand U16741 (N_16741,N_16278,N_16452);
or U16742 (N_16742,N_16267,N_16462);
nand U16743 (N_16743,N_16314,N_16307);
and U16744 (N_16744,N_16325,N_16303);
or U16745 (N_16745,N_16425,N_16364);
and U16746 (N_16746,N_16230,N_16400);
and U16747 (N_16747,N_16410,N_16498);
or U16748 (N_16748,N_16345,N_16211);
xor U16749 (N_16749,N_16490,N_16426);
nor U16750 (N_16750,N_16281,N_16347);
nand U16751 (N_16751,N_16474,N_16223);
nand U16752 (N_16752,N_16388,N_16409);
xnor U16753 (N_16753,N_16477,N_16234);
nor U16754 (N_16754,N_16300,N_16474);
nor U16755 (N_16755,N_16279,N_16366);
nand U16756 (N_16756,N_16484,N_16332);
nor U16757 (N_16757,N_16386,N_16266);
xnor U16758 (N_16758,N_16491,N_16312);
nor U16759 (N_16759,N_16422,N_16203);
xor U16760 (N_16760,N_16263,N_16246);
or U16761 (N_16761,N_16208,N_16485);
nand U16762 (N_16762,N_16293,N_16482);
xor U16763 (N_16763,N_16248,N_16299);
nand U16764 (N_16764,N_16424,N_16387);
nor U16765 (N_16765,N_16483,N_16229);
nor U16766 (N_16766,N_16353,N_16245);
nor U16767 (N_16767,N_16328,N_16486);
and U16768 (N_16768,N_16386,N_16292);
and U16769 (N_16769,N_16404,N_16388);
and U16770 (N_16770,N_16348,N_16233);
or U16771 (N_16771,N_16354,N_16449);
or U16772 (N_16772,N_16414,N_16256);
nand U16773 (N_16773,N_16270,N_16237);
xnor U16774 (N_16774,N_16340,N_16222);
nand U16775 (N_16775,N_16443,N_16460);
nand U16776 (N_16776,N_16326,N_16379);
xor U16777 (N_16777,N_16413,N_16246);
nand U16778 (N_16778,N_16329,N_16495);
and U16779 (N_16779,N_16277,N_16216);
or U16780 (N_16780,N_16425,N_16479);
nor U16781 (N_16781,N_16417,N_16388);
xor U16782 (N_16782,N_16202,N_16267);
or U16783 (N_16783,N_16393,N_16336);
or U16784 (N_16784,N_16223,N_16320);
or U16785 (N_16785,N_16355,N_16296);
or U16786 (N_16786,N_16425,N_16206);
and U16787 (N_16787,N_16255,N_16366);
and U16788 (N_16788,N_16494,N_16276);
xnor U16789 (N_16789,N_16246,N_16376);
and U16790 (N_16790,N_16475,N_16328);
nor U16791 (N_16791,N_16231,N_16411);
xor U16792 (N_16792,N_16252,N_16373);
xor U16793 (N_16793,N_16497,N_16307);
or U16794 (N_16794,N_16252,N_16282);
and U16795 (N_16795,N_16442,N_16448);
nor U16796 (N_16796,N_16218,N_16279);
nor U16797 (N_16797,N_16242,N_16210);
xor U16798 (N_16798,N_16447,N_16266);
or U16799 (N_16799,N_16369,N_16232);
xor U16800 (N_16800,N_16773,N_16628);
and U16801 (N_16801,N_16639,N_16621);
nor U16802 (N_16802,N_16502,N_16602);
and U16803 (N_16803,N_16721,N_16515);
or U16804 (N_16804,N_16747,N_16665);
nor U16805 (N_16805,N_16505,N_16730);
or U16806 (N_16806,N_16589,N_16618);
nand U16807 (N_16807,N_16526,N_16561);
and U16808 (N_16808,N_16736,N_16764);
nor U16809 (N_16809,N_16507,N_16658);
or U16810 (N_16810,N_16694,N_16574);
nand U16811 (N_16811,N_16788,N_16701);
xnor U16812 (N_16812,N_16546,N_16751);
nor U16813 (N_16813,N_16514,N_16604);
nor U16814 (N_16814,N_16655,N_16672);
nand U16815 (N_16815,N_16785,N_16793);
nand U16816 (N_16816,N_16552,N_16758);
nor U16817 (N_16817,N_16620,N_16740);
and U16818 (N_16818,N_16714,N_16642);
nand U16819 (N_16819,N_16743,N_16682);
and U16820 (N_16820,N_16738,N_16709);
or U16821 (N_16821,N_16799,N_16622);
and U16822 (N_16822,N_16616,N_16756);
and U16823 (N_16823,N_16518,N_16568);
nor U16824 (N_16824,N_16791,N_16543);
and U16825 (N_16825,N_16650,N_16713);
or U16826 (N_16826,N_16702,N_16549);
nor U16827 (N_16827,N_16688,N_16733);
xor U16828 (N_16828,N_16767,N_16661);
xor U16829 (N_16829,N_16557,N_16741);
xor U16830 (N_16830,N_16653,N_16536);
or U16831 (N_16831,N_16573,N_16582);
nor U16832 (N_16832,N_16725,N_16748);
and U16833 (N_16833,N_16731,N_16699);
and U16834 (N_16834,N_16648,N_16664);
nand U16835 (N_16835,N_16692,N_16676);
xor U16836 (N_16836,N_16600,N_16592);
nor U16837 (N_16837,N_16757,N_16569);
and U16838 (N_16838,N_16601,N_16584);
and U16839 (N_16839,N_16563,N_16691);
nor U16840 (N_16840,N_16529,N_16698);
nand U16841 (N_16841,N_16558,N_16525);
xnor U16842 (N_16842,N_16739,N_16707);
nand U16843 (N_16843,N_16774,N_16528);
and U16844 (N_16844,N_16723,N_16689);
and U16845 (N_16845,N_16541,N_16567);
xor U16846 (N_16846,N_16542,N_16570);
xnor U16847 (N_16847,N_16660,N_16645);
xnor U16848 (N_16848,N_16704,N_16718);
and U16849 (N_16849,N_16717,N_16555);
and U16850 (N_16850,N_16797,N_16624);
or U16851 (N_16851,N_16706,N_16777);
or U16852 (N_16852,N_16548,N_16535);
nand U16853 (N_16853,N_16551,N_16609);
xor U16854 (N_16854,N_16783,N_16659);
nor U16855 (N_16855,N_16632,N_16790);
or U16856 (N_16856,N_16629,N_16610);
xor U16857 (N_16857,N_16564,N_16786);
xor U16858 (N_16858,N_16781,N_16550);
xor U16859 (N_16859,N_16657,N_16695);
or U16860 (N_16860,N_16735,N_16680);
and U16861 (N_16861,N_16517,N_16575);
and U16862 (N_16862,N_16670,N_16571);
and U16863 (N_16863,N_16605,N_16510);
and U16864 (N_16864,N_16651,N_16649);
nand U16865 (N_16865,N_16681,N_16583);
nand U16866 (N_16866,N_16656,N_16627);
or U16867 (N_16867,N_16727,N_16544);
nand U16868 (N_16868,N_16646,N_16522);
nor U16869 (N_16869,N_16673,N_16782);
nor U16870 (N_16870,N_16641,N_16608);
or U16871 (N_16871,N_16690,N_16539);
or U16872 (N_16872,N_16524,N_16623);
or U16873 (N_16873,N_16637,N_16588);
nand U16874 (N_16874,N_16662,N_16780);
and U16875 (N_16875,N_16719,N_16615);
xnor U16876 (N_16876,N_16532,N_16565);
nor U16877 (N_16877,N_16737,N_16652);
nor U16878 (N_16878,N_16679,N_16769);
xor U16879 (N_16879,N_16590,N_16547);
or U16880 (N_16880,N_16722,N_16697);
xor U16881 (N_16881,N_16511,N_16766);
nor U16882 (N_16882,N_16603,N_16531);
nor U16883 (N_16883,N_16716,N_16579);
and U16884 (N_16884,N_16753,N_16634);
and U16885 (N_16885,N_16776,N_16765);
nand U16886 (N_16886,N_16527,N_16729);
nand U16887 (N_16887,N_16724,N_16626);
nand U16888 (N_16888,N_16668,N_16761);
xor U16889 (N_16889,N_16612,N_16734);
and U16890 (N_16890,N_16644,N_16666);
xor U16891 (N_16891,N_16566,N_16554);
nand U16892 (N_16892,N_16763,N_16770);
nor U16893 (N_16893,N_16674,N_16576);
xor U16894 (N_16894,N_16631,N_16562);
xor U16895 (N_16895,N_16708,N_16560);
and U16896 (N_16896,N_16762,N_16710);
xnor U16897 (N_16897,N_16586,N_16556);
nand U16898 (N_16898,N_16503,N_16508);
nor U16899 (N_16899,N_16611,N_16537);
and U16900 (N_16900,N_16768,N_16684);
and U16901 (N_16901,N_16696,N_16572);
xnor U16902 (N_16902,N_16669,N_16501);
and U16903 (N_16903,N_16760,N_16654);
or U16904 (N_16904,N_16530,N_16521);
and U16905 (N_16905,N_16752,N_16686);
xnor U16906 (N_16906,N_16726,N_16509);
nand U16907 (N_16907,N_16771,N_16540);
xnor U16908 (N_16908,N_16607,N_16678);
and U16909 (N_16909,N_16593,N_16640);
and U16910 (N_16910,N_16591,N_16712);
nand U16911 (N_16911,N_16580,N_16513);
xnor U16912 (N_16912,N_16784,N_16772);
nand U16913 (N_16913,N_16789,N_16630);
nand U16914 (N_16914,N_16545,N_16643);
nor U16915 (N_16915,N_16559,N_16625);
or U16916 (N_16916,N_16534,N_16705);
nor U16917 (N_16917,N_16581,N_16500);
nand U16918 (N_16918,N_16796,N_16671);
or U16919 (N_16919,N_16750,N_16663);
nand U16920 (N_16920,N_16596,N_16595);
or U16921 (N_16921,N_16597,N_16614);
and U16922 (N_16922,N_16599,N_16746);
or U16923 (N_16923,N_16720,N_16728);
or U16924 (N_16924,N_16617,N_16598);
nor U16925 (N_16925,N_16755,N_16693);
nand U16926 (N_16926,N_16744,N_16578);
or U16927 (N_16927,N_16647,N_16754);
xnor U16928 (N_16928,N_16533,N_16538);
xor U16929 (N_16929,N_16606,N_16506);
nand U16930 (N_16930,N_16700,N_16520);
nand U16931 (N_16931,N_16795,N_16779);
xor U16932 (N_16932,N_16685,N_16778);
or U16933 (N_16933,N_16635,N_16577);
xnor U16934 (N_16934,N_16636,N_16504);
nor U16935 (N_16935,N_16775,N_16794);
or U16936 (N_16936,N_16553,N_16798);
and U16937 (N_16937,N_16633,N_16745);
nor U16938 (N_16938,N_16749,N_16677);
xor U16939 (N_16939,N_16742,N_16759);
or U16940 (N_16940,N_16523,N_16613);
or U16941 (N_16941,N_16594,N_16711);
xnor U16942 (N_16942,N_16638,N_16675);
nand U16943 (N_16943,N_16703,N_16687);
xor U16944 (N_16944,N_16619,N_16516);
nor U16945 (N_16945,N_16519,N_16683);
xor U16946 (N_16946,N_16667,N_16585);
or U16947 (N_16947,N_16715,N_16512);
nand U16948 (N_16948,N_16587,N_16732);
or U16949 (N_16949,N_16787,N_16792);
or U16950 (N_16950,N_16592,N_16551);
or U16951 (N_16951,N_16563,N_16795);
and U16952 (N_16952,N_16628,N_16562);
nor U16953 (N_16953,N_16795,N_16682);
xnor U16954 (N_16954,N_16580,N_16693);
or U16955 (N_16955,N_16592,N_16635);
and U16956 (N_16956,N_16537,N_16739);
nor U16957 (N_16957,N_16568,N_16576);
xnor U16958 (N_16958,N_16554,N_16783);
nand U16959 (N_16959,N_16730,N_16749);
and U16960 (N_16960,N_16766,N_16759);
xnor U16961 (N_16961,N_16716,N_16692);
nand U16962 (N_16962,N_16540,N_16510);
and U16963 (N_16963,N_16649,N_16507);
xnor U16964 (N_16964,N_16586,N_16581);
or U16965 (N_16965,N_16704,N_16735);
xor U16966 (N_16966,N_16525,N_16695);
or U16967 (N_16967,N_16530,N_16758);
nand U16968 (N_16968,N_16512,N_16644);
and U16969 (N_16969,N_16571,N_16651);
nand U16970 (N_16970,N_16594,N_16569);
xnor U16971 (N_16971,N_16742,N_16616);
nor U16972 (N_16972,N_16546,N_16531);
nor U16973 (N_16973,N_16661,N_16590);
or U16974 (N_16974,N_16700,N_16670);
or U16975 (N_16975,N_16590,N_16707);
nand U16976 (N_16976,N_16783,N_16747);
nand U16977 (N_16977,N_16641,N_16530);
or U16978 (N_16978,N_16577,N_16646);
nand U16979 (N_16979,N_16669,N_16568);
and U16980 (N_16980,N_16512,N_16711);
nor U16981 (N_16981,N_16529,N_16671);
nor U16982 (N_16982,N_16637,N_16669);
or U16983 (N_16983,N_16692,N_16697);
and U16984 (N_16984,N_16669,N_16606);
and U16985 (N_16985,N_16524,N_16691);
nand U16986 (N_16986,N_16537,N_16715);
nor U16987 (N_16987,N_16549,N_16625);
xor U16988 (N_16988,N_16524,N_16614);
and U16989 (N_16989,N_16696,N_16618);
or U16990 (N_16990,N_16577,N_16659);
nand U16991 (N_16991,N_16574,N_16680);
nand U16992 (N_16992,N_16686,N_16695);
nand U16993 (N_16993,N_16695,N_16541);
nor U16994 (N_16994,N_16736,N_16500);
or U16995 (N_16995,N_16634,N_16608);
xnor U16996 (N_16996,N_16543,N_16618);
nand U16997 (N_16997,N_16671,N_16595);
xnor U16998 (N_16998,N_16703,N_16562);
xor U16999 (N_16999,N_16576,N_16657);
xor U17000 (N_17000,N_16525,N_16762);
or U17001 (N_17001,N_16544,N_16565);
nand U17002 (N_17002,N_16628,N_16665);
xor U17003 (N_17003,N_16568,N_16655);
nand U17004 (N_17004,N_16583,N_16540);
and U17005 (N_17005,N_16764,N_16556);
and U17006 (N_17006,N_16682,N_16768);
and U17007 (N_17007,N_16643,N_16669);
and U17008 (N_17008,N_16525,N_16680);
xor U17009 (N_17009,N_16660,N_16541);
or U17010 (N_17010,N_16612,N_16666);
nand U17011 (N_17011,N_16598,N_16566);
nand U17012 (N_17012,N_16534,N_16592);
nor U17013 (N_17013,N_16601,N_16585);
nor U17014 (N_17014,N_16534,N_16686);
nand U17015 (N_17015,N_16640,N_16790);
xnor U17016 (N_17016,N_16709,N_16626);
nand U17017 (N_17017,N_16695,N_16565);
xor U17018 (N_17018,N_16774,N_16715);
xor U17019 (N_17019,N_16587,N_16563);
and U17020 (N_17020,N_16574,N_16553);
and U17021 (N_17021,N_16682,N_16551);
and U17022 (N_17022,N_16646,N_16562);
nand U17023 (N_17023,N_16796,N_16718);
nor U17024 (N_17024,N_16609,N_16798);
nand U17025 (N_17025,N_16627,N_16698);
xor U17026 (N_17026,N_16786,N_16739);
xor U17027 (N_17027,N_16709,N_16727);
or U17028 (N_17028,N_16657,N_16621);
xnor U17029 (N_17029,N_16642,N_16718);
or U17030 (N_17030,N_16598,N_16660);
nor U17031 (N_17031,N_16784,N_16613);
nand U17032 (N_17032,N_16629,N_16609);
nor U17033 (N_17033,N_16609,N_16745);
or U17034 (N_17034,N_16640,N_16562);
nor U17035 (N_17035,N_16694,N_16579);
xor U17036 (N_17036,N_16575,N_16576);
nor U17037 (N_17037,N_16764,N_16661);
and U17038 (N_17038,N_16706,N_16575);
nand U17039 (N_17039,N_16673,N_16531);
and U17040 (N_17040,N_16581,N_16658);
xor U17041 (N_17041,N_16519,N_16660);
nor U17042 (N_17042,N_16652,N_16717);
and U17043 (N_17043,N_16739,N_16549);
xor U17044 (N_17044,N_16582,N_16656);
nand U17045 (N_17045,N_16770,N_16713);
xnor U17046 (N_17046,N_16795,N_16586);
nand U17047 (N_17047,N_16691,N_16623);
xnor U17048 (N_17048,N_16626,N_16563);
xnor U17049 (N_17049,N_16549,N_16505);
nor U17050 (N_17050,N_16606,N_16672);
nor U17051 (N_17051,N_16639,N_16605);
nor U17052 (N_17052,N_16657,N_16724);
or U17053 (N_17053,N_16569,N_16598);
nand U17054 (N_17054,N_16784,N_16687);
nand U17055 (N_17055,N_16540,N_16799);
nor U17056 (N_17056,N_16589,N_16504);
nor U17057 (N_17057,N_16570,N_16538);
nand U17058 (N_17058,N_16632,N_16552);
or U17059 (N_17059,N_16537,N_16538);
xnor U17060 (N_17060,N_16718,N_16696);
nand U17061 (N_17061,N_16723,N_16570);
xnor U17062 (N_17062,N_16536,N_16696);
or U17063 (N_17063,N_16755,N_16684);
nand U17064 (N_17064,N_16782,N_16637);
nor U17065 (N_17065,N_16722,N_16744);
nand U17066 (N_17066,N_16631,N_16561);
xnor U17067 (N_17067,N_16561,N_16656);
xor U17068 (N_17068,N_16656,N_16659);
nand U17069 (N_17069,N_16622,N_16522);
nor U17070 (N_17070,N_16561,N_16717);
and U17071 (N_17071,N_16650,N_16620);
or U17072 (N_17072,N_16792,N_16629);
and U17073 (N_17073,N_16669,N_16521);
and U17074 (N_17074,N_16609,N_16502);
nand U17075 (N_17075,N_16636,N_16716);
or U17076 (N_17076,N_16520,N_16529);
and U17077 (N_17077,N_16584,N_16750);
or U17078 (N_17078,N_16765,N_16780);
nor U17079 (N_17079,N_16679,N_16735);
xor U17080 (N_17080,N_16796,N_16522);
or U17081 (N_17081,N_16580,N_16770);
nand U17082 (N_17082,N_16549,N_16556);
or U17083 (N_17083,N_16619,N_16681);
nand U17084 (N_17084,N_16739,N_16669);
or U17085 (N_17085,N_16553,N_16563);
nand U17086 (N_17086,N_16714,N_16538);
and U17087 (N_17087,N_16712,N_16751);
nor U17088 (N_17088,N_16505,N_16718);
xnor U17089 (N_17089,N_16521,N_16650);
and U17090 (N_17090,N_16638,N_16731);
nand U17091 (N_17091,N_16540,N_16525);
or U17092 (N_17092,N_16705,N_16771);
nand U17093 (N_17093,N_16579,N_16646);
xor U17094 (N_17094,N_16580,N_16568);
or U17095 (N_17095,N_16688,N_16703);
or U17096 (N_17096,N_16585,N_16622);
nor U17097 (N_17097,N_16528,N_16630);
xor U17098 (N_17098,N_16577,N_16643);
xnor U17099 (N_17099,N_16608,N_16549);
nand U17100 (N_17100,N_17031,N_17059);
nand U17101 (N_17101,N_16909,N_16953);
or U17102 (N_17102,N_16824,N_17082);
xor U17103 (N_17103,N_17001,N_16809);
nor U17104 (N_17104,N_16859,N_16955);
and U17105 (N_17105,N_16971,N_17045);
or U17106 (N_17106,N_16991,N_16902);
nor U17107 (N_17107,N_17053,N_16911);
and U17108 (N_17108,N_17021,N_16869);
nand U17109 (N_17109,N_17050,N_17039);
nor U17110 (N_17110,N_16881,N_16973);
nor U17111 (N_17111,N_17016,N_17099);
xor U17112 (N_17112,N_17074,N_16999);
or U17113 (N_17113,N_16862,N_17097);
xnor U17114 (N_17114,N_16867,N_16908);
xnor U17115 (N_17115,N_16906,N_16967);
nor U17116 (N_17116,N_16884,N_16885);
xnor U17117 (N_17117,N_16961,N_16812);
nor U17118 (N_17118,N_16913,N_17005);
or U17119 (N_17119,N_16870,N_16849);
or U17120 (N_17120,N_17000,N_17095);
and U17121 (N_17121,N_16817,N_17042);
nor U17122 (N_17122,N_17060,N_16982);
and U17123 (N_17123,N_17062,N_16868);
nand U17124 (N_17124,N_16806,N_17035);
nand U17125 (N_17125,N_17024,N_16843);
nor U17126 (N_17126,N_16924,N_17029);
nor U17127 (N_17127,N_16887,N_16994);
nor U17128 (N_17128,N_16993,N_16872);
xnor U17129 (N_17129,N_17058,N_17033);
and U17130 (N_17130,N_16990,N_16851);
and U17131 (N_17131,N_16828,N_16941);
and U17132 (N_17132,N_16893,N_17073);
nor U17133 (N_17133,N_17046,N_16840);
xor U17134 (N_17134,N_16957,N_17048);
nor U17135 (N_17135,N_17098,N_16878);
and U17136 (N_17136,N_16904,N_17084);
nand U17137 (N_17137,N_16880,N_16853);
nor U17138 (N_17138,N_16834,N_16842);
xor U17139 (N_17139,N_16861,N_16916);
or U17140 (N_17140,N_16979,N_16947);
xor U17141 (N_17141,N_17034,N_16845);
or U17142 (N_17142,N_16949,N_17022);
and U17143 (N_17143,N_17003,N_16960);
xnor U17144 (N_17144,N_16925,N_17094);
nor U17145 (N_17145,N_17085,N_16899);
and U17146 (N_17146,N_16841,N_17040);
nor U17147 (N_17147,N_17087,N_16968);
xnor U17148 (N_17148,N_16896,N_16831);
and U17149 (N_17149,N_16980,N_17066);
nand U17150 (N_17150,N_16879,N_16966);
or U17151 (N_17151,N_16830,N_16901);
xor U17152 (N_17152,N_17043,N_16929);
and U17153 (N_17153,N_16813,N_16937);
or U17154 (N_17154,N_16915,N_16965);
nand U17155 (N_17155,N_16846,N_16989);
and U17156 (N_17156,N_16958,N_17054);
nor U17157 (N_17157,N_17025,N_16964);
nand U17158 (N_17158,N_16921,N_16950);
or U17159 (N_17159,N_17061,N_17044);
nor U17160 (N_17160,N_16818,N_16956);
nand U17161 (N_17161,N_16912,N_16832);
nor U17162 (N_17162,N_16873,N_16850);
and U17163 (N_17163,N_16827,N_17041);
or U17164 (N_17164,N_16829,N_17083);
or U17165 (N_17165,N_16936,N_16839);
or U17166 (N_17166,N_16836,N_16926);
nor U17167 (N_17167,N_16981,N_16805);
and U17168 (N_17168,N_17019,N_17067);
and U17169 (N_17169,N_17006,N_16821);
nand U17170 (N_17170,N_17030,N_17010);
or U17171 (N_17171,N_16808,N_16892);
xor U17172 (N_17172,N_17071,N_16833);
nor U17173 (N_17173,N_16954,N_16985);
nor U17174 (N_17174,N_16814,N_16882);
nor U17175 (N_17175,N_17014,N_16920);
nor U17176 (N_17176,N_16959,N_16876);
and U17177 (N_17177,N_16938,N_17011);
and U17178 (N_17178,N_17091,N_16871);
xnor U17179 (N_17179,N_16835,N_17086);
or U17180 (N_17180,N_16946,N_16847);
nand U17181 (N_17181,N_16826,N_16988);
nor U17182 (N_17182,N_16883,N_17069);
and U17183 (N_17183,N_16939,N_16823);
or U17184 (N_17184,N_17090,N_16919);
and U17185 (N_17185,N_16951,N_17036);
and U17186 (N_17186,N_16927,N_16998);
or U17187 (N_17187,N_16860,N_16837);
and U17188 (N_17188,N_16866,N_16935);
nand U17189 (N_17189,N_16977,N_16903);
xor U17190 (N_17190,N_17049,N_17004);
or U17191 (N_17191,N_16811,N_16969);
xor U17192 (N_17192,N_16931,N_17096);
nand U17193 (N_17193,N_16810,N_16838);
and U17194 (N_17194,N_17078,N_16907);
nor U17195 (N_17195,N_17008,N_16864);
xor U17196 (N_17196,N_16865,N_17081);
or U17197 (N_17197,N_17020,N_16963);
nand U17198 (N_17198,N_17038,N_16975);
and U17199 (N_17199,N_16984,N_16891);
xnor U17200 (N_17200,N_17079,N_16905);
or U17201 (N_17201,N_17013,N_17051);
xnor U17202 (N_17202,N_16945,N_17027);
and U17203 (N_17203,N_16948,N_16804);
and U17204 (N_17204,N_16874,N_16923);
nand U17205 (N_17205,N_17077,N_16888);
xor U17206 (N_17206,N_16942,N_16886);
or U17207 (N_17207,N_16962,N_16848);
or U17208 (N_17208,N_17063,N_16819);
xnor U17209 (N_17209,N_16972,N_16934);
or U17210 (N_17210,N_16943,N_17089);
xnor U17211 (N_17211,N_17028,N_17015);
nor U17212 (N_17212,N_16922,N_17018);
xnor U17213 (N_17213,N_16930,N_16825);
or U17214 (N_17214,N_16890,N_16854);
xor U17215 (N_17215,N_16875,N_16974);
nand U17216 (N_17216,N_17023,N_16918);
xor U17217 (N_17217,N_16910,N_16857);
and U17218 (N_17218,N_16970,N_16816);
or U17219 (N_17219,N_17055,N_16803);
nor U17220 (N_17220,N_17092,N_16801);
nor U17221 (N_17221,N_16952,N_16815);
xnor U17222 (N_17222,N_16822,N_17070);
and U17223 (N_17223,N_16900,N_16940);
nor U17224 (N_17224,N_16983,N_16844);
and U17225 (N_17225,N_16996,N_17080);
xor U17226 (N_17226,N_16894,N_16856);
xnor U17227 (N_17227,N_16995,N_16914);
xnor U17228 (N_17228,N_17026,N_17065);
nor U17229 (N_17229,N_17052,N_16897);
or U17230 (N_17230,N_16986,N_17056);
or U17231 (N_17231,N_17032,N_17002);
nand U17232 (N_17232,N_17012,N_17093);
and U17233 (N_17233,N_16898,N_16877);
xor U17234 (N_17234,N_17007,N_16917);
or U17235 (N_17235,N_16852,N_16928);
nand U17236 (N_17236,N_17009,N_17064);
xor U17237 (N_17237,N_16987,N_17068);
or U17238 (N_17238,N_16800,N_17088);
nand U17239 (N_17239,N_16976,N_16944);
and U17240 (N_17240,N_17072,N_17037);
or U17241 (N_17241,N_16997,N_16889);
nor U17242 (N_17242,N_16807,N_16978);
or U17243 (N_17243,N_17017,N_17057);
or U17244 (N_17244,N_16863,N_16858);
nand U17245 (N_17245,N_16855,N_16992);
and U17246 (N_17246,N_16895,N_16933);
nand U17247 (N_17247,N_16802,N_17075);
and U17248 (N_17248,N_17076,N_16932);
or U17249 (N_17249,N_16820,N_17047);
xnor U17250 (N_17250,N_16957,N_17064);
and U17251 (N_17251,N_16953,N_16986);
nor U17252 (N_17252,N_17018,N_16830);
or U17253 (N_17253,N_17058,N_17092);
xnor U17254 (N_17254,N_16998,N_16844);
xnor U17255 (N_17255,N_17026,N_16813);
and U17256 (N_17256,N_17066,N_17032);
and U17257 (N_17257,N_16985,N_16951);
and U17258 (N_17258,N_16934,N_17059);
xnor U17259 (N_17259,N_16969,N_16817);
nor U17260 (N_17260,N_17036,N_16816);
xnor U17261 (N_17261,N_16876,N_16911);
nor U17262 (N_17262,N_17086,N_16950);
and U17263 (N_17263,N_17075,N_16993);
xor U17264 (N_17264,N_16842,N_16883);
or U17265 (N_17265,N_16862,N_16913);
nand U17266 (N_17266,N_17080,N_17082);
xnor U17267 (N_17267,N_16916,N_17059);
nand U17268 (N_17268,N_17047,N_16834);
nand U17269 (N_17269,N_16912,N_16966);
xnor U17270 (N_17270,N_16974,N_16931);
and U17271 (N_17271,N_16812,N_16864);
xnor U17272 (N_17272,N_17000,N_16945);
nand U17273 (N_17273,N_16980,N_16996);
xor U17274 (N_17274,N_16943,N_16902);
nor U17275 (N_17275,N_16951,N_17064);
xnor U17276 (N_17276,N_16804,N_16878);
nor U17277 (N_17277,N_16978,N_17031);
xor U17278 (N_17278,N_16942,N_16857);
and U17279 (N_17279,N_16833,N_16923);
nand U17280 (N_17280,N_16858,N_16912);
and U17281 (N_17281,N_16850,N_17018);
and U17282 (N_17282,N_17065,N_16969);
xnor U17283 (N_17283,N_16875,N_17070);
nand U17284 (N_17284,N_17091,N_16981);
and U17285 (N_17285,N_17050,N_16972);
xnor U17286 (N_17286,N_16873,N_16981);
nand U17287 (N_17287,N_16954,N_17059);
nand U17288 (N_17288,N_17024,N_16915);
and U17289 (N_17289,N_16944,N_16895);
nor U17290 (N_17290,N_17036,N_16962);
xor U17291 (N_17291,N_16899,N_16898);
xor U17292 (N_17292,N_17058,N_17024);
or U17293 (N_17293,N_16893,N_17016);
or U17294 (N_17294,N_16878,N_16806);
nor U17295 (N_17295,N_16872,N_16932);
nor U17296 (N_17296,N_16831,N_17084);
and U17297 (N_17297,N_16894,N_16826);
and U17298 (N_17298,N_16915,N_16988);
xor U17299 (N_17299,N_16924,N_17025);
xnor U17300 (N_17300,N_17035,N_16895);
or U17301 (N_17301,N_17055,N_16842);
or U17302 (N_17302,N_16831,N_17060);
nor U17303 (N_17303,N_16821,N_16935);
and U17304 (N_17304,N_17079,N_17015);
and U17305 (N_17305,N_17011,N_16836);
xnor U17306 (N_17306,N_16824,N_17076);
nand U17307 (N_17307,N_16891,N_17091);
nor U17308 (N_17308,N_17041,N_16925);
xor U17309 (N_17309,N_17052,N_16941);
nor U17310 (N_17310,N_17028,N_17011);
nor U17311 (N_17311,N_16898,N_16913);
or U17312 (N_17312,N_16889,N_17051);
nor U17313 (N_17313,N_16891,N_16847);
xor U17314 (N_17314,N_16974,N_16968);
and U17315 (N_17315,N_17075,N_17054);
nand U17316 (N_17316,N_16997,N_16988);
and U17317 (N_17317,N_16843,N_17063);
and U17318 (N_17318,N_17007,N_16962);
nor U17319 (N_17319,N_17022,N_16987);
and U17320 (N_17320,N_17051,N_16959);
nor U17321 (N_17321,N_17016,N_17057);
nand U17322 (N_17322,N_17024,N_17086);
xnor U17323 (N_17323,N_16804,N_16903);
or U17324 (N_17324,N_16816,N_16849);
nand U17325 (N_17325,N_16882,N_17075);
nor U17326 (N_17326,N_17093,N_16847);
or U17327 (N_17327,N_16992,N_16817);
nand U17328 (N_17328,N_17070,N_16886);
and U17329 (N_17329,N_17036,N_16946);
nor U17330 (N_17330,N_16833,N_17088);
xor U17331 (N_17331,N_16830,N_16882);
or U17332 (N_17332,N_16819,N_17062);
and U17333 (N_17333,N_17049,N_16943);
nor U17334 (N_17334,N_17052,N_16881);
nor U17335 (N_17335,N_16829,N_16823);
xor U17336 (N_17336,N_16901,N_16957);
or U17337 (N_17337,N_16865,N_17099);
nor U17338 (N_17338,N_16972,N_17065);
nor U17339 (N_17339,N_17064,N_16938);
nand U17340 (N_17340,N_16854,N_16855);
nor U17341 (N_17341,N_17068,N_16829);
or U17342 (N_17342,N_16939,N_17044);
nand U17343 (N_17343,N_17083,N_17059);
and U17344 (N_17344,N_16858,N_16840);
or U17345 (N_17345,N_17001,N_16823);
and U17346 (N_17346,N_16933,N_17032);
or U17347 (N_17347,N_16984,N_17075);
nor U17348 (N_17348,N_16900,N_16985);
xor U17349 (N_17349,N_16859,N_16976);
or U17350 (N_17350,N_16999,N_16899);
and U17351 (N_17351,N_16806,N_16843);
nand U17352 (N_17352,N_16850,N_16803);
or U17353 (N_17353,N_17005,N_16816);
and U17354 (N_17354,N_16887,N_17040);
nand U17355 (N_17355,N_16901,N_16818);
xor U17356 (N_17356,N_16928,N_17084);
or U17357 (N_17357,N_16845,N_16945);
and U17358 (N_17358,N_17039,N_17048);
nor U17359 (N_17359,N_16904,N_17056);
and U17360 (N_17360,N_17044,N_16936);
nor U17361 (N_17361,N_17098,N_17085);
or U17362 (N_17362,N_16820,N_16814);
or U17363 (N_17363,N_17092,N_16966);
nand U17364 (N_17364,N_17070,N_16819);
nand U17365 (N_17365,N_16904,N_16927);
xor U17366 (N_17366,N_16902,N_16885);
or U17367 (N_17367,N_16883,N_17019);
or U17368 (N_17368,N_16987,N_17043);
nor U17369 (N_17369,N_16834,N_16976);
nor U17370 (N_17370,N_17017,N_16957);
xor U17371 (N_17371,N_16818,N_17049);
xnor U17372 (N_17372,N_16856,N_16885);
and U17373 (N_17373,N_17001,N_17054);
xor U17374 (N_17374,N_16822,N_17066);
nor U17375 (N_17375,N_16815,N_16985);
or U17376 (N_17376,N_17037,N_16946);
xor U17377 (N_17377,N_16844,N_16941);
and U17378 (N_17378,N_17014,N_17015);
xor U17379 (N_17379,N_16884,N_17023);
nor U17380 (N_17380,N_16926,N_16809);
nand U17381 (N_17381,N_17010,N_16921);
xnor U17382 (N_17382,N_16971,N_16803);
and U17383 (N_17383,N_16899,N_16939);
or U17384 (N_17384,N_17055,N_16930);
xnor U17385 (N_17385,N_16871,N_16973);
and U17386 (N_17386,N_16993,N_16861);
xor U17387 (N_17387,N_17040,N_16840);
xor U17388 (N_17388,N_16971,N_16874);
or U17389 (N_17389,N_17060,N_16813);
nand U17390 (N_17390,N_16803,N_17026);
nand U17391 (N_17391,N_17049,N_16813);
nor U17392 (N_17392,N_16926,N_16931);
and U17393 (N_17393,N_16828,N_16924);
nand U17394 (N_17394,N_16836,N_17048);
nand U17395 (N_17395,N_16915,N_17011);
xor U17396 (N_17396,N_16926,N_16839);
and U17397 (N_17397,N_17045,N_16850);
and U17398 (N_17398,N_16987,N_16908);
xor U17399 (N_17399,N_16937,N_16814);
and U17400 (N_17400,N_17379,N_17187);
or U17401 (N_17401,N_17256,N_17137);
nor U17402 (N_17402,N_17126,N_17165);
or U17403 (N_17403,N_17396,N_17291);
and U17404 (N_17404,N_17221,N_17166);
nor U17405 (N_17405,N_17283,N_17348);
nand U17406 (N_17406,N_17334,N_17275);
or U17407 (N_17407,N_17131,N_17344);
nor U17408 (N_17408,N_17229,N_17257);
and U17409 (N_17409,N_17101,N_17398);
or U17410 (N_17410,N_17176,N_17231);
nor U17411 (N_17411,N_17173,N_17282);
nor U17412 (N_17412,N_17136,N_17163);
xor U17413 (N_17413,N_17203,N_17274);
xnor U17414 (N_17414,N_17251,N_17271);
nand U17415 (N_17415,N_17337,N_17242);
and U17416 (N_17416,N_17252,N_17366);
nor U17417 (N_17417,N_17304,N_17299);
and U17418 (N_17418,N_17360,N_17389);
nor U17419 (N_17419,N_17109,N_17182);
xnor U17420 (N_17420,N_17189,N_17354);
nor U17421 (N_17421,N_17152,N_17111);
or U17422 (N_17422,N_17106,N_17273);
nand U17423 (N_17423,N_17172,N_17325);
or U17424 (N_17424,N_17116,N_17162);
or U17425 (N_17425,N_17292,N_17356);
or U17426 (N_17426,N_17365,N_17159);
and U17427 (N_17427,N_17142,N_17193);
xnor U17428 (N_17428,N_17324,N_17160);
or U17429 (N_17429,N_17175,N_17181);
xnor U17430 (N_17430,N_17248,N_17349);
nand U17431 (N_17431,N_17154,N_17388);
nand U17432 (N_17432,N_17371,N_17297);
xnor U17433 (N_17433,N_17140,N_17335);
and U17434 (N_17434,N_17112,N_17372);
or U17435 (N_17435,N_17276,N_17293);
xor U17436 (N_17436,N_17202,N_17121);
and U17437 (N_17437,N_17170,N_17208);
nand U17438 (N_17438,N_17153,N_17183);
nor U17439 (N_17439,N_17262,N_17359);
xor U17440 (N_17440,N_17345,N_17213);
or U17441 (N_17441,N_17215,N_17322);
xor U17442 (N_17442,N_17307,N_17122);
or U17443 (N_17443,N_17373,N_17285);
xor U17444 (N_17444,N_17341,N_17155);
xnor U17445 (N_17445,N_17323,N_17386);
nor U17446 (N_17446,N_17377,N_17331);
and U17447 (N_17447,N_17279,N_17357);
nor U17448 (N_17448,N_17258,N_17261);
xnor U17449 (N_17449,N_17178,N_17117);
or U17450 (N_17450,N_17199,N_17194);
or U17451 (N_17451,N_17306,N_17198);
xnor U17452 (N_17452,N_17316,N_17287);
and U17453 (N_17453,N_17151,N_17267);
nor U17454 (N_17454,N_17222,N_17207);
nand U17455 (N_17455,N_17336,N_17281);
xnor U17456 (N_17456,N_17192,N_17133);
nor U17457 (N_17457,N_17353,N_17288);
xor U17458 (N_17458,N_17327,N_17171);
nor U17459 (N_17459,N_17216,N_17168);
nand U17460 (N_17460,N_17390,N_17370);
nor U17461 (N_17461,N_17232,N_17135);
nor U17462 (N_17462,N_17141,N_17150);
nand U17463 (N_17463,N_17332,N_17329);
and U17464 (N_17464,N_17104,N_17362);
nand U17465 (N_17465,N_17355,N_17394);
nand U17466 (N_17466,N_17119,N_17266);
and U17467 (N_17467,N_17378,N_17164);
and U17468 (N_17468,N_17149,N_17290);
and U17469 (N_17469,N_17308,N_17206);
xnor U17470 (N_17470,N_17108,N_17161);
nand U17471 (N_17471,N_17205,N_17220);
or U17472 (N_17472,N_17384,N_17103);
or U17473 (N_17473,N_17277,N_17300);
xor U17474 (N_17474,N_17338,N_17144);
nor U17475 (N_17475,N_17265,N_17247);
and U17476 (N_17476,N_17115,N_17369);
nand U17477 (N_17477,N_17139,N_17224);
nor U17478 (N_17478,N_17328,N_17201);
xnor U17479 (N_17479,N_17387,N_17125);
and U17480 (N_17480,N_17367,N_17295);
nand U17481 (N_17481,N_17185,N_17312);
nor U17482 (N_17482,N_17114,N_17110);
nand U17483 (N_17483,N_17228,N_17249);
or U17484 (N_17484,N_17120,N_17393);
nand U17485 (N_17485,N_17167,N_17234);
nor U17486 (N_17486,N_17330,N_17244);
nand U17487 (N_17487,N_17156,N_17204);
and U17488 (N_17488,N_17333,N_17280);
nor U17489 (N_17489,N_17347,N_17113);
xor U17490 (N_17490,N_17180,N_17218);
xnor U17491 (N_17491,N_17268,N_17399);
nor U17492 (N_17492,N_17264,N_17177);
nand U17493 (N_17493,N_17395,N_17246);
or U17494 (N_17494,N_17259,N_17303);
and U17495 (N_17495,N_17364,N_17385);
nand U17496 (N_17496,N_17239,N_17250);
nand U17497 (N_17497,N_17255,N_17343);
nor U17498 (N_17498,N_17269,N_17100);
and U17499 (N_17499,N_17241,N_17313);
or U17500 (N_17500,N_17105,N_17315);
xnor U17501 (N_17501,N_17107,N_17186);
nand U17502 (N_17502,N_17226,N_17191);
nor U17503 (N_17503,N_17146,N_17236);
nand U17504 (N_17504,N_17294,N_17227);
nand U17505 (N_17505,N_17169,N_17289);
or U17506 (N_17506,N_17158,N_17254);
and U17507 (N_17507,N_17301,N_17240);
or U17508 (N_17508,N_17129,N_17284);
and U17509 (N_17509,N_17342,N_17319);
nor U17510 (N_17510,N_17363,N_17147);
and U17511 (N_17511,N_17223,N_17298);
nand U17512 (N_17512,N_17296,N_17217);
nor U17513 (N_17513,N_17358,N_17381);
xnor U17514 (N_17514,N_17368,N_17188);
nor U17515 (N_17515,N_17143,N_17130);
and U17516 (N_17516,N_17253,N_17145);
xor U17517 (N_17517,N_17243,N_17124);
or U17518 (N_17518,N_17317,N_17380);
xnor U17519 (N_17519,N_17397,N_17238);
and U17520 (N_17520,N_17179,N_17174);
nor U17521 (N_17521,N_17157,N_17361);
or U17522 (N_17522,N_17235,N_17326);
and U17523 (N_17523,N_17245,N_17272);
xor U17524 (N_17524,N_17102,N_17340);
and U17525 (N_17525,N_17318,N_17196);
nand U17526 (N_17526,N_17233,N_17270);
xnor U17527 (N_17527,N_17138,N_17128);
xor U17528 (N_17528,N_17383,N_17350);
nand U17529 (N_17529,N_17184,N_17392);
nand U17530 (N_17530,N_17123,N_17352);
nand U17531 (N_17531,N_17339,N_17260);
xnor U17532 (N_17532,N_17375,N_17210);
or U17533 (N_17533,N_17209,N_17219);
xnor U17534 (N_17534,N_17230,N_17197);
and U17535 (N_17535,N_17382,N_17346);
xor U17536 (N_17536,N_17314,N_17225);
nor U17537 (N_17537,N_17351,N_17214);
nand U17538 (N_17538,N_17200,N_17321);
nand U17539 (N_17539,N_17134,N_17278);
or U17540 (N_17540,N_17305,N_17309);
xor U17541 (N_17541,N_17118,N_17376);
xor U17542 (N_17542,N_17263,N_17132);
xnor U17543 (N_17543,N_17302,N_17195);
nand U17544 (N_17544,N_17310,N_17212);
or U17545 (N_17545,N_17190,N_17127);
nor U17546 (N_17546,N_17374,N_17211);
and U17547 (N_17547,N_17391,N_17320);
and U17548 (N_17548,N_17148,N_17311);
nand U17549 (N_17549,N_17286,N_17237);
xor U17550 (N_17550,N_17353,N_17376);
xnor U17551 (N_17551,N_17237,N_17202);
or U17552 (N_17552,N_17281,N_17160);
or U17553 (N_17553,N_17268,N_17356);
nor U17554 (N_17554,N_17321,N_17281);
xnor U17555 (N_17555,N_17147,N_17109);
nor U17556 (N_17556,N_17331,N_17359);
and U17557 (N_17557,N_17165,N_17142);
nor U17558 (N_17558,N_17350,N_17368);
and U17559 (N_17559,N_17226,N_17319);
and U17560 (N_17560,N_17343,N_17396);
nand U17561 (N_17561,N_17113,N_17245);
or U17562 (N_17562,N_17105,N_17308);
and U17563 (N_17563,N_17391,N_17353);
nor U17564 (N_17564,N_17114,N_17334);
and U17565 (N_17565,N_17307,N_17117);
and U17566 (N_17566,N_17235,N_17362);
nor U17567 (N_17567,N_17156,N_17265);
or U17568 (N_17568,N_17311,N_17342);
or U17569 (N_17569,N_17219,N_17261);
nand U17570 (N_17570,N_17128,N_17311);
nand U17571 (N_17571,N_17283,N_17344);
nand U17572 (N_17572,N_17160,N_17144);
or U17573 (N_17573,N_17306,N_17192);
and U17574 (N_17574,N_17288,N_17333);
nor U17575 (N_17575,N_17376,N_17339);
or U17576 (N_17576,N_17306,N_17174);
and U17577 (N_17577,N_17360,N_17290);
and U17578 (N_17578,N_17160,N_17176);
nand U17579 (N_17579,N_17217,N_17183);
nor U17580 (N_17580,N_17137,N_17261);
and U17581 (N_17581,N_17363,N_17103);
or U17582 (N_17582,N_17189,N_17231);
and U17583 (N_17583,N_17359,N_17115);
xnor U17584 (N_17584,N_17254,N_17189);
nand U17585 (N_17585,N_17134,N_17156);
or U17586 (N_17586,N_17397,N_17242);
and U17587 (N_17587,N_17280,N_17390);
nor U17588 (N_17588,N_17321,N_17363);
or U17589 (N_17589,N_17132,N_17136);
xnor U17590 (N_17590,N_17233,N_17134);
and U17591 (N_17591,N_17397,N_17312);
or U17592 (N_17592,N_17378,N_17318);
nand U17593 (N_17593,N_17253,N_17396);
and U17594 (N_17594,N_17363,N_17168);
nand U17595 (N_17595,N_17125,N_17392);
nor U17596 (N_17596,N_17181,N_17362);
xor U17597 (N_17597,N_17233,N_17302);
nor U17598 (N_17598,N_17257,N_17125);
or U17599 (N_17599,N_17380,N_17195);
or U17600 (N_17600,N_17105,N_17397);
nand U17601 (N_17601,N_17135,N_17109);
xnor U17602 (N_17602,N_17376,N_17236);
nor U17603 (N_17603,N_17268,N_17305);
and U17604 (N_17604,N_17332,N_17142);
nand U17605 (N_17605,N_17289,N_17286);
xor U17606 (N_17606,N_17170,N_17346);
nor U17607 (N_17607,N_17123,N_17385);
nor U17608 (N_17608,N_17295,N_17233);
and U17609 (N_17609,N_17118,N_17101);
xnor U17610 (N_17610,N_17325,N_17306);
or U17611 (N_17611,N_17120,N_17340);
and U17612 (N_17612,N_17135,N_17220);
xnor U17613 (N_17613,N_17385,N_17326);
xor U17614 (N_17614,N_17100,N_17217);
and U17615 (N_17615,N_17344,N_17258);
nor U17616 (N_17616,N_17237,N_17290);
or U17617 (N_17617,N_17233,N_17279);
or U17618 (N_17618,N_17126,N_17192);
and U17619 (N_17619,N_17386,N_17103);
nor U17620 (N_17620,N_17156,N_17270);
and U17621 (N_17621,N_17180,N_17187);
nor U17622 (N_17622,N_17328,N_17264);
or U17623 (N_17623,N_17341,N_17154);
and U17624 (N_17624,N_17245,N_17343);
nor U17625 (N_17625,N_17347,N_17262);
xnor U17626 (N_17626,N_17311,N_17210);
or U17627 (N_17627,N_17261,N_17279);
xnor U17628 (N_17628,N_17368,N_17121);
nand U17629 (N_17629,N_17110,N_17330);
nand U17630 (N_17630,N_17139,N_17156);
or U17631 (N_17631,N_17168,N_17166);
xnor U17632 (N_17632,N_17103,N_17145);
or U17633 (N_17633,N_17359,N_17231);
xor U17634 (N_17634,N_17383,N_17254);
xnor U17635 (N_17635,N_17189,N_17210);
and U17636 (N_17636,N_17349,N_17337);
nand U17637 (N_17637,N_17367,N_17160);
xnor U17638 (N_17638,N_17113,N_17243);
and U17639 (N_17639,N_17304,N_17378);
nand U17640 (N_17640,N_17330,N_17289);
xor U17641 (N_17641,N_17142,N_17190);
or U17642 (N_17642,N_17115,N_17188);
or U17643 (N_17643,N_17328,N_17185);
and U17644 (N_17644,N_17265,N_17196);
and U17645 (N_17645,N_17103,N_17317);
nor U17646 (N_17646,N_17155,N_17359);
nand U17647 (N_17647,N_17153,N_17161);
or U17648 (N_17648,N_17368,N_17237);
or U17649 (N_17649,N_17386,N_17204);
nand U17650 (N_17650,N_17188,N_17133);
nor U17651 (N_17651,N_17200,N_17272);
and U17652 (N_17652,N_17305,N_17380);
and U17653 (N_17653,N_17261,N_17349);
or U17654 (N_17654,N_17382,N_17185);
nor U17655 (N_17655,N_17294,N_17308);
xnor U17656 (N_17656,N_17313,N_17168);
or U17657 (N_17657,N_17280,N_17350);
nor U17658 (N_17658,N_17301,N_17179);
nor U17659 (N_17659,N_17274,N_17334);
nand U17660 (N_17660,N_17131,N_17386);
nor U17661 (N_17661,N_17269,N_17202);
nand U17662 (N_17662,N_17304,N_17139);
nand U17663 (N_17663,N_17129,N_17193);
xor U17664 (N_17664,N_17307,N_17184);
xor U17665 (N_17665,N_17192,N_17100);
nand U17666 (N_17666,N_17242,N_17188);
nor U17667 (N_17667,N_17173,N_17116);
nor U17668 (N_17668,N_17121,N_17181);
or U17669 (N_17669,N_17125,N_17190);
nand U17670 (N_17670,N_17351,N_17131);
nor U17671 (N_17671,N_17212,N_17369);
or U17672 (N_17672,N_17229,N_17238);
or U17673 (N_17673,N_17315,N_17200);
nor U17674 (N_17674,N_17398,N_17333);
xnor U17675 (N_17675,N_17131,N_17396);
nand U17676 (N_17676,N_17249,N_17126);
or U17677 (N_17677,N_17344,N_17391);
or U17678 (N_17678,N_17168,N_17129);
and U17679 (N_17679,N_17385,N_17304);
or U17680 (N_17680,N_17316,N_17170);
and U17681 (N_17681,N_17222,N_17111);
xnor U17682 (N_17682,N_17243,N_17151);
xor U17683 (N_17683,N_17153,N_17252);
or U17684 (N_17684,N_17355,N_17298);
nand U17685 (N_17685,N_17320,N_17380);
nand U17686 (N_17686,N_17297,N_17128);
nor U17687 (N_17687,N_17384,N_17126);
xnor U17688 (N_17688,N_17138,N_17153);
nor U17689 (N_17689,N_17299,N_17177);
or U17690 (N_17690,N_17319,N_17356);
or U17691 (N_17691,N_17372,N_17211);
and U17692 (N_17692,N_17168,N_17126);
or U17693 (N_17693,N_17345,N_17283);
nand U17694 (N_17694,N_17160,N_17161);
nor U17695 (N_17695,N_17138,N_17270);
nor U17696 (N_17696,N_17312,N_17290);
nor U17697 (N_17697,N_17334,N_17248);
nand U17698 (N_17698,N_17396,N_17135);
xor U17699 (N_17699,N_17344,N_17292);
xnor U17700 (N_17700,N_17499,N_17581);
nand U17701 (N_17701,N_17539,N_17505);
xnor U17702 (N_17702,N_17532,N_17682);
nor U17703 (N_17703,N_17409,N_17444);
or U17704 (N_17704,N_17578,N_17625);
nor U17705 (N_17705,N_17549,N_17420);
or U17706 (N_17706,N_17551,N_17494);
nor U17707 (N_17707,N_17543,N_17589);
xnor U17708 (N_17708,N_17656,N_17611);
and U17709 (N_17709,N_17662,N_17458);
nand U17710 (N_17710,N_17452,N_17677);
or U17711 (N_17711,N_17429,N_17674);
xnor U17712 (N_17712,N_17546,N_17424);
and U17713 (N_17713,N_17561,N_17618);
or U17714 (N_17714,N_17473,N_17520);
nand U17715 (N_17715,N_17435,N_17482);
and U17716 (N_17716,N_17560,N_17684);
xor U17717 (N_17717,N_17547,N_17580);
nand U17718 (N_17718,N_17640,N_17510);
and U17719 (N_17719,N_17531,N_17615);
nor U17720 (N_17720,N_17418,N_17571);
or U17721 (N_17721,N_17408,N_17471);
nand U17722 (N_17722,N_17638,N_17526);
nand U17723 (N_17723,N_17699,N_17462);
and U17724 (N_17724,N_17566,N_17517);
nor U17725 (N_17725,N_17565,N_17481);
and U17726 (N_17726,N_17415,N_17590);
or U17727 (N_17727,N_17600,N_17417);
or U17728 (N_17728,N_17502,N_17465);
nor U17729 (N_17729,N_17649,N_17511);
nor U17730 (N_17730,N_17513,N_17689);
nand U17731 (N_17731,N_17617,N_17425);
nand U17732 (N_17732,N_17515,N_17642);
xor U17733 (N_17733,N_17688,N_17599);
xor U17734 (N_17734,N_17533,N_17512);
or U17735 (N_17735,N_17574,N_17623);
or U17736 (N_17736,N_17664,N_17667);
and U17737 (N_17737,N_17647,N_17440);
xnor U17738 (N_17738,N_17643,N_17498);
xnor U17739 (N_17739,N_17427,N_17404);
and U17740 (N_17740,N_17562,N_17636);
or U17741 (N_17741,N_17423,N_17443);
or U17742 (N_17742,N_17654,N_17609);
or U17743 (N_17743,N_17619,N_17605);
and U17744 (N_17744,N_17448,N_17493);
nand U17745 (N_17745,N_17601,N_17430);
nand U17746 (N_17746,N_17535,N_17434);
and U17747 (N_17747,N_17610,N_17504);
and U17748 (N_17748,N_17530,N_17495);
xor U17749 (N_17749,N_17472,N_17541);
or U17750 (N_17750,N_17613,N_17529);
and U17751 (N_17751,N_17487,N_17478);
nand U17752 (N_17752,N_17542,N_17419);
nor U17753 (N_17753,N_17557,N_17540);
and U17754 (N_17754,N_17608,N_17407);
xnor U17755 (N_17755,N_17606,N_17519);
nand U17756 (N_17756,N_17413,N_17428);
nand U17757 (N_17757,N_17631,N_17657);
or U17758 (N_17758,N_17678,N_17676);
nor U17759 (N_17759,N_17421,N_17523);
xor U17760 (N_17760,N_17690,N_17594);
and U17761 (N_17761,N_17641,N_17485);
nand U17762 (N_17762,N_17463,N_17506);
nand U17763 (N_17763,N_17476,N_17414);
xnor U17764 (N_17764,N_17460,N_17441);
xor U17765 (N_17765,N_17489,N_17537);
nor U17766 (N_17766,N_17470,N_17445);
nand U17767 (N_17767,N_17544,N_17439);
or U17768 (N_17768,N_17572,N_17669);
or U17769 (N_17769,N_17450,N_17595);
xor U17770 (N_17770,N_17570,N_17621);
nand U17771 (N_17771,N_17469,N_17692);
nand U17772 (N_17772,N_17576,N_17545);
nand U17773 (N_17773,N_17693,N_17695);
xor U17774 (N_17774,N_17401,N_17436);
nand U17775 (N_17775,N_17516,N_17646);
nand U17776 (N_17776,N_17490,N_17593);
xor U17777 (N_17777,N_17671,N_17672);
nor U17778 (N_17778,N_17488,N_17582);
and U17779 (N_17779,N_17412,N_17586);
xnor U17780 (N_17780,N_17597,N_17585);
and U17781 (N_17781,N_17538,N_17588);
or U17782 (N_17782,N_17634,N_17534);
nand U17783 (N_17783,N_17496,N_17563);
xnor U17784 (N_17784,N_17577,N_17607);
and U17785 (N_17785,N_17624,N_17675);
or U17786 (N_17786,N_17698,N_17591);
or U17787 (N_17787,N_17518,N_17637);
nand U17788 (N_17788,N_17666,N_17527);
nand U17789 (N_17789,N_17468,N_17645);
nor U17790 (N_17790,N_17522,N_17620);
nor U17791 (N_17791,N_17602,N_17457);
or U17792 (N_17792,N_17426,N_17622);
and U17793 (N_17793,N_17652,N_17697);
nor U17794 (N_17794,N_17558,N_17564);
xor U17795 (N_17795,N_17668,N_17616);
nor U17796 (N_17796,N_17449,N_17579);
xor U17797 (N_17797,N_17648,N_17501);
nor U17798 (N_17798,N_17480,N_17670);
or U17799 (N_17799,N_17453,N_17681);
nor U17800 (N_17800,N_17524,N_17486);
xnor U17801 (N_17801,N_17442,N_17644);
or U17802 (N_17802,N_17630,N_17660);
nand U17803 (N_17803,N_17567,N_17687);
xor U17804 (N_17804,N_17403,N_17653);
nand U17805 (N_17805,N_17658,N_17604);
nor U17806 (N_17806,N_17691,N_17433);
or U17807 (N_17807,N_17573,N_17402);
nor U17808 (N_17808,N_17603,N_17628);
or U17809 (N_17809,N_17437,N_17556);
and U17810 (N_17810,N_17497,N_17492);
or U17811 (N_17811,N_17614,N_17612);
nand U17812 (N_17812,N_17466,N_17467);
and U17813 (N_17813,N_17528,N_17694);
and U17814 (N_17814,N_17451,N_17559);
xnor U17815 (N_17815,N_17659,N_17665);
xnor U17816 (N_17816,N_17679,N_17553);
xor U17817 (N_17817,N_17596,N_17632);
and U17818 (N_17818,N_17410,N_17555);
nor U17819 (N_17819,N_17598,N_17406);
or U17820 (N_17820,N_17456,N_17461);
nor U17821 (N_17821,N_17509,N_17474);
or U17822 (N_17822,N_17483,N_17548);
nand U17823 (N_17823,N_17491,N_17507);
and U17824 (N_17824,N_17680,N_17626);
and U17825 (N_17825,N_17447,N_17454);
xor U17826 (N_17826,N_17411,N_17400);
nand U17827 (N_17827,N_17477,N_17405);
or U17828 (N_17828,N_17629,N_17661);
or U17829 (N_17829,N_17432,N_17696);
and U17830 (N_17830,N_17569,N_17633);
and U17831 (N_17831,N_17416,N_17650);
and U17832 (N_17832,N_17627,N_17639);
xnor U17833 (N_17833,N_17484,N_17431);
and U17834 (N_17834,N_17655,N_17673);
xor U17835 (N_17835,N_17446,N_17651);
nand U17836 (N_17836,N_17584,N_17475);
nor U17837 (N_17837,N_17554,N_17686);
xnor U17838 (N_17838,N_17514,N_17568);
nand U17839 (N_17839,N_17592,N_17583);
or U17840 (N_17840,N_17479,N_17500);
and U17841 (N_17841,N_17459,N_17503);
nor U17842 (N_17842,N_17508,N_17525);
xnor U17843 (N_17843,N_17635,N_17575);
xnor U17844 (N_17844,N_17683,N_17685);
nor U17845 (N_17845,N_17550,N_17521);
nand U17846 (N_17846,N_17536,N_17587);
nand U17847 (N_17847,N_17438,N_17464);
or U17848 (N_17848,N_17663,N_17422);
and U17849 (N_17849,N_17455,N_17552);
nand U17850 (N_17850,N_17472,N_17407);
nand U17851 (N_17851,N_17690,N_17505);
nor U17852 (N_17852,N_17419,N_17579);
xor U17853 (N_17853,N_17571,N_17608);
nand U17854 (N_17854,N_17402,N_17605);
nand U17855 (N_17855,N_17524,N_17630);
nand U17856 (N_17856,N_17646,N_17436);
nor U17857 (N_17857,N_17692,N_17517);
nand U17858 (N_17858,N_17554,N_17438);
or U17859 (N_17859,N_17452,N_17675);
and U17860 (N_17860,N_17623,N_17567);
nand U17861 (N_17861,N_17491,N_17495);
nand U17862 (N_17862,N_17477,N_17683);
or U17863 (N_17863,N_17576,N_17409);
nor U17864 (N_17864,N_17497,N_17548);
nand U17865 (N_17865,N_17679,N_17549);
nand U17866 (N_17866,N_17547,N_17674);
or U17867 (N_17867,N_17675,N_17605);
nand U17868 (N_17868,N_17547,N_17530);
xnor U17869 (N_17869,N_17651,N_17537);
nand U17870 (N_17870,N_17409,N_17453);
xor U17871 (N_17871,N_17423,N_17450);
and U17872 (N_17872,N_17674,N_17616);
nand U17873 (N_17873,N_17450,N_17410);
nand U17874 (N_17874,N_17416,N_17434);
xnor U17875 (N_17875,N_17682,N_17668);
xnor U17876 (N_17876,N_17694,N_17557);
nand U17877 (N_17877,N_17443,N_17664);
or U17878 (N_17878,N_17535,N_17496);
xnor U17879 (N_17879,N_17653,N_17587);
xor U17880 (N_17880,N_17455,N_17472);
nor U17881 (N_17881,N_17570,N_17470);
xor U17882 (N_17882,N_17408,N_17426);
and U17883 (N_17883,N_17626,N_17490);
nand U17884 (N_17884,N_17603,N_17520);
and U17885 (N_17885,N_17406,N_17658);
or U17886 (N_17886,N_17619,N_17423);
nor U17887 (N_17887,N_17582,N_17591);
or U17888 (N_17888,N_17562,N_17651);
and U17889 (N_17889,N_17474,N_17451);
and U17890 (N_17890,N_17578,N_17512);
nor U17891 (N_17891,N_17643,N_17591);
or U17892 (N_17892,N_17469,N_17648);
nor U17893 (N_17893,N_17545,N_17525);
nor U17894 (N_17894,N_17627,N_17689);
nand U17895 (N_17895,N_17623,N_17558);
and U17896 (N_17896,N_17462,N_17645);
nor U17897 (N_17897,N_17611,N_17466);
or U17898 (N_17898,N_17626,N_17497);
or U17899 (N_17899,N_17599,N_17524);
or U17900 (N_17900,N_17410,N_17537);
xnor U17901 (N_17901,N_17667,N_17643);
nor U17902 (N_17902,N_17423,N_17593);
nand U17903 (N_17903,N_17488,N_17494);
nor U17904 (N_17904,N_17498,N_17457);
xnor U17905 (N_17905,N_17574,N_17612);
nor U17906 (N_17906,N_17690,N_17589);
xor U17907 (N_17907,N_17421,N_17605);
or U17908 (N_17908,N_17401,N_17482);
nor U17909 (N_17909,N_17505,N_17454);
and U17910 (N_17910,N_17678,N_17664);
nand U17911 (N_17911,N_17445,N_17474);
nor U17912 (N_17912,N_17414,N_17409);
nand U17913 (N_17913,N_17653,N_17636);
or U17914 (N_17914,N_17528,N_17495);
nor U17915 (N_17915,N_17580,N_17437);
and U17916 (N_17916,N_17436,N_17644);
xor U17917 (N_17917,N_17639,N_17506);
nor U17918 (N_17918,N_17548,N_17441);
xor U17919 (N_17919,N_17674,N_17627);
xor U17920 (N_17920,N_17548,N_17613);
nor U17921 (N_17921,N_17588,N_17515);
nor U17922 (N_17922,N_17436,N_17675);
and U17923 (N_17923,N_17489,N_17599);
nor U17924 (N_17924,N_17591,N_17431);
nand U17925 (N_17925,N_17579,N_17586);
and U17926 (N_17926,N_17553,N_17650);
nor U17927 (N_17927,N_17649,N_17643);
and U17928 (N_17928,N_17401,N_17554);
and U17929 (N_17929,N_17539,N_17603);
nand U17930 (N_17930,N_17628,N_17626);
nand U17931 (N_17931,N_17593,N_17506);
nand U17932 (N_17932,N_17529,N_17567);
and U17933 (N_17933,N_17682,N_17579);
and U17934 (N_17934,N_17535,N_17407);
and U17935 (N_17935,N_17570,N_17614);
xnor U17936 (N_17936,N_17425,N_17630);
or U17937 (N_17937,N_17499,N_17626);
nor U17938 (N_17938,N_17560,N_17429);
or U17939 (N_17939,N_17534,N_17691);
xor U17940 (N_17940,N_17513,N_17571);
xnor U17941 (N_17941,N_17634,N_17424);
nor U17942 (N_17942,N_17450,N_17427);
nand U17943 (N_17943,N_17642,N_17545);
and U17944 (N_17944,N_17523,N_17429);
xnor U17945 (N_17945,N_17466,N_17482);
and U17946 (N_17946,N_17541,N_17558);
or U17947 (N_17947,N_17676,N_17503);
nor U17948 (N_17948,N_17678,N_17493);
nor U17949 (N_17949,N_17660,N_17676);
xnor U17950 (N_17950,N_17645,N_17413);
or U17951 (N_17951,N_17458,N_17486);
nand U17952 (N_17952,N_17693,N_17473);
and U17953 (N_17953,N_17652,N_17545);
nand U17954 (N_17954,N_17418,N_17433);
xnor U17955 (N_17955,N_17674,N_17457);
xor U17956 (N_17956,N_17508,N_17491);
nand U17957 (N_17957,N_17562,N_17576);
and U17958 (N_17958,N_17525,N_17685);
xnor U17959 (N_17959,N_17581,N_17451);
or U17960 (N_17960,N_17567,N_17579);
nor U17961 (N_17961,N_17492,N_17692);
and U17962 (N_17962,N_17591,N_17473);
nand U17963 (N_17963,N_17608,N_17406);
xor U17964 (N_17964,N_17563,N_17474);
and U17965 (N_17965,N_17572,N_17515);
xnor U17966 (N_17966,N_17477,N_17565);
and U17967 (N_17967,N_17429,N_17402);
xor U17968 (N_17968,N_17408,N_17431);
or U17969 (N_17969,N_17617,N_17606);
or U17970 (N_17970,N_17551,N_17689);
xor U17971 (N_17971,N_17491,N_17575);
nand U17972 (N_17972,N_17490,N_17574);
xor U17973 (N_17973,N_17432,N_17491);
xor U17974 (N_17974,N_17599,N_17689);
or U17975 (N_17975,N_17450,N_17506);
or U17976 (N_17976,N_17572,N_17453);
and U17977 (N_17977,N_17603,N_17413);
and U17978 (N_17978,N_17670,N_17428);
and U17979 (N_17979,N_17486,N_17589);
nand U17980 (N_17980,N_17451,N_17692);
xor U17981 (N_17981,N_17466,N_17699);
nor U17982 (N_17982,N_17489,N_17487);
and U17983 (N_17983,N_17495,N_17526);
or U17984 (N_17984,N_17443,N_17616);
and U17985 (N_17985,N_17444,N_17668);
xor U17986 (N_17986,N_17543,N_17537);
xor U17987 (N_17987,N_17680,N_17421);
nand U17988 (N_17988,N_17695,N_17467);
xnor U17989 (N_17989,N_17691,N_17407);
nor U17990 (N_17990,N_17472,N_17631);
nand U17991 (N_17991,N_17440,N_17536);
and U17992 (N_17992,N_17625,N_17471);
nand U17993 (N_17993,N_17550,N_17537);
nand U17994 (N_17994,N_17410,N_17575);
nor U17995 (N_17995,N_17579,N_17613);
xnor U17996 (N_17996,N_17639,N_17637);
and U17997 (N_17997,N_17630,N_17522);
xor U17998 (N_17998,N_17502,N_17423);
or U17999 (N_17999,N_17434,N_17610);
nand U18000 (N_18000,N_17749,N_17704);
nand U18001 (N_18001,N_17725,N_17939);
and U18002 (N_18002,N_17879,N_17733);
nor U18003 (N_18003,N_17887,N_17950);
and U18004 (N_18004,N_17884,N_17730);
xor U18005 (N_18005,N_17721,N_17997);
nand U18006 (N_18006,N_17754,N_17738);
nand U18007 (N_18007,N_17974,N_17720);
xor U18008 (N_18008,N_17750,N_17760);
or U18009 (N_18009,N_17813,N_17954);
or U18010 (N_18010,N_17827,N_17743);
xnor U18011 (N_18011,N_17739,N_17755);
nand U18012 (N_18012,N_17967,N_17800);
or U18013 (N_18013,N_17716,N_17710);
and U18014 (N_18014,N_17870,N_17834);
nor U18015 (N_18015,N_17938,N_17971);
xnor U18016 (N_18016,N_17890,N_17751);
nand U18017 (N_18017,N_17776,N_17968);
and U18018 (N_18018,N_17944,N_17972);
or U18019 (N_18019,N_17765,N_17898);
and U18020 (N_18020,N_17909,N_17708);
nor U18021 (N_18021,N_17881,N_17724);
nor U18022 (N_18022,N_17780,N_17839);
nand U18023 (N_18023,N_17978,N_17878);
or U18024 (N_18024,N_17953,N_17923);
and U18025 (N_18025,N_17844,N_17975);
and U18026 (N_18026,N_17863,N_17762);
xnor U18027 (N_18027,N_17703,N_17894);
nand U18028 (N_18028,N_17920,N_17719);
nor U18029 (N_18029,N_17828,N_17790);
xor U18030 (N_18030,N_17919,N_17701);
xnor U18031 (N_18031,N_17847,N_17940);
nand U18032 (N_18032,N_17767,N_17914);
nand U18033 (N_18033,N_17963,N_17857);
or U18034 (N_18034,N_17866,N_17726);
xor U18035 (N_18035,N_17900,N_17785);
or U18036 (N_18036,N_17883,N_17927);
and U18037 (N_18037,N_17849,N_17805);
xor U18038 (N_18038,N_17998,N_17711);
or U18039 (N_18039,N_17769,N_17921);
or U18040 (N_18040,N_17917,N_17826);
and U18041 (N_18041,N_17807,N_17753);
nand U18042 (N_18042,N_17862,N_17741);
nand U18043 (N_18043,N_17949,N_17740);
xor U18044 (N_18044,N_17875,N_17843);
xnor U18045 (N_18045,N_17745,N_17709);
or U18046 (N_18046,N_17775,N_17868);
or U18047 (N_18047,N_17951,N_17744);
nor U18048 (N_18048,N_17853,N_17845);
xor U18049 (N_18049,N_17908,N_17731);
nor U18050 (N_18050,N_17816,N_17803);
or U18051 (N_18051,N_17912,N_17988);
nand U18052 (N_18052,N_17916,N_17994);
nand U18053 (N_18053,N_17934,N_17903);
and U18054 (N_18054,N_17802,N_17722);
and U18055 (N_18055,N_17779,N_17999);
nand U18056 (N_18056,N_17865,N_17757);
nor U18057 (N_18057,N_17788,N_17764);
nand U18058 (N_18058,N_17990,N_17925);
nand U18059 (N_18059,N_17871,N_17985);
nand U18060 (N_18060,N_17861,N_17897);
nand U18061 (N_18061,N_17987,N_17929);
nor U18062 (N_18062,N_17906,N_17892);
and U18063 (N_18063,N_17713,N_17746);
and U18064 (N_18064,N_17918,N_17789);
xnor U18065 (N_18065,N_17854,N_17804);
nor U18066 (N_18066,N_17763,N_17822);
or U18067 (N_18067,N_17706,N_17993);
and U18068 (N_18068,N_17831,N_17941);
nor U18069 (N_18069,N_17984,N_17814);
and U18070 (N_18070,N_17809,N_17966);
and U18071 (N_18071,N_17806,N_17735);
and U18072 (N_18072,N_17889,N_17979);
or U18073 (N_18073,N_17957,N_17896);
nor U18074 (N_18074,N_17799,N_17820);
or U18075 (N_18075,N_17825,N_17756);
nand U18076 (N_18076,N_17782,N_17937);
nand U18077 (N_18077,N_17983,N_17742);
or U18078 (N_18078,N_17964,N_17946);
nand U18079 (N_18079,N_17715,N_17712);
xor U18080 (N_18080,N_17836,N_17833);
nor U18081 (N_18081,N_17933,N_17734);
nor U18082 (N_18082,N_17876,N_17787);
xnor U18083 (N_18083,N_17924,N_17702);
nor U18084 (N_18084,N_17996,N_17811);
nand U18085 (N_18085,N_17783,N_17856);
nand U18086 (N_18086,N_17960,N_17959);
nor U18087 (N_18087,N_17848,N_17815);
xor U18088 (N_18088,N_17705,N_17932);
and U18089 (N_18089,N_17913,N_17895);
xor U18090 (N_18090,N_17748,N_17723);
and U18091 (N_18091,N_17936,N_17922);
nor U18092 (N_18092,N_17948,N_17819);
or U18093 (N_18093,N_17801,N_17886);
or U18094 (N_18094,N_17714,N_17794);
xor U18095 (N_18095,N_17829,N_17880);
nor U18096 (N_18096,N_17995,N_17793);
xnor U18097 (N_18097,N_17882,N_17874);
nand U18098 (N_18098,N_17935,N_17942);
nand U18099 (N_18099,N_17774,N_17926);
or U18100 (N_18100,N_17791,N_17877);
and U18101 (N_18101,N_17947,N_17832);
and U18102 (N_18102,N_17817,N_17992);
and U18103 (N_18103,N_17777,N_17770);
and U18104 (N_18104,N_17928,N_17945);
and U18105 (N_18105,N_17905,N_17792);
and U18106 (N_18106,N_17980,N_17797);
nor U18107 (N_18107,N_17781,N_17812);
nor U18108 (N_18108,N_17773,N_17904);
nand U18109 (N_18109,N_17842,N_17956);
and U18110 (N_18110,N_17700,N_17747);
or U18111 (N_18111,N_17821,N_17810);
or U18112 (N_18112,N_17798,N_17915);
and U18113 (N_18113,N_17795,N_17717);
xnor U18114 (N_18114,N_17732,N_17893);
nand U18115 (N_18115,N_17952,N_17962);
nor U18116 (N_18116,N_17768,N_17867);
or U18117 (N_18117,N_17796,N_17986);
or U18118 (N_18118,N_17855,N_17977);
xor U18119 (N_18119,N_17728,N_17981);
and U18120 (N_18120,N_17784,N_17761);
and U18121 (N_18121,N_17902,N_17823);
and U18122 (N_18122,N_17888,N_17850);
and U18123 (N_18123,N_17846,N_17707);
or U18124 (N_18124,N_17737,N_17899);
or U18125 (N_18125,N_17965,N_17772);
nor U18126 (N_18126,N_17835,N_17958);
nor U18127 (N_18127,N_17869,N_17840);
nor U18128 (N_18128,N_17969,N_17837);
xnor U18129 (N_18129,N_17910,N_17930);
xor U18130 (N_18130,N_17872,N_17859);
nand U18131 (N_18131,N_17961,N_17970);
and U18132 (N_18132,N_17907,N_17864);
and U18133 (N_18133,N_17729,N_17851);
xnor U18134 (N_18134,N_17873,N_17891);
and U18135 (N_18135,N_17766,N_17885);
or U18136 (N_18136,N_17852,N_17818);
xnor U18137 (N_18137,N_17718,N_17752);
or U18138 (N_18138,N_17955,N_17841);
nand U18139 (N_18139,N_17973,N_17991);
nand U18140 (N_18140,N_17860,N_17758);
or U18141 (N_18141,N_17736,N_17989);
nor U18142 (N_18142,N_17786,N_17901);
xnor U18143 (N_18143,N_17771,N_17931);
nor U18144 (N_18144,N_17759,N_17808);
and U18145 (N_18145,N_17838,N_17727);
and U18146 (N_18146,N_17830,N_17858);
nand U18147 (N_18147,N_17824,N_17911);
xor U18148 (N_18148,N_17778,N_17976);
nand U18149 (N_18149,N_17982,N_17943);
and U18150 (N_18150,N_17987,N_17970);
or U18151 (N_18151,N_17810,N_17844);
xor U18152 (N_18152,N_17836,N_17812);
or U18153 (N_18153,N_17868,N_17914);
or U18154 (N_18154,N_17951,N_17734);
nor U18155 (N_18155,N_17725,N_17849);
and U18156 (N_18156,N_17929,N_17870);
nor U18157 (N_18157,N_17962,N_17717);
or U18158 (N_18158,N_17858,N_17915);
xor U18159 (N_18159,N_17830,N_17746);
nor U18160 (N_18160,N_17739,N_17942);
nor U18161 (N_18161,N_17819,N_17759);
and U18162 (N_18162,N_17733,N_17875);
nand U18163 (N_18163,N_17708,N_17858);
nand U18164 (N_18164,N_17749,N_17847);
nand U18165 (N_18165,N_17985,N_17736);
and U18166 (N_18166,N_17991,N_17789);
nor U18167 (N_18167,N_17874,N_17908);
and U18168 (N_18168,N_17753,N_17896);
xor U18169 (N_18169,N_17908,N_17898);
xnor U18170 (N_18170,N_17970,N_17849);
and U18171 (N_18171,N_17786,N_17843);
or U18172 (N_18172,N_17811,N_17894);
nand U18173 (N_18173,N_17994,N_17887);
or U18174 (N_18174,N_17711,N_17883);
and U18175 (N_18175,N_17972,N_17814);
nor U18176 (N_18176,N_17816,N_17881);
xor U18177 (N_18177,N_17987,N_17746);
and U18178 (N_18178,N_17945,N_17827);
nand U18179 (N_18179,N_17893,N_17904);
and U18180 (N_18180,N_17700,N_17887);
and U18181 (N_18181,N_17873,N_17718);
nand U18182 (N_18182,N_17801,N_17899);
and U18183 (N_18183,N_17700,N_17804);
xnor U18184 (N_18184,N_17912,N_17830);
xnor U18185 (N_18185,N_17786,N_17743);
nor U18186 (N_18186,N_17758,N_17741);
or U18187 (N_18187,N_17763,N_17962);
or U18188 (N_18188,N_17979,N_17842);
and U18189 (N_18189,N_17860,N_17903);
and U18190 (N_18190,N_17754,N_17737);
and U18191 (N_18191,N_17704,N_17952);
nor U18192 (N_18192,N_17855,N_17826);
xor U18193 (N_18193,N_17911,N_17833);
nor U18194 (N_18194,N_17920,N_17914);
nand U18195 (N_18195,N_17972,N_17900);
or U18196 (N_18196,N_17882,N_17780);
nand U18197 (N_18197,N_17956,N_17927);
nand U18198 (N_18198,N_17966,N_17793);
xnor U18199 (N_18199,N_17770,N_17810);
nor U18200 (N_18200,N_17805,N_17982);
and U18201 (N_18201,N_17973,N_17990);
nor U18202 (N_18202,N_17827,N_17770);
nor U18203 (N_18203,N_17839,N_17834);
and U18204 (N_18204,N_17964,N_17888);
nor U18205 (N_18205,N_17808,N_17953);
or U18206 (N_18206,N_17952,N_17917);
nand U18207 (N_18207,N_17897,N_17860);
and U18208 (N_18208,N_17801,N_17913);
and U18209 (N_18209,N_17922,N_17714);
and U18210 (N_18210,N_17895,N_17771);
nand U18211 (N_18211,N_17899,N_17706);
nand U18212 (N_18212,N_17784,N_17932);
nor U18213 (N_18213,N_17743,N_17710);
nor U18214 (N_18214,N_17762,N_17903);
and U18215 (N_18215,N_17733,N_17911);
nand U18216 (N_18216,N_17830,N_17937);
or U18217 (N_18217,N_17968,N_17938);
and U18218 (N_18218,N_17845,N_17769);
or U18219 (N_18219,N_17783,N_17808);
or U18220 (N_18220,N_17756,N_17833);
xor U18221 (N_18221,N_17840,N_17820);
or U18222 (N_18222,N_17893,N_17772);
and U18223 (N_18223,N_17765,N_17788);
or U18224 (N_18224,N_17791,N_17722);
xnor U18225 (N_18225,N_17887,N_17882);
or U18226 (N_18226,N_17808,N_17930);
nor U18227 (N_18227,N_17749,N_17828);
xnor U18228 (N_18228,N_17894,N_17968);
nor U18229 (N_18229,N_17917,N_17896);
xnor U18230 (N_18230,N_17934,N_17912);
nand U18231 (N_18231,N_17995,N_17771);
nor U18232 (N_18232,N_17954,N_17906);
and U18233 (N_18233,N_17758,N_17946);
xor U18234 (N_18234,N_17987,N_17921);
nand U18235 (N_18235,N_17939,N_17970);
and U18236 (N_18236,N_17793,N_17753);
nand U18237 (N_18237,N_17928,N_17884);
nand U18238 (N_18238,N_17968,N_17756);
nand U18239 (N_18239,N_17881,N_17821);
nand U18240 (N_18240,N_17703,N_17937);
xnor U18241 (N_18241,N_17853,N_17952);
xor U18242 (N_18242,N_17927,N_17731);
or U18243 (N_18243,N_17814,N_17714);
nor U18244 (N_18244,N_17893,N_17891);
or U18245 (N_18245,N_17988,N_17786);
xnor U18246 (N_18246,N_17986,N_17851);
and U18247 (N_18247,N_17874,N_17731);
or U18248 (N_18248,N_17780,N_17738);
nand U18249 (N_18249,N_17834,N_17976);
xor U18250 (N_18250,N_17923,N_17947);
and U18251 (N_18251,N_17821,N_17709);
xor U18252 (N_18252,N_17965,N_17726);
or U18253 (N_18253,N_17740,N_17995);
xor U18254 (N_18254,N_17710,N_17976);
nor U18255 (N_18255,N_17904,N_17918);
and U18256 (N_18256,N_17873,N_17797);
or U18257 (N_18257,N_17947,N_17985);
and U18258 (N_18258,N_17739,N_17737);
nor U18259 (N_18259,N_17854,N_17714);
or U18260 (N_18260,N_17826,N_17982);
xnor U18261 (N_18261,N_17871,N_17760);
or U18262 (N_18262,N_17757,N_17721);
or U18263 (N_18263,N_17812,N_17882);
xor U18264 (N_18264,N_17997,N_17815);
xnor U18265 (N_18265,N_17869,N_17998);
or U18266 (N_18266,N_17817,N_17993);
and U18267 (N_18267,N_17980,N_17750);
nand U18268 (N_18268,N_17814,N_17916);
or U18269 (N_18269,N_17739,N_17803);
or U18270 (N_18270,N_17702,N_17842);
nor U18271 (N_18271,N_17797,N_17915);
and U18272 (N_18272,N_17877,N_17858);
xnor U18273 (N_18273,N_17776,N_17822);
xnor U18274 (N_18274,N_17935,N_17905);
and U18275 (N_18275,N_17947,N_17735);
nand U18276 (N_18276,N_17846,N_17960);
xnor U18277 (N_18277,N_17881,N_17939);
and U18278 (N_18278,N_17742,N_17822);
xnor U18279 (N_18279,N_17929,N_17920);
nand U18280 (N_18280,N_17905,N_17747);
nand U18281 (N_18281,N_17893,N_17915);
xor U18282 (N_18282,N_17983,N_17921);
nor U18283 (N_18283,N_17722,N_17935);
or U18284 (N_18284,N_17783,N_17736);
or U18285 (N_18285,N_17936,N_17808);
and U18286 (N_18286,N_17875,N_17973);
or U18287 (N_18287,N_17816,N_17906);
xnor U18288 (N_18288,N_17766,N_17906);
xor U18289 (N_18289,N_17857,N_17997);
xnor U18290 (N_18290,N_17892,N_17937);
nand U18291 (N_18291,N_17994,N_17874);
nand U18292 (N_18292,N_17946,N_17788);
and U18293 (N_18293,N_17910,N_17847);
xor U18294 (N_18294,N_17964,N_17902);
nor U18295 (N_18295,N_17986,N_17701);
xor U18296 (N_18296,N_17780,N_17910);
or U18297 (N_18297,N_17970,N_17793);
and U18298 (N_18298,N_17827,N_17871);
and U18299 (N_18299,N_17870,N_17777);
nand U18300 (N_18300,N_18256,N_18112);
and U18301 (N_18301,N_18145,N_18187);
and U18302 (N_18302,N_18011,N_18063);
or U18303 (N_18303,N_18090,N_18023);
and U18304 (N_18304,N_18213,N_18097);
nand U18305 (N_18305,N_18053,N_18235);
nand U18306 (N_18306,N_18284,N_18052);
nor U18307 (N_18307,N_18272,N_18206);
xor U18308 (N_18308,N_18008,N_18222);
or U18309 (N_18309,N_18226,N_18022);
xnor U18310 (N_18310,N_18263,N_18133);
xnor U18311 (N_18311,N_18177,N_18050);
nor U18312 (N_18312,N_18179,N_18082);
nand U18313 (N_18313,N_18104,N_18246);
xor U18314 (N_18314,N_18231,N_18121);
nor U18315 (N_18315,N_18054,N_18149);
or U18316 (N_18316,N_18280,N_18016);
nor U18317 (N_18317,N_18026,N_18227);
xnor U18318 (N_18318,N_18183,N_18076);
nand U18319 (N_18319,N_18276,N_18119);
nand U18320 (N_18320,N_18293,N_18068);
nor U18321 (N_18321,N_18220,N_18135);
and U18322 (N_18322,N_18249,N_18048);
or U18323 (N_18323,N_18169,N_18283);
and U18324 (N_18324,N_18165,N_18018);
xor U18325 (N_18325,N_18230,N_18266);
nand U18326 (N_18326,N_18139,N_18003);
nor U18327 (N_18327,N_18225,N_18209);
or U18328 (N_18328,N_18241,N_18056);
xor U18329 (N_18329,N_18277,N_18282);
or U18330 (N_18330,N_18089,N_18116);
nand U18331 (N_18331,N_18221,N_18094);
and U18332 (N_18332,N_18142,N_18057);
or U18333 (N_18333,N_18204,N_18191);
nand U18334 (N_18334,N_18049,N_18025);
or U18335 (N_18335,N_18130,N_18137);
xnor U18336 (N_18336,N_18105,N_18152);
or U18337 (N_18337,N_18035,N_18158);
nand U18338 (N_18338,N_18066,N_18147);
xnor U18339 (N_18339,N_18136,N_18084);
nor U18340 (N_18340,N_18113,N_18170);
nand U18341 (N_18341,N_18101,N_18194);
nand U18342 (N_18342,N_18117,N_18155);
nand U18343 (N_18343,N_18217,N_18238);
xor U18344 (N_18344,N_18193,N_18037);
or U18345 (N_18345,N_18143,N_18093);
nor U18346 (N_18346,N_18019,N_18168);
or U18347 (N_18347,N_18207,N_18186);
and U18348 (N_18348,N_18058,N_18123);
and U18349 (N_18349,N_18297,N_18219);
and U18350 (N_18350,N_18013,N_18007);
and U18351 (N_18351,N_18218,N_18012);
xnor U18352 (N_18352,N_18108,N_18120);
nand U18353 (N_18353,N_18296,N_18188);
or U18354 (N_18354,N_18087,N_18279);
nor U18355 (N_18355,N_18131,N_18128);
xnor U18356 (N_18356,N_18159,N_18281);
and U18357 (N_18357,N_18138,N_18072);
or U18358 (N_18358,N_18181,N_18242);
xnor U18359 (N_18359,N_18212,N_18028);
nor U18360 (N_18360,N_18125,N_18247);
nand U18361 (N_18361,N_18260,N_18033);
or U18362 (N_18362,N_18189,N_18255);
nand U18363 (N_18363,N_18288,N_18254);
nor U18364 (N_18364,N_18092,N_18294);
nand U18365 (N_18365,N_18059,N_18267);
and U18366 (N_18366,N_18000,N_18109);
and U18367 (N_18367,N_18010,N_18286);
or U18368 (N_18368,N_18009,N_18151);
or U18369 (N_18369,N_18197,N_18110);
nor U18370 (N_18370,N_18083,N_18224);
nand U18371 (N_18371,N_18234,N_18073);
and U18372 (N_18372,N_18215,N_18268);
and U18373 (N_18373,N_18103,N_18040);
nand U18374 (N_18374,N_18166,N_18160);
and U18375 (N_18375,N_18292,N_18172);
nor U18376 (N_18376,N_18144,N_18192);
and U18377 (N_18377,N_18257,N_18253);
xor U18378 (N_18378,N_18069,N_18027);
nand U18379 (N_18379,N_18111,N_18100);
xnor U18380 (N_18380,N_18299,N_18259);
nor U18381 (N_18381,N_18102,N_18006);
nor U18382 (N_18382,N_18248,N_18150);
xor U18383 (N_18383,N_18201,N_18038);
nor U18384 (N_18384,N_18030,N_18132);
nor U18385 (N_18385,N_18034,N_18167);
xor U18386 (N_18386,N_18252,N_18001);
nand U18387 (N_18387,N_18126,N_18020);
or U18388 (N_18388,N_18262,N_18243);
nor U18389 (N_18389,N_18196,N_18229);
nand U18390 (N_18390,N_18062,N_18122);
nand U18391 (N_18391,N_18210,N_18129);
or U18392 (N_18392,N_18041,N_18127);
nor U18393 (N_18393,N_18140,N_18156);
nor U18394 (N_18394,N_18067,N_18232);
nand U18395 (N_18395,N_18075,N_18021);
or U18396 (N_18396,N_18216,N_18285);
or U18397 (N_18397,N_18065,N_18047);
and U18398 (N_18398,N_18261,N_18236);
nor U18399 (N_18399,N_18269,N_18039);
xor U18400 (N_18400,N_18161,N_18290);
nand U18401 (N_18401,N_18198,N_18184);
and U18402 (N_18402,N_18185,N_18244);
nand U18403 (N_18403,N_18265,N_18044);
xnor U18404 (N_18404,N_18061,N_18042);
and U18405 (N_18405,N_18163,N_18173);
and U18406 (N_18406,N_18287,N_18154);
nor U18407 (N_18407,N_18291,N_18202);
nor U18408 (N_18408,N_18153,N_18078);
xor U18409 (N_18409,N_18182,N_18014);
nor U18410 (N_18410,N_18180,N_18029);
and U18411 (N_18411,N_18245,N_18199);
nor U18412 (N_18412,N_18055,N_18045);
nand U18413 (N_18413,N_18205,N_18091);
nand U18414 (N_18414,N_18298,N_18174);
or U18415 (N_18415,N_18043,N_18031);
nor U18416 (N_18416,N_18079,N_18148);
or U18417 (N_18417,N_18118,N_18002);
nor U18418 (N_18418,N_18074,N_18141);
nor U18419 (N_18419,N_18278,N_18095);
nor U18420 (N_18420,N_18200,N_18250);
or U18421 (N_18421,N_18015,N_18264);
xor U18422 (N_18422,N_18070,N_18046);
xnor U18423 (N_18423,N_18178,N_18270);
nand U18424 (N_18424,N_18274,N_18157);
or U18425 (N_18425,N_18190,N_18115);
xor U18426 (N_18426,N_18295,N_18032);
and U18427 (N_18427,N_18195,N_18024);
or U18428 (N_18428,N_18077,N_18233);
xnor U18429 (N_18429,N_18146,N_18211);
or U18430 (N_18430,N_18134,N_18124);
xor U18431 (N_18431,N_18071,N_18258);
xor U18432 (N_18432,N_18088,N_18004);
xor U18433 (N_18433,N_18223,N_18208);
nand U18434 (N_18434,N_18251,N_18051);
nor U18435 (N_18435,N_18086,N_18017);
and U18436 (N_18436,N_18237,N_18080);
nor U18437 (N_18437,N_18228,N_18162);
or U18438 (N_18438,N_18098,N_18005);
nand U18439 (N_18439,N_18239,N_18289);
and U18440 (N_18440,N_18036,N_18275);
xor U18441 (N_18441,N_18106,N_18060);
nand U18442 (N_18442,N_18096,N_18164);
and U18443 (N_18443,N_18273,N_18064);
and U18444 (N_18444,N_18081,N_18085);
xnor U18445 (N_18445,N_18240,N_18107);
and U18446 (N_18446,N_18271,N_18203);
nor U18447 (N_18447,N_18171,N_18214);
and U18448 (N_18448,N_18176,N_18099);
or U18449 (N_18449,N_18175,N_18114);
nor U18450 (N_18450,N_18013,N_18125);
nor U18451 (N_18451,N_18105,N_18265);
or U18452 (N_18452,N_18201,N_18237);
nand U18453 (N_18453,N_18210,N_18153);
nand U18454 (N_18454,N_18027,N_18287);
and U18455 (N_18455,N_18042,N_18122);
nand U18456 (N_18456,N_18003,N_18253);
xor U18457 (N_18457,N_18120,N_18123);
nand U18458 (N_18458,N_18166,N_18042);
xnor U18459 (N_18459,N_18210,N_18110);
nor U18460 (N_18460,N_18227,N_18047);
xor U18461 (N_18461,N_18177,N_18162);
nand U18462 (N_18462,N_18253,N_18234);
xor U18463 (N_18463,N_18028,N_18007);
nor U18464 (N_18464,N_18065,N_18077);
nand U18465 (N_18465,N_18256,N_18156);
xor U18466 (N_18466,N_18245,N_18109);
nand U18467 (N_18467,N_18178,N_18077);
and U18468 (N_18468,N_18139,N_18054);
nor U18469 (N_18469,N_18020,N_18062);
nand U18470 (N_18470,N_18258,N_18276);
nor U18471 (N_18471,N_18104,N_18299);
and U18472 (N_18472,N_18111,N_18224);
and U18473 (N_18473,N_18190,N_18107);
nor U18474 (N_18474,N_18163,N_18045);
nand U18475 (N_18475,N_18072,N_18199);
nand U18476 (N_18476,N_18115,N_18111);
xor U18477 (N_18477,N_18093,N_18076);
xnor U18478 (N_18478,N_18165,N_18199);
xor U18479 (N_18479,N_18137,N_18187);
nand U18480 (N_18480,N_18075,N_18071);
xor U18481 (N_18481,N_18251,N_18140);
nand U18482 (N_18482,N_18050,N_18092);
or U18483 (N_18483,N_18175,N_18219);
nand U18484 (N_18484,N_18140,N_18085);
and U18485 (N_18485,N_18247,N_18040);
or U18486 (N_18486,N_18265,N_18056);
or U18487 (N_18487,N_18127,N_18266);
xnor U18488 (N_18488,N_18014,N_18292);
or U18489 (N_18489,N_18177,N_18200);
xnor U18490 (N_18490,N_18108,N_18289);
xnor U18491 (N_18491,N_18130,N_18243);
or U18492 (N_18492,N_18063,N_18248);
and U18493 (N_18493,N_18277,N_18133);
xnor U18494 (N_18494,N_18012,N_18150);
or U18495 (N_18495,N_18067,N_18114);
or U18496 (N_18496,N_18118,N_18225);
nand U18497 (N_18497,N_18290,N_18233);
nand U18498 (N_18498,N_18141,N_18037);
and U18499 (N_18499,N_18279,N_18206);
or U18500 (N_18500,N_18064,N_18009);
nor U18501 (N_18501,N_18126,N_18047);
or U18502 (N_18502,N_18128,N_18134);
or U18503 (N_18503,N_18003,N_18275);
and U18504 (N_18504,N_18036,N_18154);
and U18505 (N_18505,N_18181,N_18073);
xnor U18506 (N_18506,N_18097,N_18055);
and U18507 (N_18507,N_18015,N_18194);
or U18508 (N_18508,N_18272,N_18202);
nor U18509 (N_18509,N_18007,N_18030);
or U18510 (N_18510,N_18259,N_18180);
xnor U18511 (N_18511,N_18026,N_18145);
and U18512 (N_18512,N_18016,N_18023);
xnor U18513 (N_18513,N_18145,N_18097);
nand U18514 (N_18514,N_18284,N_18217);
nand U18515 (N_18515,N_18093,N_18201);
xnor U18516 (N_18516,N_18005,N_18029);
nand U18517 (N_18517,N_18183,N_18262);
xnor U18518 (N_18518,N_18179,N_18217);
and U18519 (N_18519,N_18161,N_18063);
or U18520 (N_18520,N_18101,N_18144);
or U18521 (N_18521,N_18210,N_18294);
xor U18522 (N_18522,N_18137,N_18085);
nand U18523 (N_18523,N_18024,N_18263);
xnor U18524 (N_18524,N_18126,N_18247);
xnor U18525 (N_18525,N_18211,N_18064);
nand U18526 (N_18526,N_18173,N_18133);
or U18527 (N_18527,N_18060,N_18030);
or U18528 (N_18528,N_18082,N_18225);
nor U18529 (N_18529,N_18261,N_18149);
or U18530 (N_18530,N_18152,N_18268);
nand U18531 (N_18531,N_18138,N_18204);
xnor U18532 (N_18532,N_18026,N_18162);
nor U18533 (N_18533,N_18284,N_18114);
and U18534 (N_18534,N_18155,N_18209);
and U18535 (N_18535,N_18112,N_18139);
nand U18536 (N_18536,N_18293,N_18087);
xor U18537 (N_18537,N_18197,N_18120);
or U18538 (N_18538,N_18143,N_18028);
xor U18539 (N_18539,N_18287,N_18037);
and U18540 (N_18540,N_18295,N_18185);
or U18541 (N_18541,N_18269,N_18278);
and U18542 (N_18542,N_18081,N_18062);
nand U18543 (N_18543,N_18047,N_18235);
nor U18544 (N_18544,N_18000,N_18192);
and U18545 (N_18545,N_18135,N_18095);
nor U18546 (N_18546,N_18116,N_18144);
nor U18547 (N_18547,N_18073,N_18256);
nor U18548 (N_18548,N_18137,N_18177);
xnor U18549 (N_18549,N_18057,N_18152);
xor U18550 (N_18550,N_18169,N_18136);
xor U18551 (N_18551,N_18137,N_18102);
or U18552 (N_18552,N_18002,N_18290);
xnor U18553 (N_18553,N_18252,N_18250);
xor U18554 (N_18554,N_18203,N_18016);
or U18555 (N_18555,N_18281,N_18270);
xnor U18556 (N_18556,N_18142,N_18033);
or U18557 (N_18557,N_18221,N_18009);
and U18558 (N_18558,N_18040,N_18173);
nor U18559 (N_18559,N_18281,N_18273);
and U18560 (N_18560,N_18158,N_18188);
and U18561 (N_18561,N_18164,N_18141);
or U18562 (N_18562,N_18283,N_18268);
nand U18563 (N_18563,N_18045,N_18248);
or U18564 (N_18564,N_18289,N_18199);
nand U18565 (N_18565,N_18168,N_18189);
and U18566 (N_18566,N_18156,N_18131);
and U18567 (N_18567,N_18018,N_18065);
nand U18568 (N_18568,N_18237,N_18169);
or U18569 (N_18569,N_18006,N_18118);
and U18570 (N_18570,N_18134,N_18225);
and U18571 (N_18571,N_18130,N_18200);
nor U18572 (N_18572,N_18288,N_18157);
nand U18573 (N_18573,N_18205,N_18251);
or U18574 (N_18574,N_18084,N_18083);
nand U18575 (N_18575,N_18249,N_18010);
or U18576 (N_18576,N_18200,N_18270);
and U18577 (N_18577,N_18192,N_18060);
or U18578 (N_18578,N_18298,N_18226);
xor U18579 (N_18579,N_18020,N_18246);
nand U18580 (N_18580,N_18202,N_18022);
and U18581 (N_18581,N_18116,N_18293);
nor U18582 (N_18582,N_18089,N_18220);
nor U18583 (N_18583,N_18109,N_18077);
xor U18584 (N_18584,N_18261,N_18126);
nor U18585 (N_18585,N_18279,N_18112);
or U18586 (N_18586,N_18020,N_18096);
or U18587 (N_18587,N_18083,N_18111);
xor U18588 (N_18588,N_18272,N_18140);
or U18589 (N_18589,N_18282,N_18160);
xor U18590 (N_18590,N_18281,N_18197);
nand U18591 (N_18591,N_18177,N_18060);
or U18592 (N_18592,N_18016,N_18057);
and U18593 (N_18593,N_18231,N_18116);
and U18594 (N_18594,N_18169,N_18140);
nand U18595 (N_18595,N_18002,N_18052);
nor U18596 (N_18596,N_18122,N_18275);
and U18597 (N_18597,N_18084,N_18013);
xor U18598 (N_18598,N_18122,N_18077);
nand U18599 (N_18599,N_18297,N_18217);
nor U18600 (N_18600,N_18378,N_18308);
or U18601 (N_18601,N_18563,N_18537);
nor U18602 (N_18602,N_18581,N_18521);
or U18603 (N_18603,N_18444,N_18586);
and U18604 (N_18604,N_18369,N_18435);
and U18605 (N_18605,N_18570,N_18590);
nor U18606 (N_18606,N_18312,N_18506);
nor U18607 (N_18607,N_18485,N_18463);
xor U18608 (N_18608,N_18496,N_18382);
nor U18609 (N_18609,N_18399,N_18480);
nand U18610 (N_18610,N_18531,N_18339);
nand U18611 (N_18611,N_18388,N_18593);
nor U18612 (N_18612,N_18420,N_18386);
xnor U18613 (N_18613,N_18477,N_18458);
or U18614 (N_18614,N_18445,N_18501);
nand U18615 (N_18615,N_18589,N_18333);
xnor U18616 (N_18616,N_18542,N_18544);
nor U18617 (N_18617,N_18343,N_18498);
or U18618 (N_18618,N_18499,N_18509);
nor U18619 (N_18619,N_18440,N_18599);
xor U18620 (N_18620,N_18391,N_18331);
nand U18621 (N_18621,N_18528,N_18529);
nor U18622 (N_18622,N_18304,N_18443);
xor U18623 (N_18623,N_18527,N_18497);
nand U18624 (N_18624,N_18511,N_18494);
and U18625 (N_18625,N_18492,N_18552);
or U18626 (N_18626,N_18351,N_18533);
nor U18627 (N_18627,N_18575,N_18321);
nand U18628 (N_18628,N_18592,N_18406);
nand U18629 (N_18629,N_18488,N_18547);
xnor U18630 (N_18630,N_18394,N_18344);
xor U18631 (N_18631,N_18483,N_18522);
or U18632 (N_18632,N_18454,N_18309);
nand U18633 (N_18633,N_18517,N_18327);
or U18634 (N_18634,N_18441,N_18409);
nor U18635 (N_18635,N_18553,N_18535);
xor U18636 (N_18636,N_18461,N_18595);
xnor U18637 (N_18637,N_18433,N_18524);
nand U18638 (N_18638,N_18315,N_18389);
nor U18639 (N_18639,N_18414,N_18370);
and U18640 (N_18640,N_18324,N_18402);
nand U18641 (N_18641,N_18360,N_18512);
or U18642 (N_18642,N_18404,N_18486);
nand U18643 (N_18643,N_18548,N_18325);
nand U18644 (N_18644,N_18313,N_18419);
nand U18645 (N_18645,N_18451,N_18476);
and U18646 (N_18646,N_18436,N_18597);
or U18647 (N_18647,N_18437,N_18412);
nor U18648 (N_18648,N_18460,N_18314);
or U18649 (N_18649,N_18352,N_18596);
and U18650 (N_18650,N_18478,N_18427);
xor U18651 (N_18651,N_18532,N_18474);
nand U18652 (N_18652,N_18543,N_18561);
and U18653 (N_18653,N_18449,N_18525);
or U18654 (N_18654,N_18493,N_18362);
nor U18655 (N_18655,N_18503,N_18549);
xor U18656 (N_18656,N_18470,N_18305);
xnor U18657 (N_18657,N_18357,N_18417);
xor U18658 (N_18658,N_18408,N_18457);
or U18659 (N_18659,N_18588,N_18459);
xnor U18660 (N_18660,N_18515,N_18426);
and U18661 (N_18661,N_18585,N_18448);
nor U18662 (N_18662,N_18566,N_18395);
or U18663 (N_18663,N_18405,N_18425);
nor U18664 (N_18664,N_18371,N_18345);
nand U18665 (N_18665,N_18418,N_18484);
and U18666 (N_18666,N_18300,N_18536);
and U18667 (N_18667,N_18337,N_18573);
and U18668 (N_18668,N_18479,N_18487);
nor U18669 (N_18669,N_18349,N_18340);
nand U18670 (N_18670,N_18372,N_18567);
xnor U18671 (N_18671,N_18383,N_18350);
and U18672 (N_18672,N_18375,N_18356);
and U18673 (N_18673,N_18452,N_18385);
nor U18674 (N_18674,N_18578,N_18353);
or U18675 (N_18675,N_18554,N_18518);
nor U18676 (N_18676,N_18472,N_18541);
or U18677 (N_18677,N_18368,N_18323);
nand U18678 (N_18678,N_18450,N_18363);
nand U18679 (N_18679,N_18550,N_18513);
nand U18680 (N_18680,N_18311,N_18447);
nand U18681 (N_18681,N_18374,N_18322);
xor U18682 (N_18682,N_18576,N_18332);
and U18683 (N_18683,N_18560,N_18359);
or U18684 (N_18684,N_18401,N_18551);
and U18685 (N_18685,N_18464,N_18577);
xnor U18686 (N_18686,N_18367,N_18358);
or U18687 (N_18687,N_18455,N_18526);
xor U18688 (N_18688,N_18317,N_18456);
and U18689 (N_18689,N_18462,N_18580);
nand U18690 (N_18690,N_18502,N_18355);
and U18691 (N_18691,N_18545,N_18407);
or U18692 (N_18692,N_18316,N_18336);
xor U18693 (N_18693,N_18466,N_18428);
xnor U18694 (N_18694,N_18438,N_18432);
nor U18695 (N_18695,N_18342,N_18390);
xnor U18696 (N_18696,N_18530,N_18468);
nand U18697 (N_18697,N_18400,N_18523);
nor U18698 (N_18698,N_18446,N_18574);
and U18699 (N_18699,N_18354,N_18301);
and U18700 (N_18700,N_18565,N_18377);
nand U18701 (N_18701,N_18546,N_18397);
xnor U18702 (N_18702,N_18539,N_18594);
and U18703 (N_18703,N_18306,N_18519);
xor U18704 (N_18704,N_18334,N_18429);
and U18705 (N_18705,N_18380,N_18341);
and U18706 (N_18706,N_18411,N_18398);
xor U18707 (N_18707,N_18422,N_18557);
nor U18708 (N_18708,N_18471,N_18421);
or U18709 (N_18709,N_18500,N_18538);
and U18710 (N_18710,N_18307,N_18413);
nand U18711 (N_18711,N_18482,N_18392);
nand U18712 (N_18712,N_18582,N_18489);
nor U18713 (N_18713,N_18347,N_18366);
nor U18714 (N_18714,N_18364,N_18453);
or U18715 (N_18715,N_18584,N_18504);
nand U18716 (N_18716,N_18556,N_18328);
or U18717 (N_18717,N_18510,N_18571);
nand U18718 (N_18718,N_18520,N_18348);
and U18719 (N_18719,N_18572,N_18361);
nand U18720 (N_18720,N_18579,N_18481);
nand U18721 (N_18721,N_18583,N_18423);
xor U18722 (N_18722,N_18326,N_18424);
nand U18723 (N_18723,N_18491,N_18507);
or U18724 (N_18724,N_18318,N_18384);
or U18725 (N_18725,N_18338,N_18564);
and U18726 (N_18726,N_18376,N_18516);
nor U18727 (N_18727,N_18431,N_18562);
and U18728 (N_18728,N_18559,N_18505);
nor U18729 (N_18729,N_18469,N_18490);
xnor U18730 (N_18730,N_18346,N_18569);
and U18731 (N_18731,N_18310,N_18514);
or U18732 (N_18732,N_18534,N_18381);
nand U18733 (N_18733,N_18555,N_18598);
or U18734 (N_18734,N_18473,N_18373);
and U18735 (N_18735,N_18475,N_18320);
nor U18736 (N_18736,N_18587,N_18379);
and U18737 (N_18737,N_18302,N_18430);
nor U18738 (N_18738,N_18303,N_18442);
xnor U18739 (N_18739,N_18568,N_18465);
nor U18740 (N_18740,N_18434,N_18467);
xor U18741 (N_18741,N_18393,N_18330);
and U18742 (N_18742,N_18439,N_18415);
or U18743 (N_18743,N_18403,N_18329);
nor U18744 (N_18744,N_18508,N_18387);
xor U18745 (N_18745,N_18558,N_18540);
or U18746 (N_18746,N_18410,N_18396);
nor U18747 (N_18747,N_18591,N_18365);
xnor U18748 (N_18748,N_18319,N_18416);
or U18749 (N_18749,N_18335,N_18495);
nor U18750 (N_18750,N_18315,N_18445);
nand U18751 (N_18751,N_18323,N_18387);
nor U18752 (N_18752,N_18324,N_18326);
nor U18753 (N_18753,N_18594,N_18312);
xnor U18754 (N_18754,N_18496,N_18378);
xnor U18755 (N_18755,N_18515,N_18516);
and U18756 (N_18756,N_18441,N_18477);
nand U18757 (N_18757,N_18589,N_18339);
nand U18758 (N_18758,N_18582,N_18331);
nand U18759 (N_18759,N_18515,N_18434);
nor U18760 (N_18760,N_18523,N_18599);
or U18761 (N_18761,N_18306,N_18503);
nand U18762 (N_18762,N_18365,N_18301);
and U18763 (N_18763,N_18521,N_18381);
nand U18764 (N_18764,N_18390,N_18344);
xnor U18765 (N_18765,N_18301,N_18350);
and U18766 (N_18766,N_18544,N_18566);
or U18767 (N_18767,N_18586,N_18322);
and U18768 (N_18768,N_18533,N_18535);
or U18769 (N_18769,N_18523,N_18479);
xnor U18770 (N_18770,N_18419,N_18552);
and U18771 (N_18771,N_18304,N_18416);
nor U18772 (N_18772,N_18484,N_18526);
nor U18773 (N_18773,N_18335,N_18492);
nand U18774 (N_18774,N_18531,N_18381);
xnor U18775 (N_18775,N_18450,N_18320);
and U18776 (N_18776,N_18558,N_18317);
and U18777 (N_18777,N_18473,N_18476);
nor U18778 (N_18778,N_18438,N_18412);
and U18779 (N_18779,N_18574,N_18577);
nor U18780 (N_18780,N_18482,N_18393);
and U18781 (N_18781,N_18429,N_18475);
xnor U18782 (N_18782,N_18494,N_18586);
nand U18783 (N_18783,N_18327,N_18364);
nand U18784 (N_18784,N_18399,N_18304);
nor U18785 (N_18785,N_18347,N_18541);
or U18786 (N_18786,N_18331,N_18499);
nor U18787 (N_18787,N_18599,N_18419);
nor U18788 (N_18788,N_18304,N_18500);
nor U18789 (N_18789,N_18472,N_18549);
or U18790 (N_18790,N_18427,N_18505);
or U18791 (N_18791,N_18301,N_18386);
nand U18792 (N_18792,N_18459,N_18403);
xor U18793 (N_18793,N_18312,N_18585);
nor U18794 (N_18794,N_18561,N_18571);
or U18795 (N_18795,N_18505,N_18496);
and U18796 (N_18796,N_18357,N_18400);
or U18797 (N_18797,N_18499,N_18373);
and U18798 (N_18798,N_18527,N_18522);
xnor U18799 (N_18799,N_18366,N_18308);
and U18800 (N_18800,N_18452,N_18315);
nand U18801 (N_18801,N_18358,N_18425);
nor U18802 (N_18802,N_18568,N_18360);
xnor U18803 (N_18803,N_18418,N_18376);
or U18804 (N_18804,N_18533,N_18507);
xor U18805 (N_18805,N_18449,N_18521);
nor U18806 (N_18806,N_18411,N_18316);
nor U18807 (N_18807,N_18309,N_18305);
nand U18808 (N_18808,N_18493,N_18391);
and U18809 (N_18809,N_18461,N_18347);
nand U18810 (N_18810,N_18313,N_18504);
or U18811 (N_18811,N_18382,N_18375);
xor U18812 (N_18812,N_18560,N_18483);
or U18813 (N_18813,N_18387,N_18341);
nor U18814 (N_18814,N_18489,N_18457);
nor U18815 (N_18815,N_18336,N_18395);
nand U18816 (N_18816,N_18511,N_18401);
nand U18817 (N_18817,N_18412,N_18362);
xnor U18818 (N_18818,N_18564,N_18467);
xnor U18819 (N_18819,N_18302,N_18520);
nand U18820 (N_18820,N_18330,N_18375);
nand U18821 (N_18821,N_18365,N_18488);
and U18822 (N_18822,N_18511,N_18328);
xnor U18823 (N_18823,N_18457,N_18394);
nor U18824 (N_18824,N_18488,N_18490);
xnor U18825 (N_18825,N_18549,N_18317);
and U18826 (N_18826,N_18306,N_18449);
and U18827 (N_18827,N_18538,N_18409);
and U18828 (N_18828,N_18336,N_18559);
nor U18829 (N_18829,N_18532,N_18588);
or U18830 (N_18830,N_18435,N_18538);
nand U18831 (N_18831,N_18533,N_18357);
nor U18832 (N_18832,N_18364,N_18351);
or U18833 (N_18833,N_18542,N_18583);
xor U18834 (N_18834,N_18539,N_18496);
or U18835 (N_18835,N_18315,N_18517);
xor U18836 (N_18836,N_18590,N_18397);
or U18837 (N_18837,N_18327,N_18335);
nor U18838 (N_18838,N_18486,N_18366);
nor U18839 (N_18839,N_18343,N_18425);
nand U18840 (N_18840,N_18413,N_18559);
xor U18841 (N_18841,N_18593,N_18596);
nand U18842 (N_18842,N_18301,N_18309);
xor U18843 (N_18843,N_18314,N_18473);
nand U18844 (N_18844,N_18326,N_18579);
and U18845 (N_18845,N_18300,N_18586);
and U18846 (N_18846,N_18444,N_18568);
and U18847 (N_18847,N_18433,N_18570);
or U18848 (N_18848,N_18520,N_18501);
nor U18849 (N_18849,N_18514,N_18347);
nand U18850 (N_18850,N_18562,N_18476);
xor U18851 (N_18851,N_18303,N_18309);
and U18852 (N_18852,N_18379,N_18368);
and U18853 (N_18853,N_18388,N_18582);
and U18854 (N_18854,N_18545,N_18490);
and U18855 (N_18855,N_18317,N_18393);
and U18856 (N_18856,N_18510,N_18330);
nand U18857 (N_18857,N_18374,N_18584);
nor U18858 (N_18858,N_18302,N_18351);
nand U18859 (N_18859,N_18543,N_18567);
nand U18860 (N_18860,N_18303,N_18511);
xor U18861 (N_18861,N_18564,N_18592);
nor U18862 (N_18862,N_18391,N_18367);
or U18863 (N_18863,N_18513,N_18591);
and U18864 (N_18864,N_18458,N_18459);
nor U18865 (N_18865,N_18408,N_18508);
nor U18866 (N_18866,N_18376,N_18396);
nand U18867 (N_18867,N_18564,N_18335);
and U18868 (N_18868,N_18486,N_18479);
or U18869 (N_18869,N_18356,N_18474);
nor U18870 (N_18870,N_18530,N_18451);
xor U18871 (N_18871,N_18378,N_18559);
and U18872 (N_18872,N_18424,N_18509);
or U18873 (N_18873,N_18308,N_18304);
nand U18874 (N_18874,N_18504,N_18365);
nand U18875 (N_18875,N_18452,N_18316);
or U18876 (N_18876,N_18470,N_18457);
xor U18877 (N_18877,N_18393,N_18389);
xor U18878 (N_18878,N_18342,N_18457);
or U18879 (N_18879,N_18403,N_18560);
or U18880 (N_18880,N_18352,N_18553);
and U18881 (N_18881,N_18392,N_18395);
or U18882 (N_18882,N_18580,N_18559);
nand U18883 (N_18883,N_18509,N_18518);
and U18884 (N_18884,N_18568,N_18463);
xor U18885 (N_18885,N_18366,N_18564);
and U18886 (N_18886,N_18313,N_18408);
or U18887 (N_18887,N_18581,N_18487);
nor U18888 (N_18888,N_18338,N_18570);
nand U18889 (N_18889,N_18311,N_18440);
xor U18890 (N_18890,N_18544,N_18355);
nor U18891 (N_18891,N_18403,N_18512);
and U18892 (N_18892,N_18505,N_18404);
xnor U18893 (N_18893,N_18586,N_18489);
nor U18894 (N_18894,N_18408,N_18331);
and U18895 (N_18895,N_18326,N_18379);
nor U18896 (N_18896,N_18381,N_18410);
nand U18897 (N_18897,N_18507,N_18511);
or U18898 (N_18898,N_18503,N_18325);
and U18899 (N_18899,N_18500,N_18407);
nand U18900 (N_18900,N_18755,N_18698);
nor U18901 (N_18901,N_18677,N_18896);
xnor U18902 (N_18902,N_18888,N_18804);
and U18903 (N_18903,N_18817,N_18620);
nand U18904 (N_18904,N_18822,N_18783);
nor U18905 (N_18905,N_18812,N_18625);
nor U18906 (N_18906,N_18768,N_18671);
or U18907 (N_18907,N_18895,N_18857);
and U18908 (N_18908,N_18887,N_18645);
or U18909 (N_18909,N_18830,N_18823);
or U18910 (N_18910,N_18735,N_18655);
or U18911 (N_18911,N_18886,N_18672);
or U18912 (N_18912,N_18686,N_18719);
nor U18913 (N_18913,N_18639,N_18876);
and U18914 (N_18914,N_18856,N_18759);
nand U18915 (N_18915,N_18780,N_18687);
xor U18916 (N_18916,N_18694,N_18846);
xor U18917 (N_18917,N_18806,N_18824);
xor U18918 (N_18918,N_18853,N_18800);
nor U18919 (N_18919,N_18743,N_18633);
nand U18920 (N_18920,N_18665,N_18637);
and U18921 (N_18921,N_18730,N_18872);
nand U18922 (N_18922,N_18814,N_18722);
nor U18923 (N_18923,N_18842,N_18855);
xor U18924 (N_18924,N_18868,N_18899);
nand U18925 (N_18925,N_18852,N_18667);
or U18926 (N_18926,N_18798,N_18858);
or U18927 (N_18927,N_18769,N_18882);
or U18928 (N_18928,N_18619,N_18721);
xor U18929 (N_18929,N_18656,N_18816);
nand U18930 (N_18930,N_18675,N_18737);
xor U18931 (N_18931,N_18771,N_18713);
and U18932 (N_18932,N_18650,N_18701);
or U18933 (N_18933,N_18635,N_18708);
and U18934 (N_18934,N_18603,N_18731);
and U18935 (N_18935,N_18761,N_18794);
xnor U18936 (N_18936,N_18614,N_18851);
or U18937 (N_18937,N_18616,N_18615);
and U18938 (N_18938,N_18795,N_18765);
nand U18939 (N_18939,N_18757,N_18610);
nor U18940 (N_18940,N_18696,N_18744);
nand U18941 (N_18941,N_18600,N_18704);
or U18942 (N_18942,N_18889,N_18779);
nand U18943 (N_18943,N_18837,N_18753);
nor U18944 (N_18944,N_18683,N_18717);
and U18945 (N_18945,N_18624,N_18809);
xor U18946 (N_18946,N_18703,N_18792);
and U18947 (N_18947,N_18649,N_18734);
nand U18948 (N_18948,N_18728,N_18727);
xnor U18949 (N_18949,N_18623,N_18848);
nor U18950 (N_18950,N_18849,N_18748);
xor U18951 (N_18951,N_18775,N_18751);
and U18952 (N_18952,N_18670,N_18894);
nor U18953 (N_18953,N_18602,N_18709);
and U18954 (N_18954,N_18631,N_18838);
or U18955 (N_18955,N_18821,N_18773);
and U18956 (N_18956,N_18658,N_18636);
or U18957 (N_18957,N_18850,N_18724);
nand U18958 (N_18958,N_18705,N_18678);
nand U18959 (N_18959,N_18700,N_18844);
nand U18960 (N_18960,N_18776,N_18668);
nor U18961 (N_18961,N_18819,N_18706);
nand U18962 (N_18962,N_18787,N_18745);
xnor U18963 (N_18963,N_18766,N_18691);
and U18964 (N_18964,N_18892,N_18747);
or U18965 (N_18965,N_18750,N_18866);
or U18966 (N_18966,N_18752,N_18647);
xnor U18967 (N_18967,N_18797,N_18622);
nor U18968 (N_18968,N_18867,N_18841);
xor U18969 (N_18969,N_18786,N_18788);
nor U18970 (N_18970,N_18644,N_18738);
nor U18971 (N_18971,N_18833,N_18692);
and U18972 (N_18972,N_18638,N_18825);
and U18973 (N_18973,N_18746,N_18652);
and U18974 (N_18974,N_18865,N_18732);
nand U18975 (N_18975,N_18859,N_18653);
and U18976 (N_18976,N_18808,N_18684);
nand U18977 (N_18977,N_18789,N_18718);
nor U18978 (N_18978,N_18862,N_18818);
nand U18979 (N_18979,N_18871,N_18885);
nor U18980 (N_18980,N_18762,N_18664);
xnor U18981 (N_18981,N_18811,N_18661);
xor U18982 (N_18982,N_18836,N_18605);
nand U18983 (N_18983,N_18688,N_18720);
nor U18984 (N_18984,N_18883,N_18660);
nor U18985 (N_18985,N_18803,N_18760);
and U18986 (N_18986,N_18863,N_18891);
or U18987 (N_18987,N_18861,N_18749);
xnor U18988 (N_18988,N_18770,N_18711);
or U18989 (N_18989,N_18604,N_18831);
nand U18990 (N_18990,N_18877,N_18659);
or U18991 (N_18991,N_18707,N_18782);
and U18992 (N_18992,N_18716,N_18632);
and U18993 (N_18993,N_18695,N_18646);
xor U18994 (N_18994,N_18870,N_18893);
nand U18995 (N_18995,N_18826,N_18875);
nand U18996 (N_18996,N_18714,N_18608);
xnor U18997 (N_18997,N_18666,N_18679);
xor U18998 (N_18998,N_18642,N_18740);
or U18999 (N_18999,N_18810,N_18643);
or U19000 (N_19000,N_18606,N_18878);
nand U19001 (N_19001,N_18767,N_18777);
or U19002 (N_19002,N_18802,N_18881);
nand U19003 (N_19003,N_18725,N_18621);
nand U19004 (N_19004,N_18754,N_18827);
and U19005 (N_19005,N_18676,N_18805);
nor U19006 (N_19006,N_18880,N_18860);
or U19007 (N_19007,N_18854,N_18820);
or U19008 (N_19008,N_18685,N_18791);
or U19009 (N_19009,N_18634,N_18607);
and U19010 (N_19010,N_18726,N_18710);
nand U19011 (N_19011,N_18763,N_18807);
nor U19012 (N_19012,N_18657,N_18648);
and U19013 (N_19013,N_18674,N_18715);
and U19014 (N_19014,N_18813,N_18793);
and U19015 (N_19015,N_18879,N_18873);
xor U19016 (N_19016,N_18693,N_18617);
nor U19017 (N_19017,N_18781,N_18663);
or U19018 (N_19018,N_18640,N_18772);
xor U19019 (N_19019,N_18864,N_18758);
xor U19020 (N_19020,N_18690,N_18815);
or U19021 (N_19021,N_18682,N_18733);
nand U19022 (N_19022,N_18790,N_18785);
xor U19023 (N_19023,N_18702,N_18613);
or U19024 (N_19024,N_18778,N_18839);
nand U19025 (N_19025,N_18689,N_18840);
nor U19026 (N_19026,N_18832,N_18874);
nand U19027 (N_19027,N_18801,N_18756);
or U19028 (N_19028,N_18618,N_18669);
xor U19029 (N_19029,N_18680,N_18799);
or U19030 (N_19030,N_18662,N_18739);
nor U19031 (N_19031,N_18699,N_18884);
xor U19032 (N_19032,N_18784,N_18835);
nor U19033 (N_19033,N_18796,N_18898);
and U19034 (N_19034,N_18629,N_18626);
and U19035 (N_19035,N_18628,N_18834);
and U19036 (N_19036,N_18774,N_18729);
nor U19037 (N_19037,N_18736,N_18723);
nand U19038 (N_19038,N_18712,N_18869);
xor U19039 (N_19039,N_18845,N_18673);
nand U19040 (N_19040,N_18843,N_18697);
or U19041 (N_19041,N_18609,N_18764);
nor U19042 (N_19042,N_18654,N_18651);
and U19043 (N_19043,N_18829,N_18847);
and U19044 (N_19044,N_18742,N_18630);
xor U19045 (N_19045,N_18890,N_18627);
nand U19046 (N_19046,N_18641,N_18828);
nand U19047 (N_19047,N_18611,N_18612);
nor U19048 (N_19048,N_18741,N_18681);
nor U19049 (N_19049,N_18897,N_18601);
xnor U19050 (N_19050,N_18880,N_18818);
and U19051 (N_19051,N_18806,N_18851);
and U19052 (N_19052,N_18626,N_18745);
nand U19053 (N_19053,N_18611,N_18681);
nand U19054 (N_19054,N_18747,N_18682);
or U19055 (N_19055,N_18705,N_18730);
or U19056 (N_19056,N_18894,N_18707);
xnor U19057 (N_19057,N_18628,N_18783);
or U19058 (N_19058,N_18616,N_18895);
xnor U19059 (N_19059,N_18700,N_18875);
nand U19060 (N_19060,N_18852,N_18757);
or U19061 (N_19061,N_18656,N_18790);
nor U19062 (N_19062,N_18754,N_18739);
nand U19063 (N_19063,N_18748,N_18798);
nand U19064 (N_19064,N_18745,N_18845);
xnor U19065 (N_19065,N_18718,N_18855);
xor U19066 (N_19066,N_18611,N_18851);
nand U19067 (N_19067,N_18875,N_18726);
xor U19068 (N_19068,N_18775,N_18841);
xor U19069 (N_19069,N_18758,N_18745);
nand U19070 (N_19070,N_18817,N_18651);
and U19071 (N_19071,N_18852,N_18604);
nand U19072 (N_19072,N_18700,N_18881);
nor U19073 (N_19073,N_18716,N_18774);
nand U19074 (N_19074,N_18738,N_18836);
xor U19075 (N_19075,N_18779,N_18865);
and U19076 (N_19076,N_18776,N_18742);
or U19077 (N_19077,N_18730,N_18711);
and U19078 (N_19078,N_18757,N_18815);
nand U19079 (N_19079,N_18859,N_18693);
or U19080 (N_19080,N_18742,N_18809);
nor U19081 (N_19081,N_18665,N_18795);
nor U19082 (N_19082,N_18810,N_18695);
and U19083 (N_19083,N_18723,N_18692);
or U19084 (N_19084,N_18843,N_18871);
nor U19085 (N_19085,N_18794,N_18871);
xnor U19086 (N_19086,N_18725,N_18623);
xnor U19087 (N_19087,N_18897,N_18682);
nand U19088 (N_19088,N_18686,N_18818);
and U19089 (N_19089,N_18713,N_18824);
and U19090 (N_19090,N_18611,N_18711);
xnor U19091 (N_19091,N_18859,N_18733);
nor U19092 (N_19092,N_18884,N_18735);
and U19093 (N_19093,N_18701,N_18817);
nand U19094 (N_19094,N_18748,N_18756);
nor U19095 (N_19095,N_18643,N_18836);
and U19096 (N_19096,N_18777,N_18837);
nor U19097 (N_19097,N_18635,N_18785);
nor U19098 (N_19098,N_18887,N_18660);
xor U19099 (N_19099,N_18667,N_18820);
xnor U19100 (N_19100,N_18619,N_18679);
nand U19101 (N_19101,N_18701,N_18700);
nor U19102 (N_19102,N_18669,N_18769);
nand U19103 (N_19103,N_18714,N_18817);
nor U19104 (N_19104,N_18679,N_18775);
xor U19105 (N_19105,N_18863,N_18860);
and U19106 (N_19106,N_18745,N_18794);
xnor U19107 (N_19107,N_18855,N_18723);
nor U19108 (N_19108,N_18841,N_18872);
nand U19109 (N_19109,N_18748,N_18684);
and U19110 (N_19110,N_18814,N_18626);
or U19111 (N_19111,N_18862,N_18832);
nand U19112 (N_19112,N_18860,N_18783);
and U19113 (N_19113,N_18784,N_18871);
nand U19114 (N_19114,N_18666,N_18744);
nand U19115 (N_19115,N_18772,N_18760);
and U19116 (N_19116,N_18780,N_18833);
or U19117 (N_19117,N_18672,N_18810);
and U19118 (N_19118,N_18764,N_18854);
nor U19119 (N_19119,N_18737,N_18858);
and U19120 (N_19120,N_18812,N_18826);
nand U19121 (N_19121,N_18621,N_18834);
and U19122 (N_19122,N_18827,N_18807);
or U19123 (N_19123,N_18696,N_18642);
xor U19124 (N_19124,N_18732,N_18779);
nand U19125 (N_19125,N_18804,N_18630);
nor U19126 (N_19126,N_18752,N_18734);
and U19127 (N_19127,N_18707,N_18798);
nand U19128 (N_19128,N_18724,N_18842);
nor U19129 (N_19129,N_18840,N_18673);
and U19130 (N_19130,N_18701,N_18659);
nand U19131 (N_19131,N_18789,N_18804);
and U19132 (N_19132,N_18622,N_18719);
nand U19133 (N_19133,N_18615,N_18785);
and U19134 (N_19134,N_18676,N_18768);
or U19135 (N_19135,N_18687,N_18750);
nand U19136 (N_19136,N_18787,N_18804);
nor U19137 (N_19137,N_18722,N_18888);
and U19138 (N_19138,N_18603,N_18712);
xnor U19139 (N_19139,N_18617,N_18769);
xor U19140 (N_19140,N_18835,N_18695);
and U19141 (N_19141,N_18753,N_18604);
nand U19142 (N_19142,N_18800,N_18765);
nor U19143 (N_19143,N_18874,N_18823);
xnor U19144 (N_19144,N_18813,N_18698);
or U19145 (N_19145,N_18754,N_18691);
xor U19146 (N_19146,N_18635,N_18806);
nor U19147 (N_19147,N_18613,N_18737);
nand U19148 (N_19148,N_18850,N_18796);
nor U19149 (N_19149,N_18708,N_18742);
nor U19150 (N_19150,N_18630,N_18645);
xnor U19151 (N_19151,N_18684,N_18730);
and U19152 (N_19152,N_18694,N_18755);
or U19153 (N_19153,N_18783,N_18760);
xor U19154 (N_19154,N_18798,N_18827);
or U19155 (N_19155,N_18701,N_18804);
nor U19156 (N_19156,N_18737,N_18854);
xor U19157 (N_19157,N_18806,N_18798);
nor U19158 (N_19158,N_18688,N_18692);
xor U19159 (N_19159,N_18709,N_18811);
nand U19160 (N_19160,N_18628,N_18658);
and U19161 (N_19161,N_18683,N_18822);
and U19162 (N_19162,N_18676,N_18803);
and U19163 (N_19163,N_18841,N_18637);
or U19164 (N_19164,N_18636,N_18891);
nor U19165 (N_19165,N_18821,N_18847);
and U19166 (N_19166,N_18776,N_18722);
nor U19167 (N_19167,N_18657,N_18634);
nor U19168 (N_19168,N_18884,N_18621);
nor U19169 (N_19169,N_18893,N_18627);
nand U19170 (N_19170,N_18796,N_18825);
nand U19171 (N_19171,N_18744,N_18746);
nor U19172 (N_19172,N_18796,N_18866);
nor U19173 (N_19173,N_18697,N_18834);
xor U19174 (N_19174,N_18829,N_18736);
nand U19175 (N_19175,N_18772,N_18776);
and U19176 (N_19176,N_18655,N_18774);
nand U19177 (N_19177,N_18806,N_18692);
xor U19178 (N_19178,N_18883,N_18862);
nor U19179 (N_19179,N_18701,N_18846);
xor U19180 (N_19180,N_18767,N_18642);
or U19181 (N_19181,N_18825,N_18699);
nand U19182 (N_19182,N_18871,N_18802);
nor U19183 (N_19183,N_18634,N_18813);
or U19184 (N_19184,N_18879,N_18657);
xor U19185 (N_19185,N_18769,N_18615);
xor U19186 (N_19186,N_18823,N_18615);
and U19187 (N_19187,N_18665,N_18801);
nand U19188 (N_19188,N_18791,N_18869);
nor U19189 (N_19189,N_18707,N_18662);
nor U19190 (N_19190,N_18714,N_18843);
or U19191 (N_19191,N_18731,N_18834);
xor U19192 (N_19192,N_18891,N_18858);
or U19193 (N_19193,N_18784,N_18724);
nor U19194 (N_19194,N_18717,N_18801);
or U19195 (N_19195,N_18693,N_18857);
nand U19196 (N_19196,N_18874,N_18673);
nand U19197 (N_19197,N_18800,N_18753);
nor U19198 (N_19198,N_18774,N_18750);
nor U19199 (N_19199,N_18764,N_18698);
xnor U19200 (N_19200,N_19184,N_18901);
nand U19201 (N_19201,N_18962,N_18987);
and U19202 (N_19202,N_19196,N_19186);
or U19203 (N_19203,N_18906,N_18932);
nand U19204 (N_19204,N_18948,N_19032);
and U19205 (N_19205,N_19000,N_18963);
xor U19206 (N_19206,N_18970,N_19132);
and U19207 (N_19207,N_18974,N_19039);
or U19208 (N_19208,N_19021,N_19084);
and U19209 (N_19209,N_18973,N_19095);
nor U19210 (N_19210,N_19121,N_19042);
or U19211 (N_19211,N_19123,N_18950);
and U19212 (N_19212,N_18914,N_18916);
or U19213 (N_19213,N_19072,N_18910);
nand U19214 (N_19214,N_18991,N_19096);
nand U19215 (N_19215,N_18938,N_18903);
xor U19216 (N_19216,N_19080,N_19082);
nor U19217 (N_19217,N_19133,N_19136);
xor U19218 (N_19218,N_18917,N_18926);
and U19219 (N_19219,N_19116,N_18971);
nand U19220 (N_19220,N_19118,N_19185);
and U19221 (N_19221,N_19139,N_19059);
or U19222 (N_19222,N_19040,N_18992);
nor U19223 (N_19223,N_18993,N_18996);
nor U19224 (N_19224,N_19076,N_18995);
nand U19225 (N_19225,N_18953,N_19168);
nand U19226 (N_19226,N_19007,N_18961);
and U19227 (N_19227,N_19195,N_18942);
nor U19228 (N_19228,N_18928,N_19085);
or U19229 (N_19229,N_19112,N_18960);
nand U19230 (N_19230,N_19162,N_19051);
xor U19231 (N_19231,N_18923,N_19131);
and U19232 (N_19232,N_18977,N_19108);
or U19233 (N_19233,N_19013,N_19143);
xnor U19234 (N_19234,N_19077,N_18984);
or U19235 (N_19235,N_19026,N_19078);
nand U19236 (N_19236,N_19097,N_19089);
xor U19237 (N_19237,N_19151,N_19134);
or U19238 (N_19238,N_19154,N_18935);
nor U19239 (N_19239,N_19098,N_19020);
nor U19240 (N_19240,N_18913,N_19142);
or U19241 (N_19241,N_18997,N_18967);
nor U19242 (N_19242,N_19187,N_19093);
nand U19243 (N_19243,N_19050,N_18955);
xnor U19244 (N_19244,N_19144,N_19179);
or U19245 (N_19245,N_18933,N_19062);
nor U19246 (N_19246,N_19073,N_18975);
and U19247 (N_19247,N_19147,N_18949);
and U19248 (N_19248,N_19170,N_18947);
nand U19249 (N_19249,N_19054,N_18966);
or U19250 (N_19250,N_19028,N_19109);
or U19251 (N_19251,N_19126,N_18936);
xor U19252 (N_19252,N_19037,N_19107);
or U19253 (N_19253,N_19065,N_18907);
or U19254 (N_19254,N_18994,N_18941);
xnor U19255 (N_19255,N_19010,N_18986);
xor U19256 (N_19256,N_19091,N_19014);
or U19257 (N_19257,N_19018,N_18927);
nand U19258 (N_19258,N_19114,N_19002);
nand U19259 (N_19259,N_18912,N_19060);
nand U19260 (N_19260,N_19174,N_19180);
nand U19261 (N_19261,N_19177,N_19197);
or U19262 (N_19262,N_18954,N_19111);
nor U19263 (N_19263,N_19130,N_18924);
and U19264 (N_19264,N_18981,N_19075);
nor U19265 (N_19265,N_19066,N_19067);
nand U19266 (N_19266,N_19048,N_19165);
nand U19267 (N_19267,N_19155,N_19074);
nor U19268 (N_19268,N_18976,N_19004);
nor U19269 (N_19269,N_18908,N_19056);
xor U19270 (N_19270,N_19188,N_18968);
nand U19271 (N_19271,N_19199,N_18940);
xnor U19272 (N_19272,N_19156,N_18952);
or U19273 (N_19273,N_19083,N_19024);
nand U19274 (N_19274,N_19183,N_19079);
xor U19275 (N_19275,N_18902,N_19005);
xor U19276 (N_19276,N_19081,N_19103);
nor U19277 (N_19277,N_19058,N_19159);
or U19278 (N_19278,N_18944,N_19057);
or U19279 (N_19279,N_19046,N_19041);
or U19280 (N_19280,N_18909,N_19069);
nand U19281 (N_19281,N_19157,N_19163);
nand U19282 (N_19282,N_19172,N_19015);
xnor U19283 (N_19283,N_18919,N_19119);
or U19284 (N_19284,N_18979,N_18985);
nor U19285 (N_19285,N_18930,N_19149);
or U19286 (N_19286,N_19124,N_19053);
nor U19287 (N_19287,N_18980,N_19104);
or U19288 (N_19288,N_19164,N_19125);
or U19289 (N_19289,N_19176,N_19129);
or U19290 (N_19290,N_19106,N_18946);
nand U19291 (N_19291,N_19101,N_19063);
nand U19292 (N_19292,N_19140,N_19055);
or U19293 (N_19293,N_19158,N_19094);
or U19294 (N_19294,N_19120,N_18945);
or U19295 (N_19295,N_19017,N_19001);
nand U19296 (N_19296,N_19182,N_18957);
and U19297 (N_19297,N_19064,N_19099);
and U19298 (N_19298,N_19047,N_18988);
nor U19299 (N_19299,N_18989,N_19027);
or U19300 (N_19300,N_19193,N_19150);
nor U19301 (N_19301,N_19113,N_18904);
nand U19302 (N_19302,N_19194,N_19045);
xnor U19303 (N_19303,N_19138,N_19023);
and U19304 (N_19304,N_19038,N_19016);
or U19305 (N_19305,N_18990,N_19044);
and U19306 (N_19306,N_19006,N_19178);
and U19307 (N_19307,N_19148,N_18925);
nor U19308 (N_19308,N_18972,N_19167);
nand U19309 (N_19309,N_19122,N_18900);
and U19310 (N_19310,N_18999,N_18956);
xor U19311 (N_19311,N_18964,N_19146);
or U19312 (N_19312,N_18943,N_19086);
nand U19313 (N_19313,N_19135,N_19190);
or U19314 (N_19314,N_19189,N_19019);
and U19315 (N_19315,N_19191,N_18937);
xnor U19316 (N_19316,N_18998,N_19173);
nand U19317 (N_19317,N_19100,N_19145);
nand U19318 (N_19318,N_19070,N_19030);
nand U19319 (N_19319,N_19035,N_19029);
nand U19320 (N_19320,N_19166,N_19033);
and U19321 (N_19321,N_18939,N_18918);
and U19322 (N_19322,N_19052,N_19031);
xnor U19323 (N_19323,N_18921,N_19087);
xor U19324 (N_19324,N_19012,N_18931);
and U19325 (N_19325,N_19043,N_19025);
and U19326 (N_19326,N_18922,N_18905);
nand U19327 (N_19327,N_18934,N_19192);
or U19328 (N_19328,N_19022,N_19169);
nor U19329 (N_19329,N_19115,N_19068);
or U19330 (N_19330,N_19105,N_19034);
and U19331 (N_19331,N_19153,N_19071);
or U19332 (N_19332,N_18958,N_19036);
xnor U19333 (N_19333,N_19137,N_18951);
nor U19334 (N_19334,N_19011,N_19061);
or U19335 (N_19335,N_19049,N_19181);
or U19336 (N_19336,N_19175,N_19110);
nand U19337 (N_19337,N_18915,N_19088);
and U19338 (N_19338,N_18929,N_18982);
nor U19339 (N_19339,N_19171,N_18969);
and U19340 (N_19340,N_19161,N_19198);
xnor U19341 (N_19341,N_19009,N_19128);
nor U19342 (N_19342,N_19160,N_19008);
nor U19343 (N_19343,N_19090,N_19127);
nor U19344 (N_19344,N_18965,N_18959);
nand U19345 (N_19345,N_18983,N_19117);
or U19346 (N_19346,N_19003,N_19152);
xnor U19347 (N_19347,N_19141,N_18911);
nand U19348 (N_19348,N_19092,N_19102);
xor U19349 (N_19349,N_18978,N_18920);
or U19350 (N_19350,N_18970,N_19151);
and U19351 (N_19351,N_19160,N_18985);
or U19352 (N_19352,N_18983,N_19112);
and U19353 (N_19353,N_19039,N_18986);
or U19354 (N_19354,N_19172,N_19165);
nand U19355 (N_19355,N_19029,N_19095);
xor U19356 (N_19356,N_19027,N_19139);
nor U19357 (N_19357,N_18941,N_19100);
and U19358 (N_19358,N_19049,N_18921);
xnor U19359 (N_19359,N_18975,N_18931);
and U19360 (N_19360,N_19047,N_19085);
xnor U19361 (N_19361,N_18970,N_19031);
nor U19362 (N_19362,N_18934,N_19156);
nand U19363 (N_19363,N_18943,N_19073);
nand U19364 (N_19364,N_18911,N_18929);
xnor U19365 (N_19365,N_18935,N_19179);
xor U19366 (N_19366,N_19102,N_19122);
and U19367 (N_19367,N_19019,N_18956);
nand U19368 (N_19368,N_19022,N_19008);
and U19369 (N_19369,N_19151,N_19096);
nand U19370 (N_19370,N_18917,N_18960);
and U19371 (N_19371,N_18948,N_18906);
nor U19372 (N_19372,N_19008,N_19018);
xor U19373 (N_19373,N_18966,N_19088);
nand U19374 (N_19374,N_18903,N_18972);
and U19375 (N_19375,N_19076,N_19050);
xnor U19376 (N_19376,N_19130,N_19076);
nand U19377 (N_19377,N_19009,N_18948);
nand U19378 (N_19378,N_19194,N_19073);
nand U19379 (N_19379,N_19040,N_18905);
nand U19380 (N_19380,N_19197,N_18957);
and U19381 (N_19381,N_18971,N_19091);
or U19382 (N_19382,N_19075,N_18923);
xor U19383 (N_19383,N_18939,N_19057);
nor U19384 (N_19384,N_18982,N_19093);
xnor U19385 (N_19385,N_19048,N_19181);
nor U19386 (N_19386,N_19138,N_18902);
nand U19387 (N_19387,N_18941,N_18916);
and U19388 (N_19388,N_19125,N_18992);
nand U19389 (N_19389,N_19006,N_19050);
xnor U19390 (N_19390,N_19085,N_18992);
and U19391 (N_19391,N_18925,N_19138);
nand U19392 (N_19392,N_18914,N_19088);
nor U19393 (N_19393,N_19101,N_19107);
xnor U19394 (N_19394,N_19012,N_18951);
or U19395 (N_19395,N_19088,N_19125);
nor U19396 (N_19396,N_19193,N_18987);
and U19397 (N_19397,N_18997,N_19078);
nor U19398 (N_19398,N_19133,N_19195);
xor U19399 (N_19399,N_19132,N_18932);
nor U19400 (N_19400,N_19015,N_19157);
nor U19401 (N_19401,N_19197,N_18982);
and U19402 (N_19402,N_19173,N_18909);
nor U19403 (N_19403,N_18956,N_18982);
xor U19404 (N_19404,N_18928,N_19026);
nand U19405 (N_19405,N_19006,N_19045);
xnor U19406 (N_19406,N_19197,N_19087);
xnor U19407 (N_19407,N_18981,N_19159);
xor U19408 (N_19408,N_18909,N_18941);
nand U19409 (N_19409,N_19136,N_18971);
nor U19410 (N_19410,N_18911,N_18943);
xor U19411 (N_19411,N_19021,N_18965);
and U19412 (N_19412,N_19078,N_19159);
nor U19413 (N_19413,N_18997,N_18941);
xnor U19414 (N_19414,N_19076,N_19113);
and U19415 (N_19415,N_19046,N_19095);
or U19416 (N_19416,N_18959,N_18977);
and U19417 (N_19417,N_19006,N_19067);
nor U19418 (N_19418,N_18963,N_18934);
and U19419 (N_19419,N_18935,N_19164);
xnor U19420 (N_19420,N_19176,N_18943);
or U19421 (N_19421,N_19134,N_18934);
or U19422 (N_19422,N_19135,N_19103);
nor U19423 (N_19423,N_19145,N_18939);
and U19424 (N_19424,N_18954,N_18957);
nor U19425 (N_19425,N_18924,N_18900);
and U19426 (N_19426,N_18999,N_18971);
nand U19427 (N_19427,N_19165,N_19057);
nand U19428 (N_19428,N_19075,N_18909);
nor U19429 (N_19429,N_19099,N_19015);
xor U19430 (N_19430,N_19024,N_19127);
nor U19431 (N_19431,N_18919,N_19076);
and U19432 (N_19432,N_19194,N_19140);
or U19433 (N_19433,N_18935,N_19183);
nor U19434 (N_19434,N_19035,N_19039);
nor U19435 (N_19435,N_19135,N_18997);
and U19436 (N_19436,N_18975,N_18958);
nor U19437 (N_19437,N_18963,N_18955);
nor U19438 (N_19438,N_19165,N_18991);
nand U19439 (N_19439,N_18988,N_19013);
nand U19440 (N_19440,N_19079,N_19150);
or U19441 (N_19441,N_18950,N_19109);
or U19442 (N_19442,N_19129,N_19028);
nand U19443 (N_19443,N_18911,N_19195);
nand U19444 (N_19444,N_18926,N_19067);
xnor U19445 (N_19445,N_19161,N_19036);
xor U19446 (N_19446,N_19060,N_19062);
nor U19447 (N_19447,N_18984,N_18969);
or U19448 (N_19448,N_18909,N_19018);
xnor U19449 (N_19449,N_18952,N_18930);
nor U19450 (N_19450,N_19198,N_19167);
or U19451 (N_19451,N_18902,N_18922);
nor U19452 (N_19452,N_18972,N_19076);
nor U19453 (N_19453,N_18973,N_19001);
xnor U19454 (N_19454,N_19179,N_18977);
or U19455 (N_19455,N_19072,N_19050);
xnor U19456 (N_19456,N_18988,N_19127);
and U19457 (N_19457,N_19148,N_18975);
and U19458 (N_19458,N_19022,N_18958);
nor U19459 (N_19459,N_18942,N_19073);
nor U19460 (N_19460,N_18928,N_19195);
nand U19461 (N_19461,N_19064,N_19037);
xnor U19462 (N_19462,N_18919,N_19091);
and U19463 (N_19463,N_19029,N_19057);
nor U19464 (N_19464,N_18970,N_19002);
xnor U19465 (N_19465,N_19160,N_19115);
or U19466 (N_19466,N_19130,N_18959);
or U19467 (N_19467,N_18946,N_18940);
nand U19468 (N_19468,N_19020,N_19147);
and U19469 (N_19469,N_19128,N_19081);
and U19470 (N_19470,N_19010,N_19027);
or U19471 (N_19471,N_19138,N_18945);
nor U19472 (N_19472,N_18999,N_19175);
and U19473 (N_19473,N_19162,N_19132);
nand U19474 (N_19474,N_18924,N_19153);
and U19475 (N_19475,N_19006,N_18924);
nand U19476 (N_19476,N_19010,N_18947);
nor U19477 (N_19477,N_18959,N_18951);
nor U19478 (N_19478,N_19148,N_19017);
or U19479 (N_19479,N_18911,N_18915);
and U19480 (N_19480,N_19001,N_19111);
nor U19481 (N_19481,N_18970,N_19097);
nand U19482 (N_19482,N_19178,N_18973);
nor U19483 (N_19483,N_18963,N_18935);
nand U19484 (N_19484,N_19188,N_19082);
nand U19485 (N_19485,N_19121,N_19159);
nor U19486 (N_19486,N_18977,N_19180);
nor U19487 (N_19487,N_18903,N_18901);
xnor U19488 (N_19488,N_19163,N_19190);
nor U19489 (N_19489,N_19003,N_18952);
or U19490 (N_19490,N_18966,N_19190);
nor U19491 (N_19491,N_18970,N_19030);
or U19492 (N_19492,N_19000,N_18981);
and U19493 (N_19493,N_19061,N_19052);
nand U19494 (N_19494,N_18944,N_19068);
or U19495 (N_19495,N_19060,N_19004);
xnor U19496 (N_19496,N_18921,N_19144);
or U19497 (N_19497,N_19038,N_18946);
xnor U19498 (N_19498,N_19183,N_18963);
and U19499 (N_19499,N_19096,N_19166);
xor U19500 (N_19500,N_19326,N_19476);
nand U19501 (N_19501,N_19354,N_19364);
nor U19502 (N_19502,N_19432,N_19435);
xor U19503 (N_19503,N_19417,N_19303);
or U19504 (N_19504,N_19332,N_19335);
nor U19505 (N_19505,N_19305,N_19228);
nand U19506 (N_19506,N_19203,N_19260);
xnor U19507 (N_19507,N_19406,N_19425);
xnor U19508 (N_19508,N_19499,N_19477);
nand U19509 (N_19509,N_19398,N_19208);
nor U19510 (N_19510,N_19287,N_19424);
and U19511 (N_19511,N_19248,N_19230);
nand U19512 (N_19512,N_19297,N_19347);
nand U19513 (N_19513,N_19226,N_19227);
nor U19514 (N_19514,N_19465,N_19368);
xnor U19515 (N_19515,N_19300,N_19485);
and U19516 (N_19516,N_19263,N_19244);
or U19517 (N_19517,N_19283,N_19359);
nor U19518 (N_19518,N_19223,N_19309);
nand U19519 (N_19519,N_19270,N_19420);
nand U19520 (N_19520,N_19325,N_19258);
or U19521 (N_19521,N_19386,N_19212);
xor U19522 (N_19522,N_19429,N_19371);
or U19523 (N_19523,N_19369,N_19215);
nor U19524 (N_19524,N_19357,N_19443);
nor U19525 (N_19525,N_19239,N_19261);
and U19526 (N_19526,N_19233,N_19209);
xnor U19527 (N_19527,N_19202,N_19334);
xnor U19528 (N_19528,N_19448,N_19225);
nand U19529 (N_19529,N_19346,N_19304);
and U19530 (N_19530,N_19307,N_19264);
nand U19531 (N_19531,N_19214,N_19336);
nand U19532 (N_19532,N_19454,N_19256);
xnor U19533 (N_19533,N_19404,N_19262);
and U19534 (N_19534,N_19457,N_19391);
and U19535 (N_19535,N_19421,N_19344);
nand U19536 (N_19536,N_19373,N_19277);
and U19537 (N_19537,N_19246,N_19254);
xor U19538 (N_19538,N_19489,N_19356);
or U19539 (N_19539,N_19308,N_19343);
and U19540 (N_19540,N_19461,N_19296);
xnor U19541 (N_19541,N_19313,N_19480);
and U19542 (N_19542,N_19415,N_19205);
and U19543 (N_19543,N_19383,N_19370);
and U19544 (N_19544,N_19275,N_19232);
nand U19545 (N_19545,N_19316,N_19362);
nand U19546 (N_19546,N_19353,N_19224);
nand U19547 (N_19547,N_19234,N_19387);
xor U19548 (N_19548,N_19206,N_19222);
or U19549 (N_19549,N_19449,N_19375);
or U19550 (N_19550,N_19319,N_19471);
and U19551 (N_19551,N_19492,N_19399);
nor U19552 (N_19552,N_19253,N_19295);
nor U19553 (N_19553,N_19324,N_19470);
or U19554 (N_19554,N_19385,N_19318);
nand U19555 (N_19555,N_19446,N_19482);
nand U19556 (N_19556,N_19245,N_19410);
nor U19557 (N_19557,N_19444,N_19411);
and U19558 (N_19558,N_19452,N_19229);
nor U19559 (N_19559,N_19299,N_19496);
nand U19560 (N_19560,N_19486,N_19413);
and U19561 (N_19561,N_19345,N_19259);
and U19562 (N_19562,N_19434,N_19216);
and U19563 (N_19563,N_19294,N_19463);
nand U19564 (N_19564,N_19494,N_19393);
nor U19565 (N_19565,N_19280,N_19437);
or U19566 (N_19566,N_19498,N_19436);
xnor U19567 (N_19567,N_19451,N_19467);
nor U19568 (N_19568,N_19408,N_19221);
nor U19569 (N_19569,N_19374,N_19414);
and U19570 (N_19570,N_19442,N_19394);
or U19571 (N_19571,N_19247,N_19349);
and U19572 (N_19572,N_19407,N_19268);
nor U19573 (N_19573,N_19377,N_19487);
nand U19574 (N_19574,N_19418,N_19310);
and U19575 (N_19575,N_19323,N_19315);
nor U19576 (N_19576,N_19252,N_19472);
and U19577 (N_19577,N_19314,N_19358);
or U19578 (N_19578,N_19453,N_19372);
and U19579 (N_19579,N_19269,N_19338);
nor U19580 (N_19580,N_19378,N_19389);
or U19581 (N_19581,N_19200,N_19478);
nand U19582 (N_19582,N_19322,N_19363);
nor U19583 (N_19583,N_19381,N_19328);
nand U19584 (N_19584,N_19423,N_19455);
nor U19585 (N_19585,N_19367,N_19340);
xnor U19586 (N_19586,N_19218,N_19257);
xor U19587 (N_19587,N_19348,N_19337);
xnor U19588 (N_19588,N_19456,N_19272);
xor U19589 (N_19589,N_19361,N_19382);
nor U19590 (N_19590,N_19416,N_19213);
or U19591 (N_19591,N_19409,N_19204);
xnor U19592 (N_19592,N_19400,N_19293);
nor U19593 (N_19593,N_19458,N_19290);
nand U19594 (N_19594,N_19462,N_19475);
and U19595 (N_19595,N_19430,N_19441);
xor U19596 (N_19596,N_19438,N_19401);
nand U19597 (N_19597,N_19431,N_19392);
xnor U19598 (N_19598,N_19271,N_19330);
nor U19599 (N_19599,N_19220,N_19279);
nand U19600 (N_19600,N_19238,N_19466);
and U19601 (N_19601,N_19428,N_19274);
xor U19602 (N_19602,N_19365,N_19320);
xor U19603 (N_19603,N_19288,N_19445);
and U19604 (N_19604,N_19286,N_19265);
nor U19605 (N_19605,N_19481,N_19291);
or U19606 (N_19606,N_19267,N_19249);
nor U19607 (N_19607,N_19495,N_19474);
nand U19608 (N_19608,N_19311,N_19281);
xnor U19609 (N_19609,N_19376,N_19459);
nor U19610 (N_19610,N_19329,N_19339);
and U19611 (N_19611,N_19366,N_19384);
or U19612 (N_19612,N_19342,N_19278);
xnor U19613 (N_19613,N_19292,N_19422);
nor U19614 (N_19614,N_19201,N_19317);
nand U19615 (N_19615,N_19289,N_19396);
nand U19616 (N_19616,N_19266,N_19360);
or U19617 (N_19617,N_19243,N_19397);
and U19618 (N_19618,N_19427,N_19439);
or U19619 (N_19619,N_19473,N_19219);
and U19620 (N_19620,N_19468,N_19211);
nor U19621 (N_19621,N_19231,N_19447);
nor U19622 (N_19622,N_19355,N_19255);
nor U19623 (N_19623,N_19237,N_19491);
nor U19624 (N_19624,N_19235,N_19273);
xor U19625 (N_19625,N_19479,N_19460);
xor U19626 (N_19626,N_19433,N_19352);
nor U19627 (N_19627,N_19321,N_19379);
and U19628 (N_19628,N_19497,N_19236);
and U19629 (N_19629,N_19405,N_19412);
and U19630 (N_19630,N_19440,N_19390);
xnor U19631 (N_19631,N_19250,N_19282);
and U19632 (N_19632,N_19341,N_19240);
nor U19633 (N_19633,N_19331,N_19302);
nand U19634 (N_19634,N_19301,N_19284);
or U19635 (N_19635,N_19312,N_19402);
and U19636 (N_19636,N_19484,N_19488);
and U19637 (N_19637,N_19207,N_19298);
xor U19638 (N_19638,N_19490,N_19251);
nand U19639 (N_19639,N_19327,N_19388);
xor U19640 (N_19640,N_19285,N_19242);
or U19641 (N_19641,N_19276,N_19419);
xor U19642 (N_19642,N_19483,N_19450);
nand U19643 (N_19643,N_19464,N_19380);
nand U19644 (N_19644,N_19469,N_19403);
or U19645 (N_19645,N_19210,N_19351);
nor U19646 (N_19646,N_19241,N_19350);
nand U19647 (N_19647,N_19395,N_19306);
nor U19648 (N_19648,N_19493,N_19426);
nand U19649 (N_19649,N_19217,N_19333);
nand U19650 (N_19650,N_19304,N_19481);
or U19651 (N_19651,N_19374,N_19332);
nand U19652 (N_19652,N_19440,N_19498);
nand U19653 (N_19653,N_19395,N_19491);
nor U19654 (N_19654,N_19280,N_19326);
or U19655 (N_19655,N_19386,N_19345);
and U19656 (N_19656,N_19384,N_19472);
nor U19657 (N_19657,N_19320,N_19242);
xnor U19658 (N_19658,N_19264,N_19447);
and U19659 (N_19659,N_19493,N_19323);
nor U19660 (N_19660,N_19265,N_19280);
and U19661 (N_19661,N_19327,N_19236);
xnor U19662 (N_19662,N_19247,N_19298);
and U19663 (N_19663,N_19478,N_19234);
or U19664 (N_19664,N_19218,N_19232);
and U19665 (N_19665,N_19211,N_19296);
and U19666 (N_19666,N_19207,N_19454);
xor U19667 (N_19667,N_19445,N_19292);
or U19668 (N_19668,N_19468,N_19446);
or U19669 (N_19669,N_19237,N_19313);
or U19670 (N_19670,N_19470,N_19357);
or U19671 (N_19671,N_19415,N_19405);
xnor U19672 (N_19672,N_19324,N_19301);
xnor U19673 (N_19673,N_19241,N_19227);
xnor U19674 (N_19674,N_19406,N_19367);
nor U19675 (N_19675,N_19439,N_19333);
and U19676 (N_19676,N_19432,N_19236);
or U19677 (N_19677,N_19434,N_19297);
nor U19678 (N_19678,N_19454,N_19486);
xnor U19679 (N_19679,N_19280,N_19241);
and U19680 (N_19680,N_19445,N_19247);
xor U19681 (N_19681,N_19497,N_19419);
and U19682 (N_19682,N_19437,N_19481);
nand U19683 (N_19683,N_19342,N_19358);
and U19684 (N_19684,N_19201,N_19419);
xor U19685 (N_19685,N_19306,N_19308);
or U19686 (N_19686,N_19235,N_19448);
nand U19687 (N_19687,N_19474,N_19379);
nand U19688 (N_19688,N_19429,N_19202);
nand U19689 (N_19689,N_19314,N_19428);
and U19690 (N_19690,N_19352,N_19323);
or U19691 (N_19691,N_19385,N_19338);
xor U19692 (N_19692,N_19429,N_19475);
and U19693 (N_19693,N_19488,N_19443);
or U19694 (N_19694,N_19345,N_19229);
nor U19695 (N_19695,N_19477,N_19401);
nor U19696 (N_19696,N_19440,N_19288);
nand U19697 (N_19697,N_19214,N_19421);
nor U19698 (N_19698,N_19279,N_19464);
and U19699 (N_19699,N_19351,N_19427);
and U19700 (N_19700,N_19274,N_19335);
xnor U19701 (N_19701,N_19232,N_19472);
xor U19702 (N_19702,N_19342,N_19211);
xnor U19703 (N_19703,N_19320,N_19310);
nand U19704 (N_19704,N_19283,N_19392);
xnor U19705 (N_19705,N_19470,N_19333);
and U19706 (N_19706,N_19303,N_19411);
nor U19707 (N_19707,N_19480,N_19349);
xnor U19708 (N_19708,N_19215,N_19433);
or U19709 (N_19709,N_19366,N_19279);
and U19710 (N_19710,N_19490,N_19338);
nand U19711 (N_19711,N_19424,N_19413);
and U19712 (N_19712,N_19447,N_19244);
nor U19713 (N_19713,N_19347,N_19445);
or U19714 (N_19714,N_19322,N_19468);
and U19715 (N_19715,N_19389,N_19347);
nor U19716 (N_19716,N_19430,N_19493);
xnor U19717 (N_19717,N_19265,N_19211);
and U19718 (N_19718,N_19295,N_19402);
nand U19719 (N_19719,N_19467,N_19332);
nor U19720 (N_19720,N_19214,N_19305);
nand U19721 (N_19721,N_19414,N_19331);
nor U19722 (N_19722,N_19253,N_19308);
xor U19723 (N_19723,N_19482,N_19413);
nand U19724 (N_19724,N_19364,N_19428);
nand U19725 (N_19725,N_19241,N_19289);
and U19726 (N_19726,N_19435,N_19393);
nand U19727 (N_19727,N_19319,N_19241);
xnor U19728 (N_19728,N_19282,N_19232);
nand U19729 (N_19729,N_19239,N_19374);
and U19730 (N_19730,N_19331,N_19326);
or U19731 (N_19731,N_19303,N_19243);
and U19732 (N_19732,N_19219,N_19497);
or U19733 (N_19733,N_19218,N_19465);
nand U19734 (N_19734,N_19223,N_19326);
or U19735 (N_19735,N_19278,N_19493);
nor U19736 (N_19736,N_19258,N_19226);
nor U19737 (N_19737,N_19386,N_19450);
or U19738 (N_19738,N_19412,N_19426);
and U19739 (N_19739,N_19380,N_19482);
xor U19740 (N_19740,N_19249,N_19261);
xnor U19741 (N_19741,N_19411,N_19218);
nor U19742 (N_19742,N_19378,N_19265);
xor U19743 (N_19743,N_19486,N_19480);
or U19744 (N_19744,N_19270,N_19259);
and U19745 (N_19745,N_19203,N_19386);
and U19746 (N_19746,N_19240,N_19289);
nand U19747 (N_19747,N_19443,N_19479);
nor U19748 (N_19748,N_19441,N_19434);
nor U19749 (N_19749,N_19371,N_19448);
or U19750 (N_19750,N_19426,N_19491);
xnor U19751 (N_19751,N_19395,N_19285);
xnor U19752 (N_19752,N_19353,N_19402);
xnor U19753 (N_19753,N_19378,N_19398);
and U19754 (N_19754,N_19483,N_19499);
and U19755 (N_19755,N_19264,N_19237);
and U19756 (N_19756,N_19228,N_19458);
or U19757 (N_19757,N_19348,N_19216);
nor U19758 (N_19758,N_19272,N_19221);
or U19759 (N_19759,N_19337,N_19461);
nor U19760 (N_19760,N_19270,N_19447);
xnor U19761 (N_19761,N_19388,N_19294);
and U19762 (N_19762,N_19440,N_19327);
or U19763 (N_19763,N_19450,N_19330);
nand U19764 (N_19764,N_19470,N_19275);
and U19765 (N_19765,N_19242,N_19316);
nand U19766 (N_19766,N_19304,N_19439);
and U19767 (N_19767,N_19475,N_19339);
xor U19768 (N_19768,N_19432,N_19263);
or U19769 (N_19769,N_19449,N_19467);
or U19770 (N_19770,N_19305,N_19476);
xnor U19771 (N_19771,N_19421,N_19413);
or U19772 (N_19772,N_19386,N_19483);
and U19773 (N_19773,N_19421,N_19210);
nand U19774 (N_19774,N_19383,N_19451);
and U19775 (N_19775,N_19406,N_19395);
or U19776 (N_19776,N_19341,N_19239);
and U19777 (N_19777,N_19474,N_19335);
xnor U19778 (N_19778,N_19246,N_19466);
xor U19779 (N_19779,N_19219,N_19372);
xor U19780 (N_19780,N_19212,N_19369);
and U19781 (N_19781,N_19374,N_19329);
nand U19782 (N_19782,N_19277,N_19257);
nand U19783 (N_19783,N_19311,N_19372);
or U19784 (N_19784,N_19368,N_19309);
nand U19785 (N_19785,N_19440,N_19215);
nand U19786 (N_19786,N_19329,N_19443);
nand U19787 (N_19787,N_19350,N_19453);
nand U19788 (N_19788,N_19277,N_19263);
or U19789 (N_19789,N_19402,N_19395);
nand U19790 (N_19790,N_19225,N_19231);
and U19791 (N_19791,N_19293,N_19304);
or U19792 (N_19792,N_19339,N_19424);
xor U19793 (N_19793,N_19254,N_19303);
nor U19794 (N_19794,N_19324,N_19234);
nor U19795 (N_19795,N_19238,N_19332);
and U19796 (N_19796,N_19478,N_19445);
and U19797 (N_19797,N_19494,N_19264);
nand U19798 (N_19798,N_19428,N_19395);
nand U19799 (N_19799,N_19435,N_19410);
and U19800 (N_19800,N_19671,N_19635);
or U19801 (N_19801,N_19713,N_19677);
nand U19802 (N_19802,N_19649,N_19732);
and U19803 (N_19803,N_19669,N_19604);
and U19804 (N_19804,N_19772,N_19799);
xor U19805 (N_19805,N_19710,N_19611);
nand U19806 (N_19806,N_19720,N_19629);
nand U19807 (N_19807,N_19784,N_19587);
and U19808 (N_19808,N_19765,N_19667);
xor U19809 (N_19809,N_19771,N_19688);
nand U19810 (N_19810,N_19634,N_19500);
nor U19811 (N_19811,N_19699,N_19514);
nor U19812 (N_19812,N_19727,N_19549);
and U19813 (N_19813,N_19597,N_19664);
xnor U19814 (N_19814,N_19636,N_19749);
nand U19815 (N_19815,N_19550,N_19542);
or U19816 (N_19816,N_19525,N_19659);
xnor U19817 (N_19817,N_19683,N_19769);
and U19818 (N_19818,N_19654,N_19601);
nor U19819 (N_19819,N_19726,N_19616);
and U19820 (N_19820,N_19776,N_19589);
xnor U19821 (N_19821,N_19546,N_19735);
nand U19822 (N_19822,N_19739,N_19666);
nand U19823 (N_19823,N_19755,N_19738);
and U19824 (N_19824,N_19540,N_19670);
and U19825 (N_19825,N_19598,N_19752);
or U19826 (N_19826,N_19529,N_19526);
nor U19827 (N_19827,N_19652,N_19674);
nor U19828 (N_19828,N_19582,N_19718);
or U19829 (N_19829,N_19531,N_19653);
or U19830 (N_19830,N_19706,N_19501);
and U19831 (N_19831,N_19703,N_19797);
nand U19832 (N_19832,N_19558,N_19621);
and U19833 (N_19833,N_19605,N_19623);
and U19834 (N_19834,N_19702,N_19719);
or U19835 (N_19835,N_19606,N_19681);
or U19836 (N_19836,N_19689,N_19651);
nor U19837 (N_19837,N_19523,N_19520);
nand U19838 (N_19838,N_19524,N_19580);
nor U19839 (N_19839,N_19705,N_19569);
nand U19840 (N_19840,N_19592,N_19599);
or U19841 (N_19841,N_19657,N_19576);
and U19842 (N_19842,N_19750,N_19764);
and U19843 (N_19843,N_19579,N_19595);
xor U19844 (N_19844,N_19741,N_19762);
or U19845 (N_19845,N_19759,N_19692);
xor U19846 (N_19846,N_19515,N_19795);
and U19847 (N_19847,N_19633,N_19655);
xor U19848 (N_19848,N_19648,N_19632);
or U19849 (N_19849,N_19602,N_19638);
and U19850 (N_19850,N_19770,N_19510);
xnor U19851 (N_19851,N_19698,N_19695);
nor U19852 (N_19852,N_19748,N_19571);
and U19853 (N_19853,N_19513,N_19734);
nand U19854 (N_19854,N_19591,N_19679);
or U19855 (N_19855,N_19608,N_19613);
nand U19856 (N_19856,N_19568,N_19562);
nand U19857 (N_19857,N_19534,N_19767);
or U19858 (N_19858,N_19675,N_19768);
and U19859 (N_19859,N_19519,N_19567);
nand U19860 (N_19860,N_19796,N_19627);
nand U19861 (N_19861,N_19701,N_19612);
and U19862 (N_19862,N_19575,N_19781);
or U19863 (N_19863,N_19662,N_19642);
and U19864 (N_19864,N_19643,N_19730);
or U19865 (N_19865,N_19573,N_19521);
and U19866 (N_19866,N_19736,N_19504);
xnor U19867 (N_19867,N_19650,N_19564);
nand U19868 (N_19868,N_19619,N_19774);
or U19869 (N_19869,N_19790,N_19584);
xor U19870 (N_19870,N_19532,N_19685);
nor U19871 (N_19871,N_19716,N_19577);
nor U19872 (N_19872,N_19754,N_19761);
nand U19873 (N_19873,N_19622,N_19660);
xor U19874 (N_19874,N_19553,N_19779);
and U19875 (N_19875,N_19773,N_19548);
nand U19876 (N_19876,N_19614,N_19618);
and U19877 (N_19877,N_19509,N_19593);
or U19878 (N_19878,N_19563,N_19615);
and U19879 (N_19879,N_19539,N_19740);
nor U19880 (N_19880,N_19556,N_19617);
nand U19881 (N_19881,N_19527,N_19731);
or U19882 (N_19882,N_19712,N_19777);
xnor U19883 (N_19883,N_19787,N_19760);
and U19884 (N_19884,N_19528,N_19782);
nand U19885 (N_19885,N_19518,N_19672);
nand U19886 (N_19886,N_19552,N_19780);
xor U19887 (N_19887,N_19537,N_19555);
nand U19888 (N_19888,N_19717,N_19574);
nor U19889 (N_19889,N_19746,N_19508);
nor U19890 (N_19890,N_19758,N_19785);
or U19891 (N_19891,N_19647,N_19756);
nor U19892 (N_19892,N_19661,N_19789);
and U19893 (N_19893,N_19714,N_19751);
nand U19894 (N_19894,N_19678,N_19742);
nor U19895 (N_19895,N_19596,N_19630);
nand U19896 (N_19896,N_19733,N_19610);
nor U19897 (N_19897,N_19792,N_19778);
nand U19898 (N_19898,N_19551,N_19530);
and U19899 (N_19899,N_19503,N_19516);
or U19900 (N_19900,N_19586,N_19644);
or U19901 (N_19901,N_19625,N_19690);
nand U19902 (N_19902,N_19691,N_19572);
or U19903 (N_19903,N_19728,N_19682);
nor U19904 (N_19904,N_19533,N_19744);
nor U19905 (N_19905,N_19570,N_19665);
and U19906 (N_19906,N_19711,N_19585);
and U19907 (N_19907,N_19561,N_19668);
or U19908 (N_19908,N_19680,N_19594);
nand U19909 (N_19909,N_19583,N_19673);
or U19910 (N_19910,N_19607,N_19517);
nor U19911 (N_19911,N_19603,N_19624);
or U19912 (N_19912,N_19757,N_19788);
or U19913 (N_19913,N_19697,N_19658);
nand U19914 (N_19914,N_19753,N_19637);
nor U19915 (N_19915,N_19544,N_19559);
or U19916 (N_19916,N_19560,N_19783);
nand U19917 (N_19917,N_19707,N_19506);
nor U19918 (N_19918,N_19538,N_19609);
nor U19919 (N_19919,N_19554,N_19696);
nor U19920 (N_19920,N_19536,N_19566);
or U19921 (N_19921,N_19715,N_19676);
nor U19922 (N_19922,N_19775,N_19763);
or U19923 (N_19923,N_19547,N_19631);
nand U19924 (N_19924,N_19724,N_19708);
and U19925 (N_19925,N_19639,N_19786);
nor U19926 (N_19926,N_19745,N_19600);
nand U19927 (N_19927,N_19522,N_19590);
nand U19928 (N_19928,N_19743,N_19628);
nand U19929 (N_19929,N_19737,N_19686);
xnor U19930 (N_19930,N_19721,N_19565);
and U19931 (N_19931,N_19578,N_19747);
nand U19932 (N_19932,N_19505,N_19729);
xnor U19933 (N_19933,N_19656,N_19535);
nor U19934 (N_19934,N_19704,N_19684);
and U19935 (N_19935,N_19507,N_19588);
and U19936 (N_19936,N_19663,N_19581);
or U19937 (N_19937,N_19693,N_19709);
or U19938 (N_19938,N_19725,N_19557);
nor U19939 (N_19939,N_19511,N_19543);
nand U19940 (N_19940,N_19700,N_19620);
nor U19941 (N_19941,N_19640,N_19541);
or U19942 (N_19942,N_19791,N_19722);
or U19943 (N_19943,N_19645,N_19794);
nor U19944 (N_19944,N_19646,N_19793);
or U19945 (N_19945,N_19798,N_19512);
nor U19946 (N_19946,N_19766,N_19687);
xnor U19947 (N_19947,N_19694,N_19641);
nand U19948 (N_19948,N_19626,N_19545);
and U19949 (N_19949,N_19723,N_19502);
or U19950 (N_19950,N_19757,N_19723);
nand U19951 (N_19951,N_19578,N_19548);
and U19952 (N_19952,N_19609,N_19563);
nand U19953 (N_19953,N_19677,N_19718);
or U19954 (N_19954,N_19535,N_19766);
nand U19955 (N_19955,N_19501,N_19765);
xor U19956 (N_19956,N_19620,N_19709);
nand U19957 (N_19957,N_19710,N_19642);
nor U19958 (N_19958,N_19696,N_19589);
xnor U19959 (N_19959,N_19663,N_19502);
or U19960 (N_19960,N_19503,N_19790);
xor U19961 (N_19961,N_19559,N_19588);
nor U19962 (N_19962,N_19532,N_19611);
nor U19963 (N_19963,N_19629,N_19537);
nand U19964 (N_19964,N_19622,N_19686);
xnor U19965 (N_19965,N_19762,N_19520);
and U19966 (N_19966,N_19693,N_19552);
and U19967 (N_19967,N_19535,N_19699);
nor U19968 (N_19968,N_19716,N_19616);
and U19969 (N_19969,N_19650,N_19727);
and U19970 (N_19970,N_19732,N_19691);
or U19971 (N_19971,N_19577,N_19509);
and U19972 (N_19972,N_19789,N_19589);
and U19973 (N_19973,N_19505,N_19587);
nor U19974 (N_19974,N_19799,N_19610);
nor U19975 (N_19975,N_19674,N_19561);
nor U19976 (N_19976,N_19769,N_19664);
xnor U19977 (N_19977,N_19643,N_19545);
nand U19978 (N_19978,N_19729,N_19570);
nor U19979 (N_19979,N_19768,N_19639);
and U19980 (N_19980,N_19665,N_19783);
or U19981 (N_19981,N_19723,N_19514);
nor U19982 (N_19982,N_19517,N_19645);
nand U19983 (N_19983,N_19698,N_19510);
xor U19984 (N_19984,N_19704,N_19652);
and U19985 (N_19985,N_19540,N_19765);
and U19986 (N_19986,N_19666,N_19796);
nand U19987 (N_19987,N_19502,N_19728);
nor U19988 (N_19988,N_19500,N_19706);
xor U19989 (N_19989,N_19775,N_19712);
nand U19990 (N_19990,N_19596,N_19564);
nand U19991 (N_19991,N_19573,N_19705);
or U19992 (N_19992,N_19581,N_19753);
xor U19993 (N_19993,N_19514,N_19668);
xnor U19994 (N_19994,N_19621,N_19761);
or U19995 (N_19995,N_19643,N_19527);
or U19996 (N_19996,N_19563,N_19709);
or U19997 (N_19997,N_19793,N_19654);
xor U19998 (N_19998,N_19614,N_19686);
xnor U19999 (N_19999,N_19698,N_19675);
and U20000 (N_20000,N_19630,N_19660);
or U20001 (N_20001,N_19637,N_19717);
xnor U20002 (N_20002,N_19727,N_19512);
nor U20003 (N_20003,N_19719,N_19654);
nand U20004 (N_20004,N_19529,N_19754);
nor U20005 (N_20005,N_19708,N_19600);
and U20006 (N_20006,N_19517,N_19774);
xor U20007 (N_20007,N_19720,N_19553);
nor U20008 (N_20008,N_19589,N_19590);
nor U20009 (N_20009,N_19623,N_19629);
xnor U20010 (N_20010,N_19623,N_19544);
xor U20011 (N_20011,N_19502,N_19783);
xor U20012 (N_20012,N_19700,N_19667);
xor U20013 (N_20013,N_19703,N_19634);
nor U20014 (N_20014,N_19607,N_19698);
or U20015 (N_20015,N_19652,N_19760);
and U20016 (N_20016,N_19523,N_19641);
xor U20017 (N_20017,N_19549,N_19728);
xor U20018 (N_20018,N_19509,N_19676);
nor U20019 (N_20019,N_19507,N_19799);
nand U20020 (N_20020,N_19541,N_19754);
nor U20021 (N_20021,N_19602,N_19624);
or U20022 (N_20022,N_19662,N_19748);
or U20023 (N_20023,N_19580,N_19655);
and U20024 (N_20024,N_19565,N_19566);
or U20025 (N_20025,N_19599,N_19785);
nand U20026 (N_20026,N_19729,N_19681);
nor U20027 (N_20027,N_19555,N_19595);
and U20028 (N_20028,N_19674,N_19576);
and U20029 (N_20029,N_19648,N_19707);
nand U20030 (N_20030,N_19637,N_19766);
and U20031 (N_20031,N_19694,N_19645);
xor U20032 (N_20032,N_19616,N_19558);
nand U20033 (N_20033,N_19667,N_19723);
and U20034 (N_20034,N_19579,N_19728);
and U20035 (N_20035,N_19605,N_19517);
and U20036 (N_20036,N_19709,N_19647);
nor U20037 (N_20037,N_19526,N_19681);
and U20038 (N_20038,N_19648,N_19743);
and U20039 (N_20039,N_19615,N_19764);
and U20040 (N_20040,N_19707,N_19509);
nor U20041 (N_20041,N_19601,N_19679);
or U20042 (N_20042,N_19538,N_19582);
xor U20043 (N_20043,N_19512,N_19658);
nor U20044 (N_20044,N_19554,N_19730);
and U20045 (N_20045,N_19693,N_19781);
or U20046 (N_20046,N_19611,N_19620);
or U20047 (N_20047,N_19578,N_19724);
xnor U20048 (N_20048,N_19638,N_19560);
xnor U20049 (N_20049,N_19569,N_19524);
xor U20050 (N_20050,N_19572,N_19526);
xor U20051 (N_20051,N_19584,N_19558);
xnor U20052 (N_20052,N_19505,N_19573);
nand U20053 (N_20053,N_19558,N_19759);
nor U20054 (N_20054,N_19647,N_19567);
or U20055 (N_20055,N_19582,N_19738);
nor U20056 (N_20056,N_19784,N_19656);
or U20057 (N_20057,N_19606,N_19609);
nand U20058 (N_20058,N_19589,N_19522);
and U20059 (N_20059,N_19734,N_19798);
xnor U20060 (N_20060,N_19557,N_19764);
or U20061 (N_20061,N_19685,N_19799);
and U20062 (N_20062,N_19776,N_19504);
nor U20063 (N_20063,N_19600,N_19679);
xor U20064 (N_20064,N_19614,N_19741);
nor U20065 (N_20065,N_19611,N_19725);
nand U20066 (N_20066,N_19501,N_19609);
nor U20067 (N_20067,N_19655,N_19603);
and U20068 (N_20068,N_19724,N_19758);
nand U20069 (N_20069,N_19724,N_19682);
or U20070 (N_20070,N_19714,N_19663);
and U20071 (N_20071,N_19692,N_19502);
xnor U20072 (N_20072,N_19716,N_19798);
or U20073 (N_20073,N_19603,N_19618);
and U20074 (N_20074,N_19606,N_19572);
nor U20075 (N_20075,N_19620,N_19694);
nand U20076 (N_20076,N_19762,N_19745);
nor U20077 (N_20077,N_19565,N_19673);
or U20078 (N_20078,N_19599,N_19600);
and U20079 (N_20079,N_19543,N_19504);
xnor U20080 (N_20080,N_19673,N_19555);
nor U20081 (N_20081,N_19713,N_19717);
nand U20082 (N_20082,N_19585,N_19784);
nand U20083 (N_20083,N_19617,N_19549);
nand U20084 (N_20084,N_19765,N_19715);
nor U20085 (N_20085,N_19569,N_19682);
or U20086 (N_20086,N_19696,N_19673);
or U20087 (N_20087,N_19562,N_19607);
nor U20088 (N_20088,N_19536,N_19587);
nor U20089 (N_20089,N_19574,N_19660);
nor U20090 (N_20090,N_19788,N_19699);
xor U20091 (N_20091,N_19598,N_19525);
xor U20092 (N_20092,N_19742,N_19775);
and U20093 (N_20093,N_19600,N_19511);
nand U20094 (N_20094,N_19760,N_19519);
xnor U20095 (N_20095,N_19596,N_19676);
or U20096 (N_20096,N_19659,N_19778);
nand U20097 (N_20097,N_19745,N_19580);
nand U20098 (N_20098,N_19693,N_19758);
nor U20099 (N_20099,N_19673,N_19647);
nor U20100 (N_20100,N_19854,N_19951);
nand U20101 (N_20101,N_19805,N_19844);
xor U20102 (N_20102,N_19968,N_19959);
or U20103 (N_20103,N_19992,N_19808);
and U20104 (N_20104,N_19838,N_19975);
nand U20105 (N_20105,N_19956,N_19803);
nor U20106 (N_20106,N_19878,N_20075);
or U20107 (N_20107,N_19877,N_19866);
nor U20108 (N_20108,N_19933,N_19873);
or U20109 (N_20109,N_19934,N_19855);
or U20110 (N_20110,N_20005,N_20049);
nor U20111 (N_20111,N_19895,N_20002);
xor U20112 (N_20112,N_20090,N_20076);
nand U20113 (N_20113,N_19811,N_19955);
or U20114 (N_20114,N_19837,N_20045);
or U20115 (N_20115,N_20020,N_19957);
nand U20116 (N_20116,N_19929,N_19804);
xnor U20117 (N_20117,N_20099,N_20070);
nand U20118 (N_20118,N_19867,N_19807);
or U20119 (N_20119,N_19941,N_19919);
nand U20120 (N_20120,N_19857,N_19864);
and U20121 (N_20121,N_19853,N_19850);
nor U20122 (N_20122,N_20023,N_19823);
xor U20123 (N_20123,N_19982,N_20052);
or U20124 (N_20124,N_19921,N_20061);
and U20125 (N_20125,N_19817,N_19818);
and U20126 (N_20126,N_19827,N_19868);
or U20127 (N_20127,N_19986,N_19926);
and U20128 (N_20128,N_19860,N_20088);
nor U20129 (N_20129,N_20035,N_19922);
nand U20130 (N_20130,N_20067,N_20078);
nor U20131 (N_20131,N_19829,N_19801);
or U20132 (N_20132,N_19964,N_20072);
nor U20133 (N_20133,N_20096,N_19871);
xnor U20134 (N_20134,N_20058,N_20068);
or U20135 (N_20135,N_19961,N_19872);
and U20136 (N_20136,N_20026,N_20039);
nand U20137 (N_20137,N_20094,N_19820);
nand U20138 (N_20138,N_19812,N_20011);
nand U20139 (N_20139,N_19983,N_19996);
xnor U20140 (N_20140,N_20032,N_20007);
nor U20141 (N_20141,N_19974,N_19858);
xnor U20142 (N_20142,N_19870,N_19874);
nand U20143 (N_20143,N_19910,N_20069);
and U20144 (N_20144,N_20051,N_20015);
or U20145 (N_20145,N_19980,N_20042);
nand U20146 (N_20146,N_20065,N_19847);
xnor U20147 (N_20147,N_19806,N_20037);
nor U20148 (N_20148,N_19846,N_19948);
and U20149 (N_20149,N_19937,N_19843);
or U20150 (N_20150,N_20062,N_19822);
nand U20151 (N_20151,N_19946,N_20054);
nand U20152 (N_20152,N_19966,N_20050);
nor U20153 (N_20153,N_20055,N_20093);
nand U20154 (N_20154,N_19913,N_19840);
nor U20155 (N_20155,N_19891,N_20041);
or U20156 (N_20156,N_20074,N_19832);
nor U20157 (N_20157,N_19898,N_20073);
or U20158 (N_20158,N_19953,N_19886);
or U20159 (N_20159,N_19879,N_20031);
nor U20160 (N_20160,N_20043,N_19971);
or U20161 (N_20161,N_19821,N_20008);
nand U20162 (N_20162,N_19965,N_19816);
nor U20163 (N_20163,N_19972,N_19899);
nand U20164 (N_20164,N_19893,N_20013);
nand U20165 (N_20165,N_19912,N_19826);
xor U20166 (N_20166,N_20047,N_19813);
or U20167 (N_20167,N_19936,N_19875);
or U20168 (N_20168,N_19939,N_20085);
or U20169 (N_20169,N_19869,N_19828);
xnor U20170 (N_20170,N_19931,N_19928);
nand U20171 (N_20171,N_19800,N_19954);
or U20172 (N_20172,N_20040,N_20029);
and U20173 (N_20173,N_20025,N_19839);
nand U20174 (N_20174,N_20095,N_19920);
and U20175 (N_20175,N_20048,N_20071);
and U20176 (N_20176,N_19845,N_20046);
or U20177 (N_20177,N_19810,N_20080);
and U20178 (N_20178,N_20028,N_19815);
xor U20179 (N_20179,N_20038,N_19930);
and U20180 (N_20180,N_19962,N_20036);
or U20181 (N_20181,N_19915,N_19841);
nand U20182 (N_20182,N_20084,N_19981);
nand U20183 (N_20183,N_20056,N_20082);
nor U20184 (N_20184,N_19825,N_20027);
nand U20185 (N_20185,N_20000,N_19882);
or U20186 (N_20186,N_19849,N_19970);
xnor U20187 (N_20187,N_19863,N_19989);
xor U20188 (N_20188,N_19947,N_19967);
xnor U20189 (N_20189,N_20087,N_19987);
nor U20190 (N_20190,N_19814,N_19990);
nor U20191 (N_20191,N_19923,N_19834);
nor U20192 (N_20192,N_20063,N_19896);
or U20193 (N_20193,N_19831,N_19925);
and U20194 (N_20194,N_19977,N_19924);
nand U20195 (N_20195,N_20014,N_19884);
nand U20196 (N_20196,N_19909,N_20081);
and U20197 (N_20197,N_20077,N_20089);
xnor U20198 (N_20198,N_19861,N_19880);
xor U20199 (N_20199,N_20091,N_19802);
xor U20200 (N_20200,N_20033,N_19979);
or U20201 (N_20201,N_19830,N_19901);
xor U20202 (N_20202,N_19976,N_20016);
nor U20203 (N_20203,N_20083,N_20079);
nand U20204 (N_20204,N_19991,N_19914);
nor U20205 (N_20205,N_19876,N_20030);
nand U20206 (N_20206,N_20034,N_19894);
and U20207 (N_20207,N_19999,N_19932);
nor U20208 (N_20208,N_19993,N_19952);
or U20209 (N_20209,N_19835,N_19942);
and U20210 (N_20210,N_19885,N_20017);
or U20211 (N_20211,N_20018,N_20019);
xor U20212 (N_20212,N_19994,N_20053);
nand U20213 (N_20213,N_19940,N_19943);
and U20214 (N_20214,N_20010,N_19935);
or U20215 (N_20215,N_19998,N_20003);
and U20216 (N_20216,N_19918,N_19978);
nand U20217 (N_20217,N_20021,N_19950);
and U20218 (N_20218,N_20097,N_19958);
or U20219 (N_20219,N_19963,N_19960);
or U20220 (N_20220,N_19907,N_19865);
xor U20221 (N_20221,N_19988,N_19856);
xnor U20222 (N_20222,N_19809,N_19949);
or U20223 (N_20223,N_19905,N_20024);
xor U20224 (N_20224,N_19906,N_19881);
nor U20225 (N_20225,N_19917,N_19851);
and U20226 (N_20226,N_19889,N_19938);
nor U20227 (N_20227,N_20059,N_19944);
and U20228 (N_20228,N_20044,N_20060);
and U20229 (N_20229,N_20001,N_19908);
and U20230 (N_20230,N_20004,N_19897);
and U20231 (N_20231,N_20057,N_19852);
or U20232 (N_20232,N_19903,N_19904);
xnor U20233 (N_20233,N_19945,N_20092);
or U20234 (N_20234,N_19916,N_19973);
nand U20235 (N_20235,N_19985,N_19836);
nor U20236 (N_20236,N_19900,N_19984);
nand U20237 (N_20237,N_19819,N_19842);
or U20238 (N_20238,N_19892,N_19911);
and U20239 (N_20239,N_19995,N_19862);
xor U20240 (N_20240,N_19902,N_20066);
nor U20241 (N_20241,N_20006,N_19969);
and U20242 (N_20242,N_19824,N_19997);
and U20243 (N_20243,N_19927,N_20086);
xor U20244 (N_20244,N_20098,N_19887);
or U20245 (N_20245,N_19890,N_20064);
and U20246 (N_20246,N_19859,N_19883);
nor U20247 (N_20247,N_20022,N_19848);
nor U20248 (N_20248,N_19833,N_20009);
xnor U20249 (N_20249,N_19888,N_20012);
nand U20250 (N_20250,N_19974,N_19837);
or U20251 (N_20251,N_20074,N_19955);
or U20252 (N_20252,N_20006,N_20063);
xor U20253 (N_20253,N_20033,N_19970);
nor U20254 (N_20254,N_20037,N_19964);
xor U20255 (N_20255,N_20012,N_19840);
nand U20256 (N_20256,N_20044,N_20069);
xnor U20257 (N_20257,N_19930,N_20094);
xnor U20258 (N_20258,N_19806,N_20073);
xor U20259 (N_20259,N_19950,N_19998);
xnor U20260 (N_20260,N_19862,N_19912);
and U20261 (N_20261,N_20049,N_20062);
nor U20262 (N_20262,N_20073,N_19876);
or U20263 (N_20263,N_19857,N_19840);
nand U20264 (N_20264,N_19858,N_19816);
and U20265 (N_20265,N_19981,N_19826);
or U20266 (N_20266,N_19970,N_19855);
or U20267 (N_20267,N_19831,N_19870);
nor U20268 (N_20268,N_19947,N_19936);
xor U20269 (N_20269,N_20023,N_19806);
and U20270 (N_20270,N_19822,N_19915);
and U20271 (N_20271,N_19921,N_19846);
or U20272 (N_20272,N_19968,N_19950);
and U20273 (N_20273,N_20075,N_19874);
nand U20274 (N_20274,N_19940,N_20098);
or U20275 (N_20275,N_19956,N_19937);
and U20276 (N_20276,N_20028,N_19819);
nor U20277 (N_20277,N_19855,N_20048);
and U20278 (N_20278,N_20088,N_19869);
nor U20279 (N_20279,N_20089,N_20063);
nand U20280 (N_20280,N_20076,N_20042);
nand U20281 (N_20281,N_20092,N_20067);
or U20282 (N_20282,N_20090,N_20009);
or U20283 (N_20283,N_20079,N_19849);
xor U20284 (N_20284,N_19963,N_19967);
or U20285 (N_20285,N_19903,N_19937);
and U20286 (N_20286,N_20066,N_19968);
xor U20287 (N_20287,N_20032,N_19995);
nor U20288 (N_20288,N_20070,N_20065);
and U20289 (N_20289,N_19846,N_19900);
nor U20290 (N_20290,N_20013,N_20031);
or U20291 (N_20291,N_19881,N_20084);
and U20292 (N_20292,N_20003,N_20064);
and U20293 (N_20293,N_19947,N_19865);
and U20294 (N_20294,N_20040,N_19966);
nand U20295 (N_20295,N_20016,N_19850);
xor U20296 (N_20296,N_19996,N_19889);
and U20297 (N_20297,N_20029,N_19898);
nand U20298 (N_20298,N_20059,N_19862);
and U20299 (N_20299,N_20096,N_20005);
and U20300 (N_20300,N_19949,N_19920);
nor U20301 (N_20301,N_19993,N_19994);
or U20302 (N_20302,N_19820,N_19949);
xnor U20303 (N_20303,N_20019,N_19937);
nor U20304 (N_20304,N_19916,N_20099);
nand U20305 (N_20305,N_19901,N_20021);
and U20306 (N_20306,N_19950,N_20008);
and U20307 (N_20307,N_20091,N_19893);
or U20308 (N_20308,N_19959,N_20044);
or U20309 (N_20309,N_20065,N_19904);
and U20310 (N_20310,N_20050,N_19918);
nand U20311 (N_20311,N_20054,N_19905);
nor U20312 (N_20312,N_19988,N_19879);
or U20313 (N_20313,N_19800,N_20074);
nor U20314 (N_20314,N_19953,N_19894);
and U20315 (N_20315,N_20099,N_19831);
nor U20316 (N_20316,N_19870,N_20015);
nand U20317 (N_20317,N_19818,N_19928);
nor U20318 (N_20318,N_19929,N_19909);
and U20319 (N_20319,N_20099,N_20077);
or U20320 (N_20320,N_20072,N_19935);
nor U20321 (N_20321,N_20003,N_19912);
and U20322 (N_20322,N_20023,N_19876);
nand U20323 (N_20323,N_19948,N_19825);
nand U20324 (N_20324,N_19805,N_19954);
xnor U20325 (N_20325,N_19879,N_20093);
xnor U20326 (N_20326,N_19991,N_19926);
xor U20327 (N_20327,N_20089,N_19933);
or U20328 (N_20328,N_20007,N_19802);
or U20329 (N_20329,N_19837,N_20063);
nand U20330 (N_20330,N_19901,N_19891);
and U20331 (N_20331,N_19898,N_20046);
or U20332 (N_20332,N_19997,N_19995);
nor U20333 (N_20333,N_20074,N_20043);
nor U20334 (N_20334,N_19922,N_19996);
nor U20335 (N_20335,N_19804,N_19979);
nor U20336 (N_20336,N_19974,N_19888);
nor U20337 (N_20337,N_19858,N_20086);
nand U20338 (N_20338,N_20041,N_19821);
nand U20339 (N_20339,N_20047,N_19947);
and U20340 (N_20340,N_20037,N_20021);
or U20341 (N_20341,N_20097,N_19963);
nor U20342 (N_20342,N_20048,N_19971);
xor U20343 (N_20343,N_19944,N_20004);
or U20344 (N_20344,N_20006,N_19946);
xor U20345 (N_20345,N_19909,N_19817);
xnor U20346 (N_20346,N_19851,N_19926);
nand U20347 (N_20347,N_19887,N_19800);
nor U20348 (N_20348,N_19873,N_19831);
xnor U20349 (N_20349,N_20039,N_20056);
xnor U20350 (N_20350,N_20009,N_19946);
nor U20351 (N_20351,N_20011,N_19988);
nand U20352 (N_20352,N_19964,N_20094);
or U20353 (N_20353,N_20065,N_19817);
xor U20354 (N_20354,N_19973,N_19880);
nor U20355 (N_20355,N_19817,N_19805);
nor U20356 (N_20356,N_19811,N_19818);
nor U20357 (N_20357,N_19959,N_20026);
nor U20358 (N_20358,N_19884,N_20019);
nand U20359 (N_20359,N_19978,N_20097);
or U20360 (N_20360,N_19898,N_19843);
xor U20361 (N_20361,N_20033,N_19853);
or U20362 (N_20362,N_19966,N_20003);
xnor U20363 (N_20363,N_19969,N_19812);
and U20364 (N_20364,N_20029,N_19862);
or U20365 (N_20365,N_20040,N_19902);
nor U20366 (N_20366,N_19927,N_19830);
and U20367 (N_20367,N_19839,N_19934);
nor U20368 (N_20368,N_20022,N_20038);
nand U20369 (N_20369,N_19859,N_19831);
nor U20370 (N_20370,N_20050,N_19832);
xnor U20371 (N_20371,N_19982,N_19959);
and U20372 (N_20372,N_19943,N_20059);
and U20373 (N_20373,N_20024,N_20041);
nor U20374 (N_20374,N_20096,N_20035);
nand U20375 (N_20375,N_19998,N_19904);
or U20376 (N_20376,N_20046,N_19901);
and U20377 (N_20377,N_20036,N_19912);
or U20378 (N_20378,N_19930,N_19814);
or U20379 (N_20379,N_19814,N_20087);
xnor U20380 (N_20380,N_20019,N_19888);
xnor U20381 (N_20381,N_19905,N_19929);
or U20382 (N_20382,N_20087,N_19858);
nand U20383 (N_20383,N_20028,N_19860);
or U20384 (N_20384,N_19863,N_20016);
nor U20385 (N_20385,N_19929,N_19850);
nand U20386 (N_20386,N_19912,N_20049);
or U20387 (N_20387,N_20073,N_19920);
nor U20388 (N_20388,N_19944,N_19965);
nand U20389 (N_20389,N_19939,N_20071);
or U20390 (N_20390,N_19978,N_19957);
nand U20391 (N_20391,N_19847,N_20022);
nand U20392 (N_20392,N_19964,N_20014);
and U20393 (N_20393,N_20074,N_19941);
and U20394 (N_20394,N_19842,N_19899);
and U20395 (N_20395,N_19939,N_20024);
and U20396 (N_20396,N_20084,N_19962);
and U20397 (N_20397,N_19911,N_20044);
xor U20398 (N_20398,N_19977,N_19865);
nor U20399 (N_20399,N_19946,N_20075);
or U20400 (N_20400,N_20199,N_20367);
nor U20401 (N_20401,N_20390,N_20290);
nor U20402 (N_20402,N_20321,N_20197);
nand U20403 (N_20403,N_20135,N_20232);
xor U20404 (N_20404,N_20339,N_20107);
nor U20405 (N_20405,N_20381,N_20267);
xor U20406 (N_20406,N_20100,N_20266);
nand U20407 (N_20407,N_20349,N_20136);
and U20408 (N_20408,N_20388,N_20345);
nand U20409 (N_20409,N_20270,N_20129);
xor U20410 (N_20410,N_20278,N_20109);
or U20411 (N_20411,N_20366,N_20250);
xnor U20412 (N_20412,N_20298,N_20368);
and U20413 (N_20413,N_20263,N_20173);
nand U20414 (N_20414,N_20139,N_20149);
nor U20415 (N_20415,N_20247,N_20116);
nand U20416 (N_20416,N_20281,N_20359);
or U20417 (N_20417,N_20104,N_20279);
and U20418 (N_20418,N_20287,N_20258);
nand U20419 (N_20419,N_20260,N_20373);
and U20420 (N_20420,N_20108,N_20393);
nor U20421 (N_20421,N_20257,N_20162);
xor U20422 (N_20422,N_20307,N_20334);
nand U20423 (N_20423,N_20350,N_20315);
and U20424 (N_20424,N_20276,N_20175);
nand U20425 (N_20425,N_20120,N_20328);
or U20426 (N_20426,N_20291,N_20330);
and U20427 (N_20427,N_20374,N_20244);
xor U20428 (N_20428,N_20202,N_20382);
and U20429 (N_20429,N_20377,N_20383);
xor U20430 (N_20430,N_20180,N_20274);
nor U20431 (N_20431,N_20118,N_20165);
and U20432 (N_20432,N_20344,N_20255);
xnor U20433 (N_20433,N_20295,N_20396);
nor U20434 (N_20434,N_20204,N_20213);
nor U20435 (N_20435,N_20229,N_20314);
nand U20436 (N_20436,N_20124,N_20191);
nor U20437 (N_20437,N_20141,N_20220);
nand U20438 (N_20438,N_20233,N_20317);
nor U20439 (N_20439,N_20121,N_20379);
or U20440 (N_20440,N_20284,N_20293);
nor U20441 (N_20441,N_20361,N_20269);
nand U20442 (N_20442,N_20215,N_20217);
or U20443 (N_20443,N_20308,N_20370);
nand U20444 (N_20444,N_20203,N_20194);
nor U20445 (N_20445,N_20126,N_20256);
xnor U20446 (N_20446,N_20206,N_20117);
xor U20447 (N_20447,N_20369,N_20254);
nand U20448 (N_20448,N_20322,N_20309);
or U20449 (N_20449,N_20398,N_20242);
nand U20450 (N_20450,N_20211,N_20351);
xor U20451 (N_20451,N_20186,N_20190);
nand U20452 (N_20452,N_20205,N_20272);
nor U20453 (N_20453,N_20376,N_20185);
nand U20454 (N_20454,N_20259,N_20277);
nor U20455 (N_20455,N_20133,N_20386);
xor U20456 (N_20456,N_20354,N_20358);
nor U20457 (N_20457,N_20112,N_20360);
or U20458 (N_20458,N_20159,N_20184);
and U20459 (N_20459,N_20389,N_20289);
nand U20460 (N_20460,N_20297,N_20312);
or U20461 (N_20461,N_20391,N_20148);
or U20462 (N_20462,N_20245,N_20127);
or U20463 (N_20463,N_20337,N_20222);
or U20464 (N_20464,N_20316,N_20146);
nor U20465 (N_20465,N_20218,N_20364);
xnor U20466 (N_20466,N_20169,N_20239);
nor U20467 (N_20467,N_20236,N_20384);
nor U20468 (N_20468,N_20111,N_20134);
nor U20469 (N_20469,N_20347,N_20122);
nand U20470 (N_20470,N_20235,N_20323);
xor U20471 (N_20471,N_20338,N_20302);
or U20472 (N_20472,N_20170,N_20219);
nor U20473 (N_20473,N_20147,N_20157);
and U20474 (N_20474,N_20193,N_20226);
nand U20475 (N_20475,N_20332,N_20340);
nor U20476 (N_20476,N_20299,N_20301);
and U20477 (N_20477,N_20251,N_20252);
nand U20478 (N_20478,N_20224,N_20282);
or U20479 (N_20479,N_20192,N_20319);
xor U20480 (N_20480,N_20200,N_20285);
xor U20481 (N_20481,N_20234,N_20326);
xor U20482 (N_20482,N_20150,N_20201);
nand U20483 (N_20483,N_20140,N_20336);
nor U20484 (N_20484,N_20207,N_20198);
and U20485 (N_20485,N_20105,N_20187);
nor U20486 (N_20486,N_20294,N_20331);
and U20487 (N_20487,N_20357,N_20221);
nand U20488 (N_20488,N_20188,N_20305);
or U20489 (N_20489,N_20113,N_20304);
xor U20490 (N_20490,N_20372,N_20375);
nor U20491 (N_20491,N_20362,N_20228);
nor U20492 (N_20492,N_20310,N_20399);
and U20493 (N_20493,N_20155,N_20195);
nand U20494 (N_20494,N_20378,N_20125);
or U20495 (N_20495,N_20154,N_20318);
nor U20496 (N_20496,N_20166,N_20152);
xor U20497 (N_20497,N_20253,N_20397);
or U20498 (N_20498,N_20246,N_20212);
or U20499 (N_20499,N_20237,N_20356);
or U20500 (N_20500,N_20286,N_20352);
or U20501 (N_20501,N_20320,N_20335);
nor U20502 (N_20502,N_20160,N_20161);
xor U20503 (N_20503,N_20261,N_20128);
nor U20504 (N_20504,N_20313,N_20132);
or U20505 (N_20505,N_20167,N_20292);
nor U20506 (N_20506,N_20248,N_20262);
xor U20507 (N_20507,N_20210,N_20385);
or U20508 (N_20508,N_20392,N_20230);
nand U20509 (N_20509,N_20115,N_20243);
and U20510 (N_20510,N_20353,N_20264);
xnor U20511 (N_20511,N_20280,N_20138);
and U20512 (N_20512,N_20182,N_20153);
nand U20513 (N_20513,N_20249,N_20174);
nor U20514 (N_20514,N_20324,N_20231);
or U20515 (N_20515,N_20311,N_20164);
nand U20516 (N_20516,N_20380,N_20333);
nor U20517 (N_20517,N_20342,N_20225);
or U20518 (N_20518,N_20343,N_20163);
nor U20519 (N_20519,N_20142,N_20131);
xor U20520 (N_20520,N_20238,N_20348);
xor U20521 (N_20521,N_20179,N_20355);
and U20522 (N_20522,N_20296,N_20143);
or U20523 (N_20523,N_20273,N_20327);
nand U20524 (N_20524,N_20275,N_20106);
or U20525 (N_20525,N_20325,N_20181);
nand U20526 (N_20526,N_20208,N_20110);
nor U20527 (N_20527,N_20271,N_20183);
and U20528 (N_20528,N_20177,N_20172);
and U20529 (N_20529,N_20394,N_20114);
nor U20530 (N_20530,N_20395,N_20123);
and U20531 (N_20531,N_20214,N_20103);
nand U20532 (N_20532,N_20300,N_20341);
and U20533 (N_20533,N_20283,N_20137);
and U20534 (N_20534,N_20176,N_20130);
and U20535 (N_20535,N_20156,N_20241);
xor U20536 (N_20536,N_20365,N_20329);
xnor U20537 (N_20537,N_20119,N_20371);
and U20538 (N_20538,N_20346,N_20145);
nor U20539 (N_20539,N_20303,N_20288);
nand U20540 (N_20540,N_20144,N_20102);
and U20541 (N_20541,N_20168,N_20363);
nor U20542 (N_20542,N_20223,N_20265);
or U20543 (N_20543,N_20151,N_20158);
nor U20544 (N_20544,N_20171,N_20268);
nor U20545 (N_20545,N_20189,N_20387);
nand U20546 (N_20546,N_20178,N_20306);
nand U20547 (N_20547,N_20216,N_20227);
xor U20548 (N_20548,N_20209,N_20196);
xnor U20549 (N_20549,N_20240,N_20101);
xnor U20550 (N_20550,N_20273,N_20261);
nor U20551 (N_20551,N_20160,N_20173);
nand U20552 (N_20552,N_20142,N_20285);
nor U20553 (N_20553,N_20179,N_20351);
nand U20554 (N_20554,N_20159,N_20183);
xor U20555 (N_20555,N_20260,N_20104);
or U20556 (N_20556,N_20349,N_20217);
nand U20557 (N_20557,N_20125,N_20188);
and U20558 (N_20558,N_20185,N_20177);
xnor U20559 (N_20559,N_20152,N_20189);
or U20560 (N_20560,N_20217,N_20371);
xor U20561 (N_20561,N_20199,N_20276);
and U20562 (N_20562,N_20397,N_20219);
and U20563 (N_20563,N_20142,N_20243);
and U20564 (N_20564,N_20186,N_20333);
nand U20565 (N_20565,N_20312,N_20332);
nand U20566 (N_20566,N_20230,N_20126);
nand U20567 (N_20567,N_20280,N_20316);
nand U20568 (N_20568,N_20315,N_20129);
nand U20569 (N_20569,N_20303,N_20245);
nor U20570 (N_20570,N_20177,N_20268);
nor U20571 (N_20571,N_20141,N_20361);
xnor U20572 (N_20572,N_20300,N_20165);
xor U20573 (N_20573,N_20319,N_20285);
xnor U20574 (N_20574,N_20105,N_20169);
xnor U20575 (N_20575,N_20328,N_20129);
or U20576 (N_20576,N_20391,N_20184);
nor U20577 (N_20577,N_20344,N_20228);
nor U20578 (N_20578,N_20269,N_20335);
nand U20579 (N_20579,N_20263,N_20131);
and U20580 (N_20580,N_20189,N_20160);
and U20581 (N_20581,N_20274,N_20362);
nor U20582 (N_20582,N_20111,N_20242);
nand U20583 (N_20583,N_20122,N_20100);
nand U20584 (N_20584,N_20347,N_20307);
xor U20585 (N_20585,N_20285,N_20292);
and U20586 (N_20586,N_20396,N_20388);
xnor U20587 (N_20587,N_20349,N_20142);
and U20588 (N_20588,N_20256,N_20146);
or U20589 (N_20589,N_20390,N_20133);
xnor U20590 (N_20590,N_20265,N_20221);
nand U20591 (N_20591,N_20267,N_20176);
and U20592 (N_20592,N_20346,N_20152);
nor U20593 (N_20593,N_20323,N_20302);
nor U20594 (N_20594,N_20150,N_20283);
nand U20595 (N_20595,N_20224,N_20351);
and U20596 (N_20596,N_20308,N_20174);
nor U20597 (N_20597,N_20253,N_20155);
xnor U20598 (N_20598,N_20162,N_20121);
nand U20599 (N_20599,N_20390,N_20181);
or U20600 (N_20600,N_20156,N_20312);
nor U20601 (N_20601,N_20209,N_20219);
or U20602 (N_20602,N_20301,N_20254);
nor U20603 (N_20603,N_20362,N_20233);
nor U20604 (N_20604,N_20228,N_20198);
and U20605 (N_20605,N_20204,N_20226);
nand U20606 (N_20606,N_20398,N_20300);
nor U20607 (N_20607,N_20184,N_20293);
nand U20608 (N_20608,N_20254,N_20326);
or U20609 (N_20609,N_20213,N_20356);
or U20610 (N_20610,N_20181,N_20287);
nor U20611 (N_20611,N_20221,N_20237);
nor U20612 (N_20612,N_20304,N_20205);
xnor U20613 (N_20613,N_20327,N_20290);
nand U20614 (N_20614,N_20384,N_20130);
and U20615 (N_20615,N_20378,N_20344);
nand U20616 (N_20616,N_20263,N_20396);
nor U20617 (N_20617,N_20139,N_20302);
nor U20618 (N_20618,N_20217,N_20297);
xnor U20619 (N_20619,N_20190,N_20270);
and U20620 (N_20620,N_20193,N_20331);
xor U20621 (N_20621,N_20239,N_20238);
nor U20622 (N_20622,N_20392,N_20158);
nor U20623 (N_20623,N_20148,N_20250);
and U20624 (N_20624,N_20111,N_20372);
nand U20625 (N_20625,N_20337,N_20216);
nand U20626 (N_20626,N_20354,N_20173);
or U20627 (N_20627,N_20254,N_20232);
or U20628 (N_20628,N_20194,N_20201);
or U20629 (N_20629,N_20279,N_20183);
or U20630 (N_20630,N_20331,N_20322);
and U20631 (N_20631,N_20369,N_20290);
nor U20632 (N_20632,N_20118,N_20125);
and U20633 (N_20633,N_20371,N_20171);
nand U20634 (N_20634,N_20134,N_20312);
xor U20635 (N_20635,N_20318,N_20217);
or U20636 (N_20636,N_20368,N_20247);
xor U20637 (N_20637,N_20316,N_20296);
or U20638 (N_20638,N_20352,N_20353);
and U20639 (N_20639,N_20300,N_20330);
nand U20640 (N_20640,N_20377,N_20300);
or U20641 (N_20641,N_20162,N_20198);
and U20642 (N_20642,N_20214,N_20152);
nor U20643 (N_20643,N_20107,N_20170);
and U20644 (N_20644,N_20376,N_20171);
nand U20645 (N_20645,N_20160,N_20310);
or U20646 (N_20646,N_20249,N_20382);
and U20647 (N_20647,N_20115,N_20252);
nand U20648 (N_20648,N_20243,N_20289);
and U20649 (N_20649,N_20100,N_20220);
nand U20650 (N_20650,N_20244,N_20108);
nand U20651 (N_20651,N_20165,N_20124);
and U20652 (N_20652,N_20110,N_20383);
nor U20653 (N_20653,N_20390,N_20326);
nor U20654 (N_20654,N_20265,N_20301);
or U20655 (N_20655,N_20153,N_20206);
nand U20656 (N_20656,N_20251,N_20382);
xnor U20657 (N_20657,N_20169,N_20390);
nor U20658 (N_20658,N_20133,N_20306);
nor U20659 (N_20659,N_20289,N_20378);
nor U20660 (N_20660,N_20104,N_20258);
or U20661 (N_20661,N_20282,N_20251);
or U20662 (N_20662,N_20193,N_20162);
xor U20663 (N_20663,N_20151,N_20170);
or U20664 (N_20664,N_20321,N_20314);
or U20665 (N_20665,N_20296,N_20347);
and U20666 (N_20666,N_20234,N_20132);
nor U20667 (N_20667,N_20303,N_20277);
or U20668 (N_20668,N_20279,N_20318);
and U20669 (N_20669,N_20110,N_20216);
and U20670 (N_20670,N_20358,N_20120);
xor U20671 (N_20671,N_20208,N_20162);
or U20672 (N_20672,N_20166,N_20355);
nand U20673 (N_20673,N_20126,N_20109);
nand U20674 (N_20674,N_20213,N_20191);
and U20675 (N_20675,N_20370,N_20246);
and U20676 (N_20676,N_20111,N_20257);
and U20677 (N_20677,N_20278,N_20220);
xnor U20678 (N_20678,N_20307,N_20351);
xnor U20679 (N_20679,N_20119,N_20169);
and U20680 (N_20680,N_20231,N_20167);
xor U20681 (N_20681,N_20221,N_20184);
nand U20682 (N_20682,N_20299,N_20382);
nand U20683 (N_20683,N_20106,N_20223);
xnor U20684 (N_20684,N_20154,N_20118);
nand U20685 (N_20685,N_20239,N_20377);
and U20686 (N_20686,N_20386,N_20148);
or U20687 (N_20687,N_20133,N_20299);
or U20688 (N_20688,N_20323,N_20110);
or U20689 (N_20689,N_20315,N_20359);
or U20690 (N_20690,N_20120,N_20339);
nor U20691 (N_20691,N_20230,N_20294);
nor U20692 (N_20692,N_20291,N_20233);
nor U20693 (N_20693,N_20236,N_20347);
nand U20694 (N_20694,N_20261,N_20156);
nand U20695 (N_20695,N_20294,N_20368);
or U20696 (N_20696,N_20287,N_20351);
and U20697 (N_20697,N_20282,N_20365);
xnor U20698 (N_20698,N_20329,N_20105);
or U20699 (N_20699,N_20182,N_20224);
xor U20700 (N_20700,N_20583,N_20677);
or U20701 (N_20701,N_20531,N_20629);
nor U20702 (N_20702,N_20664,N_20460);
nand U20703 (N_20703,N_20517,N_20630);
nand U20704 (N_20704,N_20421,N_20426);
nand U20705 (N_20705,N_20642,N_20661);
nor U20706 (N_20706,N_20621,N_20488);
nand U20707 (N_20707,N_20672,N_20604);
nand U20708 (N_20708,N_20509,N_20667);
nand U20709 (N_20709,N_20571,N_20680);
or U20710 (N_20710,N_20491,N_20690);
or U20711 (N_20711,N_20648,N_20434);
or U20712 (N_20712,N_20575,N_20572);
nor U20713 (N_20713,N_20401,N_20579);
xor U20714 (N_20714,N_20526,N_20599);
nand U20715 (N_20715,N_20437,N_20469);
xnor U20716 (N_20716,N_20576,N_20515);
xor U20717 (N_20717,N_20492,N_20405);
xnor U20718 (N_20718,N_20414,N_20639);
nor U20719 (N_20719,N_20637,N_20649);
nor U20720 (N_20720,N_20679,N_20423);
and U20721 (N_20721,N_20499,N_20456);
or U20722 (N_20722,N_20502,N_20494);
nand U20723 (N_20723,N_20624,N_20605);
xnor U20724 (N_20724,N_20673,N_20597);
or U20725 (N_20725,N_20564,N_20487);
nand U20726 (N_20726,N_20429,N_20668);
nand U20727 (N_20727,N_20558,N_20631);
xor U20728 (N_20728,N_20441,N_20546);
nor U20729 (N_20729,N_20520,N_20645);
nand U20730 (N_20730,N_20547,N_20403);
nand U20731 (N_20731,N_20446,N_20692);
xnor U20732 (N_20732,N_20602,N_20620);
xnor U20733 (N_20733,N_20540,N_20698);
and U20734 (N_20734,N_20651,N_20475);
and U20735 (N_20735,N_20543,N_20574);
or U20736 (N_20736,N_20689,N_20566);
nand U20737 (N_20737,N_20686,N_20694);
nand U20738 (N_20738,N_20550,N_20527);
or U20739 (N_20739,N_20697,N_20560);
nor U20740 (N_20740,N_20640,N_20551);
or U20741 (N_20741,N_20623,N_20532);
nand U20742 (N_20742,N_20568,N_20472);
and U20743 (N_20743,N_20402,N_20610);
or U20744 (N_20744,N_20500,N_20592);
or U20745 (N_20745,N_20582,N_20656);
xnor U20746 (N_20746,N_20508,N_20495);
nand U20747 (N_20747,N_20635,N_20577);
nand U20748 (N_20748,N_20471,N_20409);
and U20749 (N_20749,N_20559,N_20554);
nor U20750 (N_20750,N_20479,N_20544);
nor U20751 (N_20751,N_20596,N_20449);
and U20752 (N_20752,N_20643,N_20563);
and U20753 (N_20753,N_20504,N_20617);
nand U20754 (N_20754,N_20658,N_20622);
xor U20755 (N_20755,N_20524,N_20486);
or U20756 (N_20756,N_20525,N_20632);
nand U20757 (N_20757,N_20611,N_20650);
xnor U20758 (N_20758,N_20534,N_20691);
and U20759 (N_20759,N_20497,N_20557);
and U20760 (N_20760,N_20687,N_20444);
and U20761 (N_20761,N_20452,N_20608);
nor U20762 (N_20762,N_20465,N_20625);
and U20763 (N_20763,N_20587,N_20607);
nor U20764 (N_20764,N_20482,N_20549);
or U20765 (N_20765,N_20514,N_20603);
nand U20766 (N_20766,N_20493,N_20503);
xnor U20767 (N_20767,N_20545,N_20669);
xor U20768 (N_20768,N_20512,N_20541);
nand U20769 (N_20769,N_20448,N_20432);
xor U20770 (N_20770,N_20454,N_20478);
and U20771 (N_20771,N_20489,N_20627);
nor U20772 (N_20772,N_20485,N_20407);
nand U20773 (N_20773,N_20511,N_20655);
and U20774 (N_20774,N_20609,N_20428);
nand U20775 (N_20775,N_20606,N_20612);
or U20776 (N_20776,N_20552,N_20430);
xnor U20777 (N_20777,N_20408,N_20418);
or U20778 (N_20778,N_20591,N_20496);
nand U20779 (N_20779,N_20684,N_20436);
and U20780 (N_20780,N_20628,N_20425);
nor U20781 (N_20781,N_20580,N_20590);
or U20782 (N_20782,N_20675,N_20638);
xor U20783 (N_20783,N_20589,N_20647);
nand U20784 (N_20784,N_20585,N_20513);
nand U20785 (N_20785,N_20450,N_20439);
or U20786 (N_20786,N_20681,N_20420);
and U20787 (N_20787,N_20613,N_20594);
nor U20788 (N_20788,N_20537,N_20474);
and U20789 (N_20789,N_20404,N_20548);
nand U20790 (N_20790,N_20696,N_20674);
nand U20791 (N_20791,N_20556,N_20483);
or U20792 (N_20792,N_20490,N_20455);
nand U20793 (N_20793,N_20411,N_20614);
or U20794 (N_20794,N_20431,N_20433);
or U20795 (N_20795,N_20657,N_20601);
nor U20796 (N_20796,N_20435,N_20676);
or U20797 (N_20797,N_20522,N_20542);
nor U20798 (N_20798,N_20466,N_20535);
and U20799 (N_20799,N_20633,N_20641);
or U20800 (N_20800,N_20682,N_20652);
nor U20801 (N_20801,N_20473,N_20442);
or U20802 (N_20802,N_20467,N_20453);
nand U20803 (N_20803,N_20413,N_20653);
and U20804 (N_20804,N_20615,N_20663);
nor U20805 (N_20805,N_20626,N_20518);
nand U20806 (N_20806,N_20459,N_20484);
xor U20807 (N_20807,N_20406,N_20538);
and U20808 (N_20808,N_20506,N_20695);
and U20809 (N_20809,N_20480,N_20419);
or U20810 (N_20810,N_20427,N_20581);
nand U20811 (N_20811,N_20660,N_20555);
or U20812 (N_20812,N_20561,N_20659);
and U20813 (N_20813,N_20445,N_20440);
or U20814 (N_20814,N_20510,N_20519);
and U20815 (N_20815,N_20464,N_20468);
and U20816 (N_20816,N_20415,N_20646);
or U20817 (N_20817,N_20619,N_20678);
nor U20818 (N_20818,N_20400,N_20593);
or U20819 (N_20819,N_20654,N_20586);
or U20820 (N_20820,N_20463,N_20670);
nand U20821 (N_20821,N_20616,N_20477);
xor U20822 (N_20822,N_20443,N_20507);
xor U20823 (N_20823,N_20476,N_20461);
nor U20824 (N_20824,N_20417,N_20412);
or U20825 (N_20825,N_20644,N_20634);
nand U20826 (N_20826,N_20588,N_20470);
and U20827 (N_20827,N_20595,N_20451);
or U20828 (N_20828,N_20521,N_20666);
or U20829 (N_20829,N_20462,N_20458);
and U20830 (N_20830,N_20533,N_20501);
nor U20831 (N_20831,N_20523,N_20578);
or U20832 (N_20832,N_20438,N_20565);
or U20833 (N_20833,N_20573,N_20584);
or U20834 (N_20834,N_20618,N_20665);
or U20835 (N_20835,N_20570,N_20598);
and U20836 (N_20836,N_20685,N_20567);
nand U20837 (N_20837,N_20671,N_20422);
or U20838 (N_20838,N_20530,N_20424);
and U20839 (N_20839,N_20539,N_20481);
xor U20840 (N_20840,N_20699,N_20536);
nand U20841 (N_20841,N_20662,N_20683);
nor U20842 (N_20842,N_20410,N_20688);
nand U20843 (N_20843,N_20693,N_20447);
and U20844 (N_20844,N_20529,N_20569);
nor U20845 (N_20845,N_20505,N_20553);
xor U20846 (N_20846,N_20528,N_20457);
or U20847 (N_20847,N_20516,N_20416);
xnor U20848 (N_20848,N_20636,N_20562);
nand U20849 (N_20849,N_20600,N_20498);
or U20850 (N_20850,N_20554,N_20468);
xnor U20851 (N_20851,N_20595,N_20577);
nand U20852 (N_20852,N_20679,N_20416);
nor U20853 (N_20853,N_20448,N_20546);
nor U20854 (N_20854,N_20568,N_20517);
nor U20855 (N_20855,N_20405,N_20668);
xor U20856 (N_20856,N_20489,N_20541);
nor U20857 (N_20857,N_20531,N_20411);
or U20858 (N_20858,N_20433,N_20488);
nor U20859 (N_20859,N_20510,N_20593);
or U20860 (N_20860,N_20443,N_20621);
or U20861 (N_20861,N_20445,N_20601);
xnor U20862 (N_20862,N_20557,N_20464);
nand U20863 (N_20863,N_20631,N_20668);
or U20864 (N_20864,N_20663,N_20623);
xor U20865 (N_20865,N_20670,N_20513);
or U20866 (N_20866,N_20622,N_20470);
nor U20867 (N_20867,N_20513,N_20652);
xnor U20868 (N_20868,N_20484,N_20590);
nand U20869 (N_20869,N_20598,N_20440);
or U20870 (N_20870,N_20429,N_20422);
xnor U20871 (N_20871,N_20427,N_20402);
xnor U20872 (N_20872,N_20654,N_20425);
nor U20873 (N_20873,N_20584,N_20660);
or U20874 (N_20874,N_20413,N_20484);
nor U20875 (N_20875,N_20515,N_20567);
or U20876 (N_20876,N_20437,N_20450);
nor U20877 (N_20877,N_20433,N_20541);
nand U20878 (N_20878,N_20696,N_20625);
nand U20879 (N_20879,N_20606,N_20572);
nor U20880 (N_20880,N_20586,N_20578);
xnor U20881 (N_20881,N_20642,N_20684);
xnor U20882 (N_20882,N_20499,N_20418);
nor U20883 (N_20883,N_20502,N_20684);
and U20884 (N_20884,N_20451,N_20498);
nor U20885 (N_20885,N_20561,N_20607);
nor U20886 (N_20886,N_20683,N_20505);
nand U20887 (N_20887,N_20680,N_20562);
and U20888 (N_20888,N_20627,N_20595);
and U20889 (N_20889,N_20678,N_20443);
and U20890 (N_20890,N_20539,N_20681);
nor U20891 (N_20891,N_20490,N_20535);
nand U20892 (N_20892,N_20476,N_20459);
nor U20893 (N_20893,N_20671,N_20442);
and U20894 (N_20894,N_20501,N_20476);
nand U20895 (N_20895,N_20633,N_20504);
and U20896 (N_20896,N_20488,N_20455);
nor U20897 (N_20897,N_20472,N_20660);
nor U20898 (N_20898,N_20660,N_20622);
or U20899 (N_20899,N_20617,N_20669);
and U20900 (N_20900,N_20586,N_20621);
nand U20901 (N_20901,N_20499,N_20689);
nor U20902 (N_20902,N_20495,N_20451);
nand U20903 (N_20903,N_20643,N_20609);
or U20904 (N_20904,N_20567,N_20536);
xnor U20905 (N_20905,N_20698,N_20530);
xnor U20906 (N_20906,N_20455,N_20476);
nor U20907 (N_20907,N_20689,N_20495);
nand U20908 (N_20908,N_20546,N_20404);
or U20909 (N_20909,N_20423,N_20412);
or U20910 (N_20910,N_20696,N_20560);
nand U20911 (N_20911,N_20628,N_20485);
xor U20912 (N_20912,N_20646,N_20638);
nand U20913 (N_20913,N_20528,N_20598);
nor U20914 (N_20914,N_20469,N_20605);
xnor U20915 (N_20915,N_20659,N_20680);
or U20916 (N_20916,N_20547,N_20695);
and U20917 (N_20917,N_20591,N_20472);
and U20918 (N_20918,N_20623,N_20631);
nand U20919 (N_20919,N_20404,N_20593);
or U20920 (N_20920,N_20420,N_20643);
and U20921 (N_20921,N_20533,N_20437);
xnor U20922 (N_20922,N_20501,N_20523);
or U20923 (N_20923,N_20587,N_20565);
xor U20924 (N_20924,N_20411,N_20555);
nor U20925 (N_20925,N_20556,N_20462);
nand U20926 (N_20926,N_20539,N_20422);
xor U20927 (N_20927,N_20584,N_20575);
nor U20928 (N_20928,N_20405,N_20414);
nand U20929 (N_20929,N_20403,N_20427);
or U20930 (N_20930,N_20561,N_20605);
xor U20931 (N_20931,N_20539,N_20678);
xnor U20932 (N_20932,N_20541,N_20416);
or U20933 (N_20933,N_20498,N_20596);
or U20934 (N_20934,N_20505,N_20524);
xor U20935 (N_20935,N_20588,N_20481);
and U20936 (N_20936,N_20621,N_20490);
and U20937 (N_20937,N_20479,N_20699);
nand U20938 (N_20938,N_20447,N_20420);
nand U20939 (N_20939,N_20419,N_20481);
xor U20940 (N_20940,N_20562,N_20575);
xor U20941 (N_20941,N_20639,N_20604);
or U20942 (N_20942,N_20666,N_20465);
nor U20943 (N_20943,N_20535,N_20480);
and U20944 (N_20944,N_20477,N_20494);
or U20945 (N_20945,N_20534,N_20593);
and U20946 (N_20946,N_20539,N_20661);
or U20947 (N_20947,N_20533,N_20643);
or U20948 (N_20948,N_20425,N_20499);
xnor U20949 (N_20949,N_20641,N_20510);
and U20950 (N_20950,N_20674,N_20550);
nand U20951 (N_20951,N_20636,N_20478);
xor U20952 (N_20952,N_20550,N_20587);
nor U20953 (N_20953,N_20688,N_20462);
and U20954 (N_20954,N_20430,N_20588);
and U20955 (N_20955,N_20408,N_20629);
or U20956 (N_20956,N_20682,N_20657);
nand U20957 (N_20957,N_20678,N_20518);
and U20958 (N_20958,N_20547,N_20422);
nand U20959 (N_20959,N_20615,N_20629);
and U20960 (N_20960,N_20628,N_20533);
or U20961 (N_20961,N_20422,N_20458);
xor U20962 (N_20962,N_20472,N_20406);
and U20963 (N_20963,N_20417,N_20618);
nor U20964 (N_20964,N_20649,N_20669);
and U20965 (N_20965,N_20665,N_20590);
or U20966 (N_20966,N_20587,N_20645);
and U20967 (N_20967,N_20512,N_20613);
and U20968 (N_20968,N_20548,N_20443);
nor U20969 (N_20969,N_20496,N_20521);
nand U20970 (N_20970,N_20647,N_20566);
and U20971 (N_20971,N_20648,N_20432);
xnor U20972 (N_20972,N_20581,N_20672);
xor U20973 (N_20973,N_20447,N_20619);
nand U20974 (N_20974,N_20465,N_20406);
or U20975 (N_20975,N_20402,N_20602);
nor U20976 (N_20976,N_20508,N_20666);
xnor U20977 (N_20977,N_20522,N_20659);
and U20978 (N_20978,N_20641,N_20485);
and U20979 (N_20979,N_20637,N_20472);
and U20980 (N_20980,N_20630,N_20655);
nand U20981 (N_20981,N_20669,N_20600);
and U20982 (N_20982,N_20650,N_20413);
xor U20983 (N_20983,N_20499,N_20597);
nor U20984 (N_20984,N_20569,N_20626);
or U20985 (N_20985,N_20691,N_20649);
or U20986 (N_20986,N_20460,N_20440);
or U20987 (N_20987,N_20559,N_20639);
nand U20988 (N_20988,N_20520,N_20684);
xor U20989 (N_20989,N_20497,N_20699);
xor U20990 (N_20990,N_20680,N_20514);
nor U20991 (N_20991,N_20436,N_20580);
or U20992 (N_20992,N_20690,N_20590);
nand U20993 (N_20993,N_20494,N_20647);
nor U20994 (N_20994,N_20509,N_20671);
nand U20995 (N_20995,N_20437,N_20504);
nor U20996 (N_20996,N_20575,N_20552);
and U20997 (N_20997,N_20684,N_20540);
nand U20998 (N_20998,N_20652,N_20574);
xor U20999 (N_20999,N_20493,N_20430);
xnor U21000 (N_21000,N_20880,N_20723);
nor U21001 (N_21001,N_20737,N_20722);
xnor U21002 (N_21002,N_20735,N_20901);
or U21003 (N_21003,N_20760,N_20958);
xor U21004 (N_21004,N_20970,N_20995);
and U21005 (N_21005,N_20892,N_20973);
or U21006 (N_21006,N_20949,N_20736);
nor U21007 (N_21007,N_20822,N_20785);
nand U21008 (N_21008,N_20777,N_20869);
and U21009 (N_21009,N_20919,N_20748);
or U21010 (N_21010,N_20939,N_20766);
and U21011 (N_21011,N_20845,N_20897);
nor U21012 (N_21012,N_20727,N_20799);
xnor U21013 (N_21013,N_20806,N_20975);
xnor U21014 (N_21014,N_20969,N_20961);
nand U21015 (N_21015,N_20933,N_20831);
nand U21016 (N_21016,N_20718,N_20786);
and U21017 (N_21017,N_20936,N_20950);
nor U21018 (N_21018,N_20765,N_20772);
or U21019 (N_21019,N_20996,N_20798);
nand U21020 (N_21020,N_20745,N_20860);
nor U21021 (N_21021,N_20854,N_20768);
nand U21022 (N_21022,N_20853,N_20856);
and U21023 (N_21023,N_20848,N_20773);
and U21024 (N_21024,N_20792,N_20755);
nor U21025 (N_21025,N_20729,N_20866);
and U21026 (N_21026,N_20867,N_20837);
xnor U21027 (N_21027,N_20721,N_20931);
or U21028 (N_21028,N_20841,N_20927);
xor U21029 (N_21029,N_20994,N_20796);
nand U21030 (N_21030,N_20700,N_20835);
or U21031 (N_21031,N_20808,N_20740);
nand U21032 (N_21032,N_20731,N_20879);
nand U21033 (N_21033,N_20813,N_20871);
nand U21034 (N_21034,N_20944,N_20708);
nor U21035 (N_21035,N_20907,N_20793);
and U21036 (N_21036,N_20713,N_20971);
xnor U21037 (N_21037,N_20929,N_20870);
xnor U21038 (N_21038,N_20703,N_20844);
and U21039 (N_21039,N_20938,N_20830);
or U21040 (N_21040,N_20937,N_20990);
nand U21041 (N_21041,N_20895,N_20805);
or U21042 (N_21042,N_20902,N_20899);
nor U21043 (N_21043,N_20797,N_20982);
nand U21044 (N_21044,N_20855,N_20826);
xor U21045 (N_21045,N_20967,N_20877);
xnor U21046 (N_21046,N_20992,N_20839);
xor U21047 (N_21047,N_20894,N_20840);
or U21048 (N_21048,N_20753,N_20842);
nand U21049 (N_21049,N_20734,N_20743);
and U21050 (N_21050,N_20955,N_20758);
or U21051 (N_21051,N_20847,N_20861);
xor U21052 (N_21052,N_20781,N_20999);
and U21053 (N_21053,N_20751,N_20956);
xnor U21054 (N_21054,N_20925,N_20882);
xnor U21055 (N_21055,N_20818,N_20834);
or U21056 (N_21056,N_20732,N_20749);
nor U21057 (N_21057,N_20779,N_20791);
xor U21058 (N_21058,N_20711,N_20885);
nor U21059 (N_21059,N_20770,N_20863);
nand U21060 (N_21060,N_20774,N_20801);
or U21061 (N_21061,N_20888,N_20966);
nand U21062 (N_21062,N_20828,N_20803);
and U21063 (N_21063,N_20780,N_20893);
nand U21064 (N_21064,N_20954,N_20726);
and U21065 (N_21065,N_20878,N_20787);
nor U21066 (N_21066,N_20701,N_20904);
nor U21067 (N_21067,N_20756,N_20940);
xnor U21068 (N_21068,N_20912,N_20788);
and U21069 (N_21069,N_20807,N_20814);
or U21070 (N_21070,N_20945,N_20960);
xor U21071 (N_21071,N_20811,N_20782);
and U21072 (N_21072,N_20794,N_20942);
or U21073 (N_21073,N_20857,N_20948);
or U21074 (N_21074,N_20819,N_20875);
xor U21075 (N_21075,N_20754,N_20930);
nor U21076 (N_21076,N_20859,N_20916);
and U21077 (N_21077,N_20928,N_20923);
and U21078 (N_21078,N_20771,N_20884);
and U21079 (N_21079,N_20997,N_20874);
nor U21080 (N_21080,N_20915,N_20769);
or U21081 (N_21081,N_20891,N_20724);
and U21082 (N_21082,N_20763,N_20715);
or U21083 (N_21083,N_20712,N_20889);
or U21084 (N_21084,N_20795,N_20738);
or U21085 (N_21085,N_20963,N_20728);
nand U21086 (N_21086,N_20984,N_20921);
or U21087 (N_21087,N_20838,N_20914);
or U21088 (N_21088,N_20935,N_20725);
or U21089 (N_21089,N_20951,N_20824);
nor U21090 (N_21090,N_20881,N_20742);
nor U21091 (N_21091,N_20993,N_20825);
nor U21092 (N_21092,N_20896,N_20908);
and U21093 (N_21093,N_20974,N_20716);
nand U21094 (N_21094,N_20764,N_20707);
xor U21095 (N_21095,N_20709,N_20823);
nand U21096 (N_21096,N_20900,N_20783);
and U21097 (N_21097,N_20829,N_20775);
and U21098 (N_21098,N_20981,N_20762);
nand U21099 (N_21099,N_20827,N_20833);
nand U21100 (N_21100,N_20964,N_20947);
xnor U21101 (N_21101,N_20864,N_20858);
xnor U21102 (N_21102,N_20702,N_20800);
nor U21103 (N_21103,N_20789,N_20920);
xor U21104 (N_21104,N_20849,N_20776);
nand U21105 (N_21105,N_20741,N_20832);
or U21106 (N_21106,N_20922,N_20810);
and U21107 (N_21107,N_20876,N_20816);
or U21108 (N_21108,N_20821,N_20784);
nand U21109 (N_21109,N_20976,N_20978);
nand U21110 (N_21110,N_20890,N_20977);
and U21111 (N_21111,N_20790,N_20979);
xor U21112 (N_21112,N_20988,N_20809);
nor U21113 (N_21113,N_20968,N_20862);
or U21114 (N_21114,N_20932,N_20957);
nor U21115 (N_21115,N_20759,N_20905);
nand U21116 (N_21116,N_20744,N_20903);
or U21117 (N_21117,N_20991,N_20911);
xnor U21118 (N_21118,N_20972,N_20917);
or U21119 (N_21119,N_20733,N_20998);
or U21120 (N_21120,N_20924,N_20815);
nor U21121 (N_21121,N_20714,N_20962);
and U21122 (N_21122,N_20872,N_20719);
nor U21123 (N_21123,N_20986,N_20868);
nand U21124 (N_21124,N_20865,N_20965);
nor U21125 (N_21125,N_20750,N_20752);
and U21126 (N_21126,N_20757,N_20873);
xnor U21127 (N_21127,N_20778,N_20706);
nor U21128 (N_21128,N_20705,N_20934);
or U21129 (N_21129,N_20851,N_20906);
and U21130 (N_21130,N_20953,N_20717);
nor U21131 (N_21131,N_20761,N_20817);
and U21132 (N_21132,N_20846,N_20812);
nor U21133 (N_21133,N_20980,N_20730);
nor U21134 (N_21134,N_20913,N_20989);
xor U21135 (N_21135,N_20710,N_20898);
and U21136 (N_21136,N_20820,N_20910);
nor U21137 (N_21137,N_20941,N_20704);
xor U21138 (N_21138,N_20952,N_20746);
nor U21139 (N_21139,N_20804,N_20767);
and U21140 (N_21140,N_20720,N_20836);
and U21141 (N_21141,N_20946,N_20985);
and U21142 (N_21142,N_20959,N_20850);
nor U21143 (N_21143,N_20852,N_20747);
nand U21144 (N_21144,N_20926,N_20943);
and U21145 (N_21145,N_20843,N_20739);
or U21146 (N_21146,N_20983,N_20886);
nand U21147 (N_21147,N_20802,N_20987);
nor U21148 (N_21148,N_20918,N_20909);
nor U21149 (N_21149,N_20887,N_20883);
xor U21150 (N_21150,N_20970,N_20739);
and U21151 (N_21151,N_20843,N_20738);
or U21152 (N_21152,N_20878,N_20987);
nor U21153 (N_21153,N_20728,N_20778);
nor U21154 (N_21154,N_20823,N_20955);
nor U21155 (N_21155,N_20876,N_20728);
nand U21156 (N_21156,N_20956,N_20994);
xor U21157 (N_21157,N_20943,N_20732);
nand U21158 (N_21158,N_20712,N_20745);
nand U21159 (N_21159,N_20912,N_20828);
or U21160 (N_21160,N_20778,N_20813);
xor U21161 (N_21161,N_20918,N_20813);
and U21162 (N_21162,N_20742,N_20826);
xnor U21163 (N_21163,N_20751,N_20960);
or U21164 (N_21164,N_20995,N_20962);
nand U21165 (N_21165,N_20959,N_20739);
nand U21166 (N_21166,N_20707,N_20756);
nor U21167 (N_21167,N_20841,N_20771);
nand U21168 (N_21168,N_20858,N_20959);
and U21169 (N_21169,N_20839,N_20786);
and U21170 (N_21170,N_20729,N_20768);
nor U21171 (N_21171,N_20758,N_20887);
and U21172 (N_21172,N_20956,N_20879);
nor U21173 (N_21173,N_20903,N_20723);
and U21174 (N_21174,N_20898,N_20800);
nor U21175 (N_21175,N_20777,N_20804);
nand U21176 (N_21176,N_20773,N_20999);
nand U21177 (N_21177,N_20829,N_20863);
or U21178 (N_21178,N_20994,N_20995);
and U21179 (N_21179,N_20821,N_20712);
nand U21180 (N_21180,N_20799,N_20786);
nand U21181 (N_21181,N_20898,N_20982);
and U21182 (N_21182,N_20979,N_20903);
nand U21183 (N_21183,N_20963,N_20775);
and U21184 (N_21184,N_20776,N_20768);
nand U21185 (N_21185,N_20810,N_20740);
nor U21186 (N_21186,N_20731,N_20843);
xnor U21187 (N_21187,N_20795,N_20993);
and U21188 (N_21188,N_20876,N_20729);
and U21189 (N_21189,N_20941,N_20953);
and U21190 (N_21190,N_20946,N_20730);
xor U21191 (N_21191,N_20707,N_20742);
and U21192 (N_21192,N_20940,N_20913);
nor U21193 (N_21193,N_20885,N_20975);
nand U21194 (N_21194,N_20981,N_20772);
nor U21195 (N_21195,N_20979,N_20977);
or U21196 (N_21196,N_20969,N_20723);
and U21197 (N_21197,N_20997,N_20856);
xor U21198 (N_21198,N_20844,N_20706);
nor U21199 (N_21199,N_20957,N_20949);
or U21200 (N_21200,N_20941,N_20823);
xnor U21201 (N_21201,N_20929,N_20722);
xor U21202 (N_21202,N_20925,N_20888);
nand U21203 (N_21203,N_20898,N_20914);
nor U21204 (N_21204,N_20702,N_20801);
nor U21205 (N_21205,N_20976,N_20948);
nand U21206 (N_21206,N_20936,N_20776);
and U21207 (N_21207,N_20715,N_20805);
xnor U21208 (N_21208,N_20865,N_20913);
and U21209 (N_21209,N_20761,N_20777);
nor U21210 (N_21210,N_20978,N_20746);
xnor U21211 (N_21211,N_20728,N_20770);
nand U21212 (N_21212,N_20976,N_20944);
and U21213 (N_21213,N_20769,N_20970);
or U21214 (N_21214,N_20934,N_20909);
and U21215 (N_21215,N_20720,N_20730);
nand U21216 (N_21216,N_20932,N_20823);
xor U21217 (N_21217,N_20731,N_20859);
nand U21218 (N_21218,N_20737,N_20839);
nor U21219 (N_21219,N_20841,N_20863);
nor U21220 (N_21220,N_20882,N_20918);
nor U21221 (N_21221,N_20730,N_20790);
or U21222 (N_21222,N_20723,N_20784);
nand U21223 (N_21223,N_20900,N_20709);
and U21224 (N_21224,N_20797,N_20814);
nand U21225 (N_21225,N_20957,N_20802);
nor U21226 (N_21226,N_20965,N_20702);
xnor U21227 (N_21227,N_20858,N_20925);
or U21228 (N_21228,N_20776,N_20707);
or U21229 (N_21229,N_20734,N_20922);
or U21230 (N_21230,N_20956,N_20882);
nor U21231 (N_21231,N_20903,N_20946);
nand U21232 (N_21232,N_20835,N_20860);
xnor U21233 (N_21233,N_20937,N_20914);
xnor U21234 (N_21234,N_20745,N_20847);
nand U21235 (N_21235,N_20773,N_20916);
or U21236 (N_21236,N_20776,N_20860);
nand U21237 (N_21237,N_20953,N_20826);
nor U21238 (N_21238,N_20957,N_20831);
nor U21239 (N_21239,N_20907,N_20778);
or U21240 (N_21240,N_20771,N_20986);
or U21241 (N_21241,N_20770,N_20832);
nor U21242 (N_21242,N_20770,N_20786);
nor U21243 (N_21243,N_20998,N_20927);
xor U21244 (N_21244,N_20717,N_20805);
nand U21245 (N_21245,N_20761,N_20779);
and U21246 (N_21246,N_20877,N_20992);
and U21247 (N_21247,N_20819,N_20983);
or U21248 (N_21248,N_20848,N_20828);
nor U21249 (N_21249,N_20716,N_20966);
and U21250 (N_21250,N_20771,N_20995);
xnor U21251 (N_21251,N_20964,N_20886);
nand U21252 (N_21252,N_20783,N_20949);
xor U21253 (N_21253,N_20784,N_20858);
nand U21254 (N_21254,N_20788,N_20702);
or U21255 (N_21255,N_20840,N_20891);
nor U21256 (N_21256,N_20977,N_20842);
nor U21257 (N_21257,N_20947,N_20879);
xnor U21258 (N_21258,N_20889,N_20705);
xor U21259 (N_21259,N_20736,N_20821);
xor U21260 (N_21260,N_20903,N_20948);
or U21261 (N_21261,N_20891,N_20877);
and U21262 (N_21262,N_20820,N_20815);
nor U21263 (N_21263,N_20831,N_20914);
nor U21264 (N_21264,N_20765,N_20867);
and U21265 (N_21265,N_20887,N_20991);
and U21266 (N_21266,N_20847,N_20771);
nor U21267 (N_21267,N_20977,N_20983);
xor U21268 (N_21268,N_20907,N_20784);
and U21269 (N_21269,N_20715,N_20884);
xor U21270 (N_21270,N_20797,N_20944);
and U21271 (N_21271,N_20709,N_20977);
xnor U21272 (N_21272,N_20767,N_20706);
or U21273 (N_21273,N_20862,N_20754);
or U21274 (N_21274,N_20762,N_20816);
xnor U21275 (N_21275,N_20725,N_20783);
and U21276 (N_21276,N_20855,N_20934);
nor U21277 (N_21277,N_20813,N_20950);
or U21278 (N_21278,N_20913,N_20841);
nand U21279 (N_21279,N_20843,N_20895);
and U21280 (N_21280,N_20934,N_20775);
or U21281 (N_21281,N_20982,N_20855);
and U21282 (N_21282,N_20894,N_20949);
nand U21283 (N_21283,N_20980,N_20945);
xor U21284 (N_21284,N_20877,N_20901);
nor U21285 (N_21285,N_20989,N_20761);
and U21286 (N_21286,N_20887,N_20750);
nor U21287 (N_21287,N_20931,N_20835);
nand U21288 (N_21288,N_20753,N_20866);
and U21289 (N_21289,N_20736,N_20706);
nor U21290 (N_21290,N_20830,N_20950);
xnor U21291 (N_21291,N_20871,N_20793);
or U21292 (N_21292,N_20935,N_20710);
nand U21293 (N_21293,N_20883,N_20748);
or U21294 (N_21294,N_20834,N_20832);
xor U21295 (N_21295,N_20832,N_20850);
xnor U21296 (N_21296,N_20856,N_20826);
nor U21297 (N_21297,N_20893,N_20830);
xnor U21298 (N_21298,N_20897,N_20797);
or U21299 (N_21299,N_20885,N_20821);
or U21300 (N_21300,N_21259,N_21253);
or U21301 (N_21301,N_21150,N_21138);
or U21302 (N_21302,N_21108,N_21143);
or U21303 (N_21303,N_21289,N_21225);
and U21304 (N_21304,N_21173,N_21181);
xnor U21305 (N_21305,N_21104,N_21023);
nor U21306 (N_21306,N_21055,N_21217);
or U21307 (N_21307,N_21050,N_21117);
and U21308 (N_21308,N_21171,N_21273);
and U21309 (N_21309,N_21030,N_21132);
nor U21310 (N_21310,N_21135,N_21003);
nand U21311 (N_21311,N_21202,N_21060);
or U21312 (N_21312,N_21158,N_21082);
or U21313 (N_21313,N_21099,N_21236);
or U21314 (N_21314,N_21064,N_21001);
xnor U21315 (N_21315,N_21269,N_21007);
or U21316 (N_21316,N_21260,N_21053);
or U21317 (N_21317,N_21027,N_21167);
and U21318 (N_21318,N_21109,N_21151);
and U21319 (N_21319,N_21268,N_21112);
xor U21320 (N_21320,N_21279,N_21069);
nand U21321 (N_21321,N_21278,N_21272);
or U21322 (N_21322,N_21221,N_21215);
and U21323 (N_21323,N_21013,N_21256);
and U21324 (N_21324,N_21098,N_21157);
or U21325 (N_21325,N_21034,N_21041);
xor U21326 (N_21326,N_21194,N_21015);
or U21327 (N_21327,N_21258,N_21089);
and U21328 (N_21328,N_21292,N_21242);
or U21329 (N_21329,N_21287,N_21125);
xor U21330 (N_21330,N_21185,N_21039);
and U21331 (N_21331,N_21239,N_21049);
nand U21332 (N_21332,N_21092,N_21263);
nand U21333 (N_21333,N_21214,N_21080);
or U21334 (N_21334,N_21190,N_21175);
and U21335 (N_21335,N_21119,N_21193);
xnor U21336 (N_21336,N_21164,N_21065);
or U21337 (N_21337,N_21101,N_21228);
or U21338 (N_21338,N_21182,N_21254);
or U21339 (N_21339,N_21203,N_21271);
nand U21340 (N_21340,N_21057,N_21029);
or U21341 (N_21341,N_21006,N_21229);
xor U21342 (N_21342,N_21111,N_21103);
xor U21343 (N_21343,N_21226,N_21154);
nor U21344 (N_21344,N_21037,N_21234);
or U21345 (N_21345,N_21142,N_21018);
nor U21346 (N_21346,N_21275,N_21146);
and U21347 (N_21347,N_21004,N_21093);
nor U21348 (N_21348,N_21245,N_21068);
xor U21349 (N_21349,N_21038,N_21116);
or U21350 (N_21350,N_21212,N_21172);
and U21351 (N_21351,N_21120,N_21243);
and U21352 (N_21352,N_21128,N_21261);
and U21353 (N_21353,N_21075,N_21085);
xnor U21354 (N_21354,N_21113,N_21024);
nand U21355 (N_21355,N_21042,N_21189);
nor U21356 (N_21356,N_21016,N_21071);
and U21357 (N_21357,N_21141,N_21086);
xnor U21358 (N_21358,N_21067,N_21293);
xor U21359 (N_21359,N_21094,N_21235);
nand U21360 (N_21360,N_21073,N_21056);
nand U21361 (N_21361,N_21161,N_21047);
nand U21362 (N_21362,N_21147,N_21148);
and U21363 (N_21363,N_21081,N_21061);
or U21364 (N_21364,N_21045,N_21284);
nand U21365 (N_21365,N_21074,N_21066);
nand U21366 (N_21366,N_21097,N_21137);
nor U21367 (N_21367,N_21241,N_21031);
and U21368 (N_21368,N_21083,N_21149);
nand U21369 (N_21369,N_21233,N_21298);
xnor U21370 (N_21370,N_21012,N_21277);
or U21371 (N_21371,N_21224,N_21204);
xor U21372 (N_21372,N_21105,N_21195);
xor U21373 (N_21373,N_21043,N_21266);
and U21374 (N_21374,N_21163,N_21197);
or U21375 (N_21375,N_21044,N_21062);
and U21376 (N_21376,N_21000,N_21145);
and U21377 (N_21377,N_21286,N_21162);
or U21378 (N_21378,N_21170,N_21238);
nor U21379 (N_21379,N_21177,N_21188);
xnor U21380 (N_21380,N_21210,N_21107);
nor U21381 (N_21381,N_21264,N_21255);
xnor U21382 (N_21382,N_21178,N_21186);
nor U21383 (N_21383,N_21088,N_21250);
or U21384 (N_21384,N_21048,N_21131);
nand U21385 (N_21385,N_21223,N_21052);
and U21386 (N_21386,N_21035,N_21232);
xnor U21387 (N_21387,N_21121,N_21096);
nor U21388 (N_21388,N_21025,N_21114);
or U21389 (N_21389,N_21072,N_21191);
or U21390 (N_21390,N_21288,N_21248);
nand U21391 (N_21391,N_21297,N_21021);
nand U21392 (N_21392,N_21227,N_21276);
or U21393 (N_21393,N_21285,N_21136);
nand U21394 (N_21394,N_21265,N_21249);
and U21395 (N_21395,N_21002,N_21010);
nor U21396 (N_21396,N_21222,N_21009);
nand U21397 (N_21397,N_21160,N_21208);
nor U21398 (N_21398,N_21198,N_21123);
nand U21399 (N_21399,N_21270,N_21246);
nor U21400 (N_21400,N_21176,N_21078);
xor U21401 (N_21401,N_21218,N_21155);
nand U21402 (N_21402,N_21187,N_21299);
and U21403 (N_21403,N_21011,N_21032);
and U21404 (N_21404,N_21207,N_21124);
and U21405 (N_21405,N_21140,N_21058);
xor U21406 (N_21406,N_21231,N_21054);
and U21407 (N_21407,N_21192,N_21184);
or U21408 (N_21408,N_21087,N_21059);
or U21409 (N_21409,N_21153,N_21280);
and U21410 (N_21410,N_21174,N_21063);
and U21411 (N_21411,N_21206,N_21166);
and U21412 (N_21412,N_21100,N_21283);
or U21413 (N_21413,N_21017,N_21077);
nand U21414 (N_21414,N_21091,N_21126);
nor U21415 (N_21415,N_21110,N_21106);
xor U21416 (N_21416,N_21040,N_21014);
nand U21417 (N_21417,N_21183,N_21294);
or U21418 (N_21418,N_21196,N_21144);
nand U21419 (N_21419,N_21282,N_21095);
or U21420 (N_21420,N_21251,N_21130);
nor U21421 (N_21421,N_21156,N_21022);
nand U21422 (N_21422,N_21252,N_21033);
or U21423 (N_21423,N_21169,N_21118);
nand U21424 (N_21424,N_21046,N_21291);
or U21425 (N_21425,N_21084,N_21019);
nor U21426 (N_21426,N_21201,N_21051);
nand U21427 (N_21427,N_21165,N_21281);
or U21428 (N_21428,N_21219,N_21216);
nand U21429 (N_21429,N_21295,N_21020);
or U21430 (N_21430,N_21026,N_21267);
nand U21431 (N_21431,N_21274,N_21079);
or U21432 (N_21432,N_21076,N_21129);
nor U21433 (N_21433,N_21247,N_21028);
nor U21434 (N_21434,N_21290,N_21159);
and U21435 (N_21435,N_21090,N_21127);
and U21436 (N_21436,N_21070,N_21296);
or U21437 (N_21437,N_21005,N_21102);
nor U21438 (N_21438,N_21257,N_21139);
and U21439 (N_21439,N_21008,N_21180);
nand U21440 (N_21440,N_21213,N_21115);
xnor U21441 (N_21441,N_21199,N_21262);
xnor U21442 (N_21442,N_21122,N_21237);
and U21443 (N_21443,N_21152,N_21133);
xor U21444 (N_21444,N_21220,N_21240);
nor U21445 (N_21445,N_21036,N_21230);
nor U21446 (N_21446,N_21211,N_21134);
xor U21447 (N_21447,N_21168,N_21244);
nand U21448 (N_21448,N_21200,N_21205);
nor U21449 (N_21449,N_21209,N_21179);
xnor U21450 (N_21450,N_21125,N_21116);
xnor U21451 (N_21451,N_21146,N_21087);
nand U21452 (N_21452,N_21154,N_21295);
nor U21453 (N_21453,N_21056,N_21219);
and U21454 (N_21454,N_21097,N_21098);
or U21455 (N_21455,N_21296,N_21291);
and U21456 (N_21456,N_21060,N_21138);
nor U21457 (N_21457,N_21060,N_21223);
or U21458 (N_21458,N_21205,N_21261);
nor U21459 (N_21459,N_21008,N_21003);
nand U21460 (N_21460,N_21040,N_21006);
and U21461 (N_21461,N_21026,N_21180);
nand U21462 (N_21462,N_21295,N_21091);
and U21463 (N_21463,N_21289,N_21187);
nand U21464 (N_21464,N_21266,N_21268);
nor U21465 (N_21465,N_21012,N_21100);
xnor U21466 (N_21466,N_21148,N_21234);
nor U21467 (N_21467,N_21110,N_21071);
or U21468 (N_21468,N_21261,N_21167);
nand U21469 (N_21469,N_21202,N_21046);
xor U21470 (N_21470,N_21166,N_21215);
xnor U21471 (N_21471,N_21160,N_21174);
nor U21472 (N_21472,N_21236,N_21234);
nor U21473 (N_21473,N_21110,N_21231);
or U21474 (N_21474,N_21197,N_21100);
nand U21475 (N_21475,N_21108,N_21169);
and U21476 (N_21476,N_21215,N_21290);
nor U21477 (N_21477,N_21069,N_21274);
xnor U21478 (N_21478,N_21100,N_21015);
xnor U21479 (N_21479,N_21208,N_21192);
nand U21480 (N_21480,N_21214,N_21207);
xnor U21481 (N_21481,N_21130,N_21026);
or U21482 (N_21482,N_21224,N_21280);
or U21483 (N_21483,N_21018,N_21190);
or U21484 (N_21484,N_21036,N_21283);
xor U21485 (N_21485,N_21025,N_21112);
or U21486 (N_21486,N_21287,N_21079);
nor U21487 (N_21487,N_21182,N_21114);
and U21488 (N_21488,N_21064,N_21006);
or U21489 (N_21489,N_21127,N_21145);
nor U21490 (N_21490,N_21173,N_21085);
and U21491 (N_21491,N_21052,N_21054);
xnor U21492 (N_21492,N_21250,N_21241);
and U21493 (N_21493,N_21127,N_21141);
xnor U21494 (N_21494,N_21140,N_21157);
xor U21495 (N_21495,N_21195,N_21140);
and U21496 (N_21496,N_21111,N_21247);
nor U21497 (N_21497,N_21057,N_21181);
nand U21498 (N_21498,N_21243,N_21202);
or U21499 (N_21499,N_21011,N_21104);
and U21500 (N_21500,N_21002,N_21210);
and U21501 (N_21501,N_21214,N_21070);
or U21502 (N_21502,N_21210,N_21101);
and U21503 (N_21503,N_21079,N_21039);
nor U21504 (N_21504,N_21063,N_21214);
and U21505 (N_21505,N_21004,N_21263);
or U21506 (N_21506,N_21091,N_21259);
nand U21507 (N_21507,N_21137,N_21132);
nor U21508 (N_21508,N_21089,N_21096);
or U21509 (N_21509,N_21152,N_21058);
xor U21510 (N_21510,N_21288,N_21011);
xnor U21511 (N_21511,N_21099,N_21220);
and U21512 (N_21512,N_21294,N_21253);
or U21513 (N_21513,N_21085,N_21257);
xor U21514 (N_21514,N_21034,N_21217);
xnor U21515 (N_21515,N_21287,N_21242);
xor U21516 (N_21516,N_21241,N_21052);
nand U21517 (N_21517,N_21026,N_21232);
nand U21518 (N_21518,N_21075,N_21254);
or U21519 (N_21519,N_21102,N_21123);
nor U21520 (N_21520,N_21087,N_21247);
and U21521 (N_21521,N_21287,N_21272);
and U21522 (N_21522,N_21167,N_21045);
or U21523 (N_21523,N_21254,N_21063);
xnor U21524 (N_21524,N_21218,N_21179);
nand U21525 (N_21525,N_21086,N_21273);
or U21526 (N_21526,N_21118,N_21275);
and U21527 (N_21527,N_21255,N_21100);
or U21528 (N_21528,N_21226,N_21007);
xnor U21529 (N_21529,N_21120,N_21169);
and U21530 (N_21530,N_21217,N_21160);
xor U21531 (N_21531,N_21004,N_21102);
xnor U21532 (N_21532,N_21117,N_21208);
nand U21533 (N_21533,N_21106,N_21242);
or U21534 (N_21534,N_21276,N_21074);
and U21535 (N_21535,N_21290,N_21282);
and U21536 (N_21536,N_21103,N_21265);
and U21537 (N_21537,N_21282,N_21006);
or U21538 (N_21538,N_21123,N_21015);
nand U21539 (N_21539,N_21106,N_21082);
nor U21540 (N_21540,N_21013,N_21135);
and U21541 (N_21541,N_21128,N_21214);
and U21542 (N_21542,N_21169,N_21274);
and U21543 (N_21543,N_21153,N_21129);
xnor U21544 (N_21544,N_21061,N_21027);
and U21545 (N_21545,N_21293,N_21093);
xor U21546 (N_21546,N_21136,N_21270);
or U21547 (N_21547,N_21096,N_21102);
nand U21548 (N_21548,N_21288,N_21066);
nand U21549 (N_21549,N_21069,N_21033);
or U21550 (N_21550,N_21265,N_21256);
xor U21551 (N_21551,N_21295,N_21299);
or U21552 (N_21552,N_21224,N_21053);
nand U21553 (N_21553,N_21260,N_21023);
nor U21554 (N_21554,N_21148,N_21206);
and U21555 (N_21555,N_21274,N_21115);
and U21556 (N_21556,N_21055,N_21250);
nand U21557 (N_21557,N_21030,N_21216);
nor U21558 (N_21558,N_21264,N_21085);
nor U21559 (N_21559,N_21215,N_21188);
and U21560 (N_21560,N_21043,N_21177);
xor U21561 (N_21561,N_21210,N_21276);
or U21562 (N_21562,N_21057,N_21280);
and U21563 (N_21563,N_21273,N_21265);
xnor U21564 (N_21564,N_21149,N_21036);
or U21565 (N_21565,N_21015,N_21198);
or U21566 (N_21566,N_21086,N_21032);
or U21567 (N_21567,N_21008,N_21221);
nor U21568 (N_21568,N_21208,N_21011);
nor U21569 (N_21569,N_21295,N_21049);
and U21570 (N_21570,N_21157,N_21160);
or U21571 (N_21571,N_21158,N_21019);
xor U21572 (N_21572,N_21119,N_21029);
xor U21573 (N_21573,N_21027,N_21248);
xnor U21574 (N_21574,N_21093,N_21059);
xnor U21575 (N_21575,N_21180,N_21036);
nand U21576 (N_21576,N_21019,N_21176);
xnor U21577 (N_21577,N_21128,N_21203);
and U21578 (N_21578,N_21217,N_21246);
nor U21579 (N_21579,N_21001,N_21253);
nand U21580 (N_21580,N_21244,N_21037);
nand U21581 (N_21581,N_21225,N_21058);
or U21582 (N_21582,N_21070,N_21256);
nand U21583 (N_21583,N_21050,N_21063);
and U21584 (N_21584,N_21243,N_21225);
nor U21585 (N_21585,N_21072,N_21049);
nor U21586 (N_21586,N_21061,N_21133);
and U21587 (N_21587,N_21132,N_21260);
nor U21588 (N_21588,N_21158,N_21253);
or U21589 (N_21589,N_21036,N_21297);
nor U21590 (N_21590,N_21114,N_21278);
nand U21591 (N_21591,N_21149,N_21299);
nor U21592 (N_21592,N_21194,N_21025);
xnor U21593 (N_21593,N_21068,N_21203);
or U21594 (N_21594,N_21067,N_21237);
xnor U21595 (N_21595,N_21122,N_21073);
nand U21596 (N_21596,N_21230,N_21216);
nor U21597 (N_21597,N_21115,N_21175);
nand U21598 (N_21598,N_21162,N_21138);
nor U21599 (N_21599,N_21164,N_21223);
and U21600 (N_21600,N_21344,N_21397);
xnor U21601 (N_21601,N_21426,N_21553);
and U21602 (N_21602,N_21548,N_21468);
or U21603 (N_21603,N_21599,N_21534);
or U21604 (N_21604,N_21424,N_21489);
and U21605 (N_21605,N_21551,N_21362);
xnor U21606 (N_21606,N_21471,N_21358);
xor U21607 (N_21607,N_21510,N_21441);
xnor U21608 (N_21608,N_21374,N_21333);
or U21609 (N_21609,N_21419,N_21525);
xor U21610 (N_21610,N_21500,N_21403);
xor U21611 (N_21611,N_21336,N_21416);
and U21612 (N_21612,N_21519,N_21452);
and U21613 (N_21613,N_21316,N_21315);
nand U21614 (N_21614,N_21428,N_21400);
nand U21615 (N_21615,N_21559,N_21409);
or U21616 (N_21616,N_21460,N_21545);
and U21617 (N_21617,N_21487,N_21483);
xor U21618 (N_21618,N_21357,N_21550);
xor U21619 (N_21619,N_21557,N_21329);
nand U21620 (N_21620,N_21466,N_21528);
nand U21621 (N_21621,N_21579,N_21445);
xor U21622 (N_21622,N_21454,N_21375);
xnor U21623 (N_21623,N_21348,N_21367);
xor U21624 (N_21624,N_21393,N_21390);
nor U21625 (N_21625,N_21461,N_21539);
xnor U21626 (N_21626,N_21598,N_21398);
or U21627 (N_21627,N_21505,N_21427);
or U21628 (N_21628,N_21351,N_21328);
nor U21629 (N_21629,N_21469,N_21490);
nor U21630 (N_21630,N_21474,N_21577);
and U21631 (N_21631,N_21514,N_21517);
or U21632 (N_21632,N_21574,N_21492);
nand U21633 (N_21633,N_21325,N_21493);
or U21634 (N_21634,N_21417,N_21582);
xor U21635 (N_21635,N_21584,N_21502);
nor U21636 (N_21636,N_21418,N_21448);
and U21637 (N_21637,N_21556,N_21463);
or U21638 (N_21638,N_21479,N_21343);
xor U21639 (N_21639,N_21453,N_21413);
or U21640 (N_21640,N_21405,N_21485);
or U21641 (N_21641,N_21533,N_21438);
and U21642 (N_21642,N_21587,N_21597);
and U21643 (N_21643,N_21381,N_21341);
and U21644 (N_21644,N_21342,N_21371);
or U21645 (N_21645,N_21303,N_21547);
or U21646 (N_21646,N_21334,N_21580);
and U21647 (N_21647,N_21421,N_21472);
nor U21648 (N_21648,N_21563,N_21464);
nand U21649 (N_21649,N_21595,N_21572);
xor U21650 (N_21650,N_21338,N_21361);
and U21651 (N_21651,N_21522,N_21414);
xnor U21652 (N_21652,N_21449,N_21564);
and U21653 (N_21653,N_21432,N_21407);
xor U21654 (N_21654,N_21327,N_21354);
or U21655 (N_21655,N_21366,N_21364);
or U21656 (N_21656,N_21495,N_21345);
nor U21657 (N_21657,N_21571,N_21496);
xnor U21658 (N_21658,N_21331,N_21350);
nor U21659 (N_21659,N_21543,N_21433);
xor U21660 (N_21660,N_21570,N_21359);
and U21661 (N_21661,N_21549,N_21305);
nand U21662 (N_21662,N_21332,N_21423);
nor U21663 (N_21663,N_21594,N_21529);
and U21664 (N_21664,N_21446,N_21450);
nor U21665 (N_21665,N_21437,N_21566);
or U21666 (N_21666,N_21581,N_21434);
nor U21667 (N_21667,N_21411,N_21356);
and U21668 (N_21668,N_21395,N_21355);
nand U21669 (N_21669,N_21515,N_21526);
and U21670 (N_21670,N_21498,N_21470);
and U21671 (N_21671,N_21412,N_21318);
nand U21672 (N_21672,N_21484,N_21365);
nand U21673 (N_21673,N_21368,N_21513);
or U21674 (N_21674,N_21389,N_21337);
xnor U21675 (N_21675,N_21494,N_21444);
and U21676 (N_21676,N_21458,N_21586);
and U21677 (N_21677,N_21565,N_21527);
and U21678 (N_21678,N_21392,N_21473);
nand U21679 (N_21679,N_21309,N_21593);
nand U21680 (N_21680,N_21541,N_21535);
nor U21681 (N_21681,N_21406,N_21387);
nor U21682 (N_21682,N_21467,N_21532);
xor U21683 (N_21683,N_21503,N_21560);
xnor U21684 (N_21684,N_21482,N_21304);
nand U21685 (N_21685,N_21317,N_21537);
nand U21686 (N_21686,N_21455,N_21319);
xnor U21687 (N_21687,N_21352,N_21308);
xnor U21688 (N_21688,N_21552,N_21314);
nand U21689 (N_21689,N_21431,N_21567);
xor U21690 (N_21690,N_21504,N_21447);
nor U21691 (N_21691,N_21380,N_21562);
xor U21692 (N_21692,N_21462,N_21596);
and U21693 (N_21693,N_21386,N_21363);
nand U21694 (N_21694,N_21373,N_21512);
nand U21695 (N_21695,N_21307,N_21475);
xnor U21696 (N_21696,N_21330,N_21478);
or U21697 (N_21697,N_21507,N_21585);
nor U21698 (N_21698,N_21391,N_21353);
nor U21699 (N_21699,N_21360,N_21506);
nand U21700 (N_21700,N_21324,N_21524);
nand U21701 (N_21701,N_21326,N_21465);
or U21702 (N_21702,N_21476,N_21396);
xor U21703 (N_21703,N_21422,N_21301);
and U21704 (N_21704,N_21546,N_21516);
or U21705 (N_21705,N_21591,N_21456);
nand U21706 (N_21706,N_21491,N_21311);
nor U21707 (N_21707,N_21302,N_21477);
and U21708 (N_21708,N_21575,N_21404);
or U21709 (N_21709,N_21312,N_21521);
and U21710 (N_21710,N_21370,N_21382);
nor U21711 (N_21711,N_21538,N_21408);
or U21712 (N_21712,N_21530,N_21536);
or U21713 (N_21713,N_21349,N_21410);
or U21714 (N_21714,N_21402,N_21488);
xor U21715 (N_21715,N_21442,N_21531);
and U21716 (N_21716,N_21430,N_21440);
xnor U21717 (N_21717,N_21578,N_21583);
and U21718 (N_21718,N_21509,N_21429);
nand U21719 (N_21719,N_21511,N_21335);
or U21720 (N_21720,N_21415,N_21540);
and U21721 (N_21721,N_21520,N_21481);
nand U21722 (N_21722,N_21544,N_21590);
nor U21723 (N_21723,N_21320,N_21401);
nor U21724 (N_21724,N_21346,N_21569);
or U21725 (N_21725,N_21435,N_21378);
and U21726 (N_21726,N_21436,N_21480);
nor U21727 (N_21727,N_21300,N_21439);
and U21728 (N_21728,N_21347,N_21443);
xnor U21729 (N_21729,N_21523,N_21542);
or U21730 (N_21730,N_21518,N_21508);
and U21731 (N_21731,N_21555,N_21394);
nand U21732 (N_21732,N_21576,N_21340);
xor U21733 (N_21733,N_21589,N_21321);
nand U21734 (N_21734,N_21383,N_21323);
xnor U21735 (N_21735,N_21486,N_21499);
nand U21736 (N_21736,N_21377,N_21457);
nor U21737 (N_21737,N_21558,N_21592);
nor U21738 (N_21738,N_21376,N_21497);
nor U21739 (N_21739,N_21568,N_21369);
nor U21740 (N_21740,N_21384,N_21425);
nand U21741 (N_21741,N_21310,N_21372);
xor U21742 (N_21742,N_21306,N_21561);
nand U21743 (N_21743,N_21379,N_21339);
xor U21744 (N_21744,N_21588,N_21554);
nand U21745 (N_21745,N_21573,N_21388);
nor U21746 (N_21746,N_21451,N_21313);
and U21747 (N_21747,N_21385,N_21459);
xnor U21748 (N_21748,N_21501,N_21420);
or U21749 (N_21749,N_21399,N_21322);
and U21750 (N_21750,N_21331,N_21570);
and U21751 (N_21751,N_21319,N_21491);
nand U21752 (N_21752,N_21452,N_21432);
nor U21753 (N_21753,N_21429,N_21449);
or U21754 (N_21754,N_21459,N_21361);
or U21755 (N_21755,N_21476,N_21524);
nand U21756 (N_21756,N_21514,N_21442);
xnor U21757 (N_21757,N_21552,N_21426);
nand U21758 (N_21758,N_21447,N_21422);
nor U21759 (N_21759,N_21526,N_21439);
and U21760 (N_21760,N_21365,N_21427);
nand U21761 (N_21761,N_21563,N_21396);
and U21762 (N_21762,N_21509,N_21356);
nand U21763 (N_21763,N_21403,N_21493);
nor U21764 (N_21764,N_21497,N_21433);
nor U21765 (N_21765,N_21446,N_21432);
nor U21766 (N_21766,N_21360,N_21448);
and U21767 (N_21767,N_21490,N_21442);
or U21768 (N_21768,N_21391,N_21483);
xnor U21769 (N_21769,N_21551,N_21321);
nor U21770 (N_21770,N_21349,N_21333);
or U21771 (N_21771,N_21453,N_21479);
or U21772 (N_21772,N_21598,N_21556);
nor U21773 (N_21773,N_21523,N_21341);
and U21774 (N_21774,N_21346,N_21351);
or U21775 (N_21775,N_21449,N_21597);
xor U21776 (N_21776,N_21445,N_21403);
or U21777 (N_21777,N_21372,N_21547);
and U21778 (N_21778,N_21345,N_21474);
or U21779 (N_21779,N_21561,N_21578);
and U21780 (N_21780,N_21567,N_21570);
and U21781 (N_21781,N_21520,N_21460);
xnor U21782 (N_21782,N_21402,N_21496);
and U21783 (N_21783,N_21408,N_21477);
and U21784 (N_21784,N_21364,N_21517);
nor U21785 (N_21785,N_21305,N_21527);
xor U21786 (N_21786,N_21523,N_21350);
and U21787 (N_21787,N_21568,N_21566);
nand U21788 (N_21788,N_21546,N_21510);
nor U21789 (N_21789,N_21499,N_21419);
nor U21790 (N_21790,N_21579,N_21393);
nand U21791 (N_21791,N_21395,N_21575);
nor U21792 (N_21792,N_21449,N_21462);
xnor U21793 (N_21793,N_21418,N_21447);
nor U21794 (N_21794,N_21584,N_21583);
nor U21795 (N_21795,N_21515,N_21458);
or U21796 (N_21796,N_21526,N_21359);
nor U21797 (N_21797,N_21488,N_21520);
xor U21798 (N_21798,N_21584,N_21421);
nor U21799 (N_21799,N_21431,N_21515);
xnor U21800 (N_21800,N_21528,N_21316);
xor U21801 (N_21801,N_21405,N_21338);
nand U21802 (N_21802,N_21317,N_21329);
or U21803 (N_21803,N_21315,N_21597);
and U21804 (N_21804,N_21397,N_21550);
xnor U21805 (N_21805,N_21471,N_21598);
and U21806 (N_21806,N_21331,N_21357);
and U21807 (N_21807,N_21553,N_21435);
xnor U21808 (N_21808,N_21546,N_21509);
and U21809 (N_21809,N_21582,N_21432);
xnor U21810 (N_21810,N_21516,N_21436);
xor U21811 (N_21811,N_21557,N_21451);
xor U21812 (N_21812,N_21399,N_21503);
nor U21813 (N_21813,N_21503,N_21423);
and U21814 (N_21814,N_21348,N_21360);
nor U21815 (N_21815,N_21351,N_21411);
nor U21816 (N_21816,N_21453,N_21494);
nor U21817 (N_21817,N_21483,N_21437);
nor U21818 (N_21818,N_21321,N_21598);
nor U21819 (N_21819,N_21565,N_21305);
nor U21820 (N_21820,N_21349,N_21318);
and U21821 (N_21821,N_21500,N_21470);
and U21822 (N_21822,N_21416,N_21377);
xor U21823 (N_21823,N_21489,N_21467);
nor U21824 (N_21824,N_21549,N_21547);
and U21825 (N_21825,N_21461,N_21309);
or U21826 (N_21826,N_21419,N_21454);
nand U21827 (N_21827,N_21557,N_21545);
and U21828 (N_21828,N_21483,N_21516);
nor U21829 (N_21829,N_21538,N_21478);
nand U21830 (N_21830,N_21572,N_21370);
nand U21831 (N_21831,N_21374,N_21416);
or U21832 (N_21832,N_21330,N_21443);
or U21833 (N_21833,N_21346,N_21501);
xnor U21834 (N_21834,N_21351,N_21489);
xnor U21835 (N_21835,N_21407,N_21468);
nor U21836 (N_21836,N_21564,N_21553);
nand U21837 (N_21837,N_21525,N_21574);
and U21838 (N_21838,N_21507,N_21524);
xor U21839 (N_21839,N_21413,N_21528);
nand U21840 (N_21840,N_21479,N_21425);
nor U21841 (N_21841,N_21433,N_21435);
xor U21842 (N_21842,N_21445,N_21458);
or U21843 (N_21843,N_21455,N_21536);
or U21844 (N_21844,N_21499,N_21442);
nand U21845 (N_21845,N_21372,N_21433);
nand U21846 (N_21846,N_21320,N_21535);
or U21847 (N_21847,N_21531,N_21394);
nor U21848 (N_21848,N_21389,N_21535);
or U21849 (N_21849,N_21546,N_21305);
or U21850 (N_21850,N_21500,N_21368);
nand U21851 (N_21851,N_21535,N_21303);
and U21852 (N_21852,N_21517,N_21486);
and U21853 (N_21853,N_21498,N_21574);
xnor U21854 (N_21854,N_21384,N_21555);
xor U21855 (N_21855,N_21323,N_21523);
xnor U21856 (N_21856,N_21571,N_21539);
or U21857 (N_21857,N_21578,N_21437);
or U21858 (N_21858,N_21501,N_21535);
and U21859 (N_21859,N_21534,N_21584);
and U21860 (N_21860,N_21441,N_21308);
xor U21861 (N_21861,N_21590,N_21454);
xnor U21862 (N_21862,N_21401,N_21307);
xor U21863 (N_21863,N_21322,N_21402);
xnor U21864 (N_21864,N_21404,N_21424);
or U21865 (N_21865,N_21559,N_21525);
and U21866 (N_21866,N_21354,N_21441);
and U21867 (N_21867,N_21527,N_21583);
xor U21868 (N_21868,N_21571,N_21383);
nor U21869 (N_21869,N_21559,N_21400);
nand U21870 (N_21870,N_21343,N_21310);
nor U21871 (N_21871,N_21559,N_21315);
or U21872 (N_21872,N_21358,N_21443);
nor U21873 (N_21873,N_21387,N_21422);
nand U21874 (N_21874,N_21301,N_21394);
nand U21875 (N_21875,N_21533,N_21543);
xor U21876 (N_21876,N_21396,N_21406);
or U21877 (N_21877,N_21558,N_21330);
xnor U21878 (N_21878,N_21346,N_21467);
nor U21879 (N_21879,N_21339,N_21408);
and U21880 (N_21880,N_21562,N_21457);
or U21881 (N_21881,N_21468,N_21412);
xnor U21882 (N_21882,N_21408,N_21366);
and U21883 (N_21883,N_21421,N_21451);
xnor U21884 (N_21884,N_21571,N_21438);
xor U21885 (N_21885,N_21490,N_21437);
or U21886 (N_21886,N_21404,N_21316);
and U21887 (N_21887,N_21346,N_21446);
nor U21888 (N_21888,N_21579,N_21447);
and U21889 (N_21889,N_21307,N_21422);
or U21890 (N_21890,N_21330,N_21554);
and U21891 (N_21891,N_21503,N_21302);
or U21892 (N_21892,N_21576,N_21378);
xnor U21893 (N_21893,N_21594,N_21428);
xnor U21894 (N_21894,N_21474,N_21569);
and U21895 (N_21895,N_21571,N_21512);
and U21896 (N_21896,N_21594,N_21337);
nand U21897 (N_21897,N_21511,N_21440);
or U21898 (N_21898,N_21595,N_21555);
xnor U21899 (N_21899,N_21474,N_21407);
xor U21900 (N_21900,N_21653,N_21849);
xnor U21901 (N_21901,N_21714,N_21655);
nor U21902 (N_21902,N_21815,N_21847);
xor U21903 (N_21903,N_21797,N_21842);
or U21904 (N_21904,N_21687,N_21616);
xnor U21905 (N_21905,N_21892,N_21817);
and U21906 (N_21906,N_21767,N_21623);
nor U21907 (N_21907,N_21723,N_21646);
xnor U21908 (N_21908,N_21874,N_21780);
nand U21909 (N_21909,N_21765,N_21869);
or U21910 (N_21910,N_21666,N_21868);
and U21911 (N_21911,N_21864,N_21753);
nand U21912 (N_21912,N_21686,N_21730);
or U21913 (N_21913,N_21751,N_21820);
and U21914 (N_21914,N_21898,N_21705);
xnor U21915 (N_21915,N_21619,N_21720);
xnor U21916 (N_21916,N_21840,N_21731);
nor U21917 (N_21917,N_21673,N_21672);
or U21918 (N_21918,N_21813,N_21657);
or U21919 (N_21919,N_21664,N_21779);
nand U21920 (N_21920,N_21644,N_21876);
and U21921 (N_21921,N_21766,N_21871);
xor U21922 (N_21922,N_21677,N_21617);
nor U21923 (N_21923,N_21811,N_21659);
and U21924 (N_21924,N_21774,N_21703);
nand U21925 (N_21925,N_21776,N_21637);
or U21926 (N_21926,N_21689,N_21846);
xor U21927 (N_21927,N_21812,N_21852);
xnor U21928 (N_21928,N_21685,N_21837);
xnor U21929 (N_21929,N_21784,N_21785);
nand U21930 (N_21930,N_21782,N_21630);
and U21931 (N_21931,N_21738,N_21661);
nor U21932 (N_21932,N_21679,N_21880);
xor U21933 (N_21933,N_21665,N_21696);
or U21934 (N_21934,N_21702,N_21640);
or U21935 (N_21935,N_21609,N_21758);
nand U21936 (N_21936,N_21642,N_21608);
and U21937 (N_21937,N_21638,N_21899);
nor U21938 (N_21938,N_21744,N_21719);
xor U21939 (N_21939,N_21724,N_21693);
nor U21940 (N_21940,N_21746,N_21773);
xnor U21941 (N_21941,N_21841,N_21628);
and U21942 (N_21942,N_21794,N_21802);
nor U21943 (N_21943,N_21631,N_21682);
and U21944 (N_21944,N_21718,N_21825);
xnor U21945 (N_21945,N_21737,N_21881);
nor U21946 (N_21946,N_21770,N_21632);
xor U21947 (N_21947,N_21889,N_21828);
nand U21948 (N_21948,N_21771,N_21742);
xor U21949 (N_21949,N_21700,N_21688);
nor U21950 (N_21950,N_21824,N_21607);
nor U21951 (N_21951,N_21883,N_21829);
and U21952 (N_21952,N_21728,N_21887);
xor U21953 (N_21953,N_21821,N_21747);
and U21954 (N_21954,N_21756,N_21894);
xnor U21955 (N_21955,N_21676,N_21804);
nand U21956 (N_21956,N_21635,N_21645);
and U21957 (N_21957,N_21854,N_21740);
xnor U21958 (N_21958,N_21610,N_21778);
nor U21959 (N_21959,N_21614,N_21835);
xnor U21960 (N_21960,N_21736,N_21888);
nor U21961 (N_21961,N_21699,N_21851);
nand U21962 (N_21962,N_21755,N_21759);
or U21963 (N_21963,N_21656,N_21629);
or U21964 (N_21964,N_21896,N_21654);
nor U21965 (N_21965,N_21805,N_21791);
or U21966 (N_21966,N_21613,N_21684);
xor U21967 (N_21967,N_21890,N_21743);
nor U21968 (N_21968,N_21816,N_21711);
nor U21969 (N_21969,N_21612,N_21763);
xnor U21970 (N_21970,N_21856,N_21748);
nand U21971 (N_21971,N_21814,N_21600);
or U21972 (N_21972,N_21663,N_21741);
or U21973 (N_21973,N_21708,N_21877);
xnor U21974 (N_21974,N_21704,N_21691);
nor U21975 (N_21975,N_21826,N_21893);
or U21976 (N_21976,N_21798,N_21818);
xnor U21977 (N_21977,N_21707,N_21709);
nor U21978 (N_21978,N_21861,N_21866);
nand U21979 (N_21979,N_21606,N_21819);
and U21980 (N_21980,N_21618,N_21884);
or U21981 (N_21981,N_21683,N_21769);
or U21982 (N_21982,N_21808,N_21694);
and U21983 (N_21983,N_21641,N_21803);
and U21984 (N_21984,N_21757,N_21671);
nor U21985 (N_21985,N_21822,N_21649);
and U21986 (N_21986,N_21674,N_21611);
and U21987 (N_21987,N_21725,N_21845);
nand U21988 (N_21988,N_21648,N_21735);
and U21989 (N_21989,N_21697,N_21858);
and U21990 (N_21990,N_21839,N_21627);
and U21991 (N_21991,N_21809,N_21810);
xnor U21992 (N_21992,N_21831,N_21726);
and U21993 (N_21993,N_21860,N_21701);
nand U21994 (N_21994,N_21692,N_21639);
nor U21995 (N_21995,N_21651,N_21625);
or U21996 (N_21996,N_21729,N_21800);
nand U21997 (N_21997,N_21790,N_21850);
nand U21998 (N_21998,N_21667,N_21867);
nor U21999 (N_21999,N_21636,N_21716);
or U22000 (N_22000,N_21690,N_21650);
and U22001 (N_22001,N_21857,N_21749);
and U22002 (N_22002,N_21750,N_21643);
or U22003 (N_22003,N_21710,N_21615);
xor U22004 (N_22004,N_21732,N_21823);
xor U22005 (N_22005,N_21768,N_21873);
and U22006 (N_22006,N_21801,N_21603);
and U22007 (N_22007,N_21715,N_21886);
nand U22008 (N_22008,N_21764,N_21806);
nor U22009 (N_22009,N_21870,N_21662);
nor U22010 (N_22010,N_21652,N_21762);
xor U22011 (N_22011,N_21604,N_21891);
or U22012 (N_22012,N_21793,N_21620);
nor U22013 (N_22013,N_21775,N_21722);
xor U22014 (N_22014,N_21675,N_21777);
xor U22015 (N_22015,N_21853,N_21875);
or U22016 (N_22016,N_21678,N_21622);
nor U22017 (N_22017,N_21633,N_21660);
nor U22018 (N_22018,N_21783,N_21838);
or U22019 (N_22019,N_21786,N_21698);
xnor U22020 (N_22020,N_21799,N_21669);
or U22021 (N_22021,N_21795,N_21897);
nand U22022 (N_22022,N_21859,N_21772);
and U22023 (N_22023,N_21727,N_21787);
nor U22024 (N_22024,N_21827,N_21872);
and U22025 (N_22025,N_21807,N_21833);
nor U22026 (N_22026,N_21621,N_21878);
or U22027 (N_22027,N_21624,N_21602);
nor U22028 (N_22028,N_21668,N_21754);
or U22029 (N_22029,N_21734,N_21862);
or U22030 (N_22030,N_21760,N_21752);
nor U22031 (N_22031,N_21658,N_21739);
nor U22032 (N_22032,N_21796,N_21848);
nor U22033 (N_22033,N_21788,N_21680);
nor U22034 (N_22034,N_21733,N_21713);
or U22035 (N_22035,N_21843,N_21717);
and U22036 (N_22036,N_21706,N_21634);
or U22037 (N_22037,N_21792,N_21781);
nand U22038 (N_22038,N_21834,N_21681);
nor U22039 (N_22039,N_21695,N_21865);
and U22040 (N_22040,N_21712,N_21879);
nor U22041 (N_22041,N_21721,N_21647);
nand U22042 (N_22042,N_21626,N_21895);
xnor U22043 (N_22043,N_21830,N_21605);
or U22044 (N_22044,N_21855,N_21670);
nand U22045 (N_22045,N_21844,N_21601);
nand U22046 (N_22046,N_21863,N_21745);
or U22047 (N_22047,N_21832,N_21885);
and U22048 (N_22048,N_21882,N_21836);
or U22049 (N_22049,N_21789,N_21761);
or U22050 (N_22050,N_21778,N_21661);
nor U22051 (N_22051,N_21649,N_21723);
and U22052 (N_22052,N_21607,N_21841);
nand U22053 (N_22053,N_21680,N_21753);
nand U22054 (N_22054,N_21831,N_21770);
and U22055 (N_22055,N_21701,N_21833);
xor U22056 (N_22056,N_21617,N_21806);
nand U22057 (N_22057,N_21717,N_21603);
nor U22058 (N_22058,N_21890,N_21853);
nor U22059 (N_22059,N_21767,N_21628);
and U22060 (N_22060,N_21781,N_21788);
and U22061 (N_22061,N_21818,N_21605);
xor U22062 (N_22062,N_21756,N_21604);
xor U22063 (N_22063,N_21858,N_21784);
nor U22064 (N_22064,N_21667,N_21770);
or U22065 (N_22065,N_21839,N_21760);
xor U22066 (N_22066,N_21817,N_21780);
or U22067 (N_22067,N_21817,N_21834);
nor U22068 (N_22068,N_21852,N_21643);
and U22069 (N_22069,N_21874,N_21887);
and U22070 (N_22070,N_21718,N_21660);
nand U22071 (N_22071,N_21721,N_21689);
nand U22072 (N_22072,N_21749,N_21693);
and U22073 (N_22073,N_21746,N_21712);
nand U22074 (N_22074,N_21703,N_21695);
nand U22075 (N_22075,N_21611,N_21655);
or U22076 (N_22076,N_21736,N_21748);
or U22077 (N_22077,N_21740,N_21790);
nor U22078 (N_22078,N_21607,N_21681);
nor U22079 (N_22079,N_21616,N_21620);
nand U22080 (N_22080,N_21766,N_21705);
and U22081 (N_22081,N_21601,N_21605);
and U22082 (N_22082,N_21656,N_21749);
nand U22083 (N_22083,N_21658,N_21620);
nor U22084 (N_22084,N_21653,N_21882);
or U22085 (N_22085,N_21629,N_21751);
or U22086 (N_22086,N_21745,N_21731);
nand U22087 (N_22087,N_21668,N_21723);
nand U22088 (N_22088,N_21655,N_21779);
nor U22089 (N_22089,N_21808,N_21702);
xor U22090 (N_22090,N_21679,N_21623);
xor U22091 (N_22091,N_21748,N_21622);
xnor U22092 (N_22092,N_21686,N_21787);
or U22093 (N_22093,N_21811,N_21812);
nor U22094 (N_22094,N_21763,N_21883);
nor U22095 (N_22095,N_21862,N_21714);
or U22096 (N_22096,N_21686,N_21862);
and U22097 (N_22097,N_21780,N_21692);
and U22098 (N_22098,N_21687,N_21843);
nand U22099 (N_22099,N_21690,N_21634);
and U22100 (N_22100,N_21780,N_21725);
xor U22101 (N_22101,N_21629,N_21759);
and U22102 (N_22102,N_21638,N_21848);
nand U22103 (N_22103,N_21624,N_21774);
nor U22104 (N_22104,N_21775,N_21899);
xnor U22105 (N_22105,N_21602,N_21803);
nor U22106 (N_22106,N_21646,N_21605);
nand U22107 (N_22107,N_21875,N_21729);
nor U22108 (N_22108,N_21855,N_21792);
nand U22109 (N_22109,N_21763,N_21684);
nand U22110 (N_22110,N_21612,N_21646);
nand U22111 (N_22111,N_21617,N_21655);
nor U22112 (N_22112,N_21816,N_21677);
xor U22113 (N_22113,N_21782,N_21717);
xor U22114 (N_22114,N_21847,N_21896);
or U22115 (N_22115,N_21855,N_21760);
and U22116 (N_22116,N_21855,N_21701);
xor U22117 (N_22117,N_21717,N_21815);
or U22118 (N_22118,N_21823,N_21719);
nand U22119 (N_22119,N_21617,N_21647);
nand U22120 (N_22120,N_21842,N_21613);
and U22121 (N_22121,N_21789,N_21867);
nand U22122 (N_22122,N_21897,N_21718);
or U22123 (N_22123,N_21836,N_21656);
xnor U22124 (N_22124,N_21827,N_21669);
nor U22125 (N_22125,N_21664,N_21656);
nand U22126 (N_22126,N_21612,N_21635);
or U22127 (N_22127,N_21674,N_21727);
xor U22128 (N_22128,N_21656,N_21699);
or U22129 (N_22129,N_21898,N_21846);
and U22130 (N_22130,N_21796,N_21655);
or U22131 (N_22131,N_21715,N_21881);
nor U22132 (N_22132,N_21808,N_21810);
nor U22133 (N_22133,N_21680,N_21621);
and U22134 (N_22134,N_21806,N_21601);
nand U22135 (N_22135,N_21686,N_21802);
or U22136 (N_22136,N_21610,N_21863);
and U22137 (N_22137,N_21640,N_21683);
nand U22138 (N_22138,N_21716,N_21659);
or U22139 (N_22139,N_21704,N_21833);
xor U22140 (N_22140,N_21820,N_21723);
xnor U22141 (N_22141,N_21710,N_21659);
nor U22142 (N_22142,N_21790,N_21653);
nand U22143 (N_22143,N_21814,N_21770);
nor U22144 (N_22144,N_21721,N_21800);
and U22145 (N_22145,N_21617,N_21610);
nand U22146 (N_22146,N_21758,N_21823);
xnor U22147 (N_22147,N_21705,N_21889);
nand U22148 (N_22148,N_21879,N_21762);
nand U22149 (N_22149,N_21777,N_21617);
and U22150 (N_22150,N_21693,N_21616);
and U22151 (N_22151,N_21773,N_21731);
nor U22152 (N_22152,N_21748,N_21847);
nand U22153 (N_22153,N_21824,N_21634);
nand U22154 (N_22154,N_21880,N_21801);
or U22155 (N_22155,N_21642,N_21817);
nand U22156 (N_22156,N_21664,N_21773);
xnor U22157 (N_22157,N_21657,N_21632);
xor U22158 (N_22158,N_21779,N_21815);
nand U22159 (N_22159,N_21613,N_21805);
nand U22160 (N_22160,N_21816,N_21664);
xnor U22161 (N_22161,N_21853,N_21701);
and U22162 (N_22162,N_21793,N_21801);
and U22163 (N_22163,N_21815,N_21895);
xnor U22164 (N_22164,N_21715,N_21764);
and U22165 (N_22165,N_21650,N_21737);
or U22166 (N_22166,N_21664,N_21734);
nor U22167 (N_22167,N_21878,N_21672);
xor U22168 (N_22168,N_21810,N_21714);
nor U22169 (N_22169,N_21784,N_21717);
nor U22170 (N_22170,N_21869,N_21872);
nand U22171 (N_22171,N_21602,N_21749);
xor U22172 (N_22172,N_21819,N_21706);
xnor U22173 (N_22173,N_21729,N_21727);
xnor U22174 (N_22174,N_21696,N_21611);
and U22175 (N_22175,N_21641,N_21744);
and U22176 (N_22176,N_21688,N_21625);
or U22177 (N_22177,N_21698,N_21847);
nor U22178 (N_22178,N_21669,N_21864);
or U22179 (N_22179,N_21727,N_21770);
nor U22180 (N_22180,N_21723,N_21789);
nand U22181 (N_22181,N_21698,N_21892);
or U22182 (N_22182,N_21821,N_21876);
xnor U22183 (N_22183,N_21892,N_21774);
or U22184 (N_22184,N_21758,N_21784);
and U22185 (N_22185,N_21603,N_21771);
or U22186 (N_22186,N_21629,N_21677);
nor U22187 (N_22187,N_21750,N_21809);
nor U22188 (N_22188,N_21867,N_21725);
or U22189 (N_22189,N_21873,N_21742);
and U22190 (N_22190,N_21797,N_21661);
nand U22191 (N_22191,N_21827,N_21825);
or U22192 (N_22192,N_21628,N_21743);
xor U22193 (N_22193,N_21681,N_21878);
and U22194 (N_22194,N_21804,N_21616);
or U22195 (N_22195,N_21810,N_21797);
or U22196 (N_22196,N_21615,N_21602);
nor U22197 (N_22197,N_21758,N_21797);
nand U22198 (N_22198,N_21828,N_21682);
nand U22199 (N_22199,N_21855,N_21663);
xnor U22200 (N_22200,N_22158,N_22147);
and U22201 (N_22201,N_22018,N_22174);
xnor U22202 (N_22202,N_21991,N_22146);
nor U22203 (N_22203,N_22003,N_21921);
nor U22204 (N_22204,N_22191,N_22017);
xnor U22205 (N_22205,N_21904,N_22130);
nor U22206 (N_22206,N_21922,N_21956);
xnor U22207 (N_22207,N_22092,N_21937);
xor U22208 (N_22208,N_22133,N_21924);
nand U22209 (N_22209,N_22060,N_22079);
xnor U22210 (N_22210,N_22198,N_21915);
nor U22211 (N_22211,N_22179,N_22048);
and U22212 (N_22212,N_22023,N_22117);
nand U22213 (N_22213,N_21923,N_22169);
or U22214 (N_22214,N_21943,N_22166);
or U22215 (N_22215,N_22046,N_22099);
or U22216 (N_22216,N_22172,N_22096);
or U22217 (N_22217,N_21962,N_21905);
or U22218 (N_22218,N_22151,N_22129);
nor U22219 (N_22219,N_22119,N_22045);
nand U22220 (N_22220,N_22034,N_22141);
nand U22221 (N_22221,N_22140,N_22190);
and U22222 (N_22222,N_22156,N_22197);
xnor U22223 (N_22223,N_22013,N_22054);
nor U22224 (N_22224,N_22101,N_22116);
nor U22225 (N_22225,N_22095,N_22136);
nor U22226 (N_22226,N_22145,N_22187);
nor U22227 (N_22227,N_21910,N_22070);
xor U22228 (N_22228,N_21911,N_21955);
xnor U22229 (N_22229,N_22075,N_22028);
nand U22230 (N_22230,N_22186,N_22143);
or U22231 (N_22231,N_22098,N_22176);
and U22232 (N_22232,N_22196,N_22001);
or U22233 (N_22233,N_21996,N_22019);
nor U22234 (N_22234,N_22039,N_21981);
and U22235 (N_22235,N_21920,N_22020);
nand U22236 (N_22236,N_22009,N_21902);
nor U22237 (N_22237,N_21926,N_21928);
nor U22238 (N_22238,N_22193,N_21933);
nor U22239 (N_22239,N_21939,N_22144);
xor U22240 (N_22240,N_21901,N_22087);
nor U22241 (N_22241,N_21990,N_22059);
xor U22242 (N_22242,N_22067,N_21972);
nor U22243 (N_22243,N_21914,N_21957);
and U22244 (N_22244,N_22157,N_21995);
or U22245 (N_22245,N_22126,N_22026);
nand U22246 (N_22246,N_21919,N_22195);
nor U22247 (N_22247,N_22061,N_22097);
nand U22248 (N_22248,N_22153,N_21934);
or U22249 (N_22249,N_22065,N_22008);
or U22250 (N_22250,N_22063,N_22047);
nand U22251 (N_22251,N_22057,N_22024);
nor U22252 (N_22252,N_21997,N_21953);
nor U22253 (N_22253,N_22052,N_22085);
nor U22254 (N_22254,N_22149,N_22037);
nor U22255 (N_22255,N_21984,N_22007);
and U22256 (N_22256,N_22121,N_22104);
nand U22257 (N_22257,N_22053,N_22029);
and U22258 (N_22258,N_22081,N_22044);
or U22259 (N_22259,N_22139,N_22058);
or U22260 (N_22260,N_22069,N_22030);
nand U22261 (N_22261,N_21935,N_22161);
and U22262 (N_22262,N_22152,N_22163);
nand U22263 (N_22263,N_21968,N_22171);
xnor U22264 (N_22264,N_22120,N_22021);
nand U22265 (N_22265,N_22135,N_22011);
or U22266 (N_22266,N_21979,N_22064);
nand U22267 (N_22267,N_22132,N_22010);
or U22268 (N_22268,N_22073,N_22175);
nand U22269 (N_22269,N_22150,N_22033);
or U22270 (N_22270,N_21999,N_22056);
nand U22271 (N_22271,N_21983,N_22167);
xnor U22272 (N_22272,N_22183,N_22016);
or U22273 (N_22273,N_22015,N_22103);
xor U22274 (N_22274,N_21978,N_21974);
nor U22275 (N_22275,N_21982,N_22012);
or U22276 (N_22276,N_22041,N_21945);
and U22277 (N_22277,N_22173,N_22014);
nor U22278 (N_22278,N_22002,N_22086);
xor U22279 (N_22279,N_21932,N_21916);
xnor U22280 (N_22280,N_22102,N_22177);
and U22281 (N_22281,N_22199,N_21929);
nand U22282 (N_22282,N_22182,N_21927);
nand U22283 (N_22283,N_22027,N_21909);
and U22284 (N_22284,N_21963,N_21908);
nand U22285 (N_22285,N_21917,N_21987);
nor U22286 (N_22286,N_22124,N_22115);
nor U22287 (N_22287,N_21989,N_22131);
xnor U22288 (N_22288,N_22051,N_22168);
or U22289 (N_22289,N_21944,N_22050);
xor U22290 (N_22290,N_21947,N_22043);
and U22291 (N_22291,N_21942,N_21941);
or U22292 (N_22292,N_21970,N_21994);
or U22293 (N_22293,N_22185,N_22137);
and U22294 (N_22294,N_22093,N_21951);
xnor U22295 (N_22295,N_22154,N_21971);
or U22296 (N_22296,N_21975,N_21938);
or U22297 (N_22297,N_21985,N_22049);
nor U22298 (N_22298,N_22000,N_22071);
nor U22299 (N_22299,N_21969,N_21977);
or U22300 (N_22300,N_22122,N_22114);
and U22301 (N_22301,N_21965,N_22066);
nand U22302 (N_22302,N_22042,N_22089);
and U22303 (N_22303,N_21952,N_22080);
xnor U22304 (N_22304,N_21931,N_21961);
xor U22305 (N_22305,N_21912,N_22192);
xor U22306 (N_22306,N_22078,N_22106);
and U22307 (N_22307,N_22022,N_22025);
or U22308 (N_22308,N_22031,N_21925);
xnor U22309 (N_22309,N_21906,N_22148);
and U22310 (N_22310,N_21967,N_22112);
and U22311 (N_22311,N_22118,N_22194);
nor U22312 (N_22312,N_22100,N_22083);
xor U22313 (N_22313,N_21950,N_21954);
xnor U22314 (N_22314,N_22091,N_22108);
xnor U22315 (N_22315,N_21900,N_21930);
or U22316 (N_22316,N_21964,N_22036);
xor U22317 (N_22317,N_21918,N_22084);
nor U22318 (N_22318,N_21936,N_21992);
nor U22319 (N_22319,N_21980,N_22178);
xnor U22320 (N_22320,N_22038,N_21973);
nand U22321 (N_22321,N_22090,N_21986);
xnor U22322 (N_22322,N_22159,N_22035);
or U22323 (N_22323,N_22170,N_21949);
and U22324 (N_22324,N_22164,N_22105);
nand U22325 (N_22325,N_22127,N_22055);
or U22326 (N_22326,N_22072,N_22125);
nor U22327 (N_22327,N_22160,N_22005);
and U22328 (N_22328,N_22188,N_21940);
nor U22329 (N_22329,N_21913,N_22040);
nor U22330 (N_22330,N_22107,N_21976);
nand U22331 (N_22331,N_22076,N_22077);
and U22332 (N_22332,N_22123,N_21946);
nand U22333 (N_22333,N_21958,N_22181);
nor U22334 (N_22334,N_22184,N_22111);
xnor U22335 (N_22335,N_22006,N_22180);
nor U22336 (N_22336,N_22189,N_22109);
and U22337 (N_22337,N_21988,N_21993);
and U22338 (N_22338,N_22138,N_22162);
xor U22339 (N_22339,N_22094,N_21948);
or U22340 (N_22340,N_22113,N_22068);
and U22341 (N_22341,N_22082,N_22032);
and U22342 (N_22342,N_21959,N_22074);
or U22343 (N_22343,N_22134,N_22062);
xnor U22344 (N_22344,N_21998,N_21903);
or U22345 (N_22345,N_22128,N_22142);
xor U22346 (N_22346,N_22165,N_22155);
xnor U22347 (N_22347,N_22004,N_22088);
nor U22348 (N_22348,N_21960,N_22110);
or U22349 (N_22349,N_21907,N_21966);
and U22350 (N_22350,N_21907,N_22130);
and U22351 (N_22351,N_22009,N_22034);
and U22352 (N_22352,N_21976,N_22093);
or U22353 (N_22353,N_22091,N_22119);
or U22354 (N_22354,N_21953,N_22094);
nor U22355 (N_22355,N_22105,N_22084);
nand U22356 (N_22356,N_22128,N_22129);
nand U22357 (N_22357,N_22133,N_21948);
nor U22358 (N_22358,N_21992,N_22063);
xnor U22359 (N_22359,N_22149,N_22028);
xnor U22360 (N_22360,N_22189,N_21903);
nor U22361 (N_22361,N_21943,N_22164);
xor U22362 (N_22362,N_22033,N_22043);
or U22363 (N_22363,N_22043,N_21985);
xor U22364 (N_22364,N_22110,N_22042);
or U22365 (N_22365,N_22005,N_22032);
and U22366 (N_22366,N_22113,N_21946);
nor U22367 (N_22367,N_22188,N_21919);
xnor U22368 (N_22368,N_21919,N_21980);
nor U22369 (N_22369,N_22130,N_22097);
or U22370 (N_22370,N_22108,N_21998);
nand U22371 (N_22371,N_22196,N_22132);
and U22372 (N_22372,N_22087,N_22062);
nand U22373 (N_22373,N_22137,N_22082);
and U22374 (N_22374,N_22032,N_22079);
xnor U22375 (N_22375,N_22013,N_21904);
nand U22376 (N_22376,N_22169,N_22186);
nand U22377 (N_22377,N_22084,N_22119);
nor U22378 (N_22378,N_22122,N_21934);
nor U22379 (N_22379,N_21940,N_22049);
and U22380 (N_22380,N_22153,N_22011);
nor U22381 (N_22381,N_22012,N_21917);
nor U22382 (N_22382,N_22187,N_21997);
xor U22383 (N_22383,N_22188,N_22076);
nor U22384 (N_22384,N_22113,N_22182);
xor U22385 (N_22385,N_22042,N_21966);
nand U22386 (N_22386,N_22115,N_22168);
xor U22387 (N_22387,N_22066,N_22117);
nand U22388 (N_22388,N_21949,N_22004);
nand U22389 (N_22389,N_22120,N_21953);
nand U22390 (N_22390,N_21978,N_22053);
nand U22391 (N_22391,N_22057,N_21948);
nand U22392 (N_22392,N_22016,N_21909);
or U22393 (N_22393,N_22100,N_22056);
nor U22394 (N_22394,N_22080,N_22138);
or U22395 (N_22395,N_21985,N_21987);
nor U22396 (N_22396,N_22059,N_21906);
nor U22397 (N_22397,N_22137,N_22062);
nand U22398 (N_22398,N_22178,N_22031);
nand U22399 (N_22399,N_22062,N_22175);
or U22400 (N_22400,N_21929,N_21978);
nor U22401 (N_22401,N_22144,N_22105);
nand U22402 (N_22402,N_21951,N_21954);
nor U22403 (N_22403,N_22185,N_22093);
nor U22404 (N_22404,N_22063,N_22010);
xor U22405 (N_22405,N_21933,N_22108);
xnor U22406 (N_22406,N_21930,N_21941);
or U22407 (N_22407,N_21964,N_21993);
nor U22408 (N_22408,N_21969,N_22061);
nor U22409 (N_22409,N_22026,N_22079);
nor U22410 (N_22410,N_21985,N_22129);
nor U22411 (N_22411,N_22168,N_22055);
xor U22412 (N_22412,N_22117,N_21928);
nor U22413 (N_22413,N_21931,N_22031);
and U22414 (N_22414,N_21935,N_22068);
and U22415 (N_22415,N_21909,N_21930);
nand U22416 (N_22416,N_22176,N_22090);
xor U22417 (N_22417,N_21957,N_21905);
nor U22418 (N_22418,N_21995,N_22040);
or U22419 (N_22419,N_21915,N_22072);
nor U22420 (N_22420,N_22081,N_21948);
nor U22421 (N_22421,N_22197,N_21943);
and U22422 (N_22422,N_22110,N_21950);
xnor U22423 (N_22423,N_21955,N_22105);
nand U22424 (N_22424,N_21942,N_22010);
nand U22425 (N_22425,N_22069,N_22195);
and U22426 (N_22426,N_22158,N_22188);
nand U22427 (N_22427,N_21995,N_22054);
and U22428 (N_22428,N_21988,N_22028);
and U22429 (N_22429,N_22105,N_22054);
and U22430 (N_22430,N_22007,N_21936);
xnor U22431 (N_22431,N_22043,N_22183);
and U22432 (N_22432,N_22147,N_22048);
nor U22433 (N_22433,N_21900,N_22080);
xnor U22434 (N_22434,N_22176,N_22077);
nor U22435 (N_22435,N_22103,N_22092);
or U22436 (N_22436,N_22050,N_21929);
and U22437 (N_22437,N_22079,N_22160);
nor U22438 (N_22438,N_22112,N_21904);
nor U22439 (N_22439,N_22003,N_21904);
and U22440 (N_22440,N_22008,N_21969);
xnor U22441 (N_22441,N_22049,N_21943);
or U22442 (N_22442,N_22100,N_21976);
or U22443 (N_22443,N_21901,N_22149);
xnor U22444 (N_22444,N_22125,N_22073);
and U22445 (N_22445,N_22152,N_22064);
and U22446 (N_22446,N_21917,N_22158);
nor U22447 (N_22447,N_21922,N_21950);
nand U22448 (N_22448,N_22096,N_22157);
or U22449 (N_22449,N_22194,N_22042);
xnor U22450 (N_22450,N_21997,N_22093);
or U22451 (N_22451,N_22110,N_21938);
or U22452 (N_22452,N_22064,N_21900);
and U22453 (N_22453,N_21931,N_22106);
and U22454 (N_22454,N_22015,N_21979);
xor U22455 (N_22455,N_22165,N_22034);
nand U22456 (N_22456,N_21935,N_21993);
nor U22457 (N_22457,N_22062,N_22050);
and U22458 (N_22458,N_22061,N_22098);
xor U22459 (N_22459,N_22010,N_21970);
xor U22460 (N_22460,N_22017,N_21945);
xnor U22461 (N_22461,N_22036,N_22019);
and U22462 (N_22462,N_22056,N_22121);
nor U22463 (N_22463,N_22041,N_22035);
xor U22464 (N_22464,N_21965,N_22120);
nand U22465 (N_22465,N_21932,N_21995);
and U22466 (N_22466,N_22033,N_21917);
and U22467 (N_22467,N_22106,N_22031);
and U22468 (N_22468,N_22020,N_22063);
xor U22469 (N_22469,N_21946,N_21913);
xnor U22470 (N_22470,N_21943,N_22079);
and U22471 (N_22471,N_22014,N_22085);
nand U22472 (N_22472,N_21965,N_21945);
and U22473 (N_22473,N_22065,N_22162);
and U22474 (N_22474,N_22003,N_22099);
and U22475 (N_22475,N_22156,N_22096);
or U22476 (N_22476,N_22143,N_21983);
or U22477 (N_22477,N_22153,N_22073);
xnor U22478 (N_22478,N_22140,N_22132);
or U22479 (N_22479,N_22060,N_22059);
and U22480 (N_22480,N_22075,N_21930);
xnor U22481 (N_22481,N_22171,N_22087);
nor U22482 (N_22482,N_22103,N_22158);
nand U22483 (N_22483,N_22128,N_22014);
xnor U22484 (N_22484,N_22019,N_22138);
nor U22485 (N_22485,N_22115,N_21987);
nor U22486 (N_22486,N_21992,N_22080);
or U22487 (N_22487,N_22141,N_21966);
or U22488 (N_22488,N_21911,N_21937);
xor U22489 (N_22489,N_22152,N_21923);
or U22490 (N_22490,N_22108,N_22061);
or U22491 (N_22491,N_22142,N_22119);
and U22492 (N_22492,N_22062,N_22095);
nor U22493 (N_22493,N_22129,N_22115);
or U22494 (N_22494,N_22038,N_22033);
nand U22495 (N_22495,N_22034,N_22022);
nand U22496 (N_22496,N_21998,N_21939);
and U22497 (N_22497,N_22044,N_22037);
nor U22498 (N_22498,N_22124,N_21910);
nand U22499 (N_22499,N_22090,N_21925);
nor U22500 (N_22500,N_22323,N_22371);
nor U22501 (N_22501,N_22353,N_22322);
nand U22502 (N_22502,N_22212,N_22204);
xnor U22503 (N_22503,N_22329,N_22447);
and U22504 (N_22504,N_22409,N_22311);
or U22505 (N_22505,N_22424,N_22232);
xor U22506 (N_22506,N_22463,N_22368);
nand U22507 (N_22507,N_22356,N_22222);
and U22508 (N_22508,N_22313,N_22396);
xor U22509 (N_22509,N_22416,N_22233);
or U22510 (N_22510,N_22317,N_22487);
nor U22511 (N_22511,N_22275,N_22474);
nand U22512 (N_22512,N_22403,N_22370);
nand U22513 (N_22513,N_22456,N_22334);
xnor U22514 (N_22514,N_22459,N_22461);
xnor U22515 (N_22515,N_22220,N_22293);
or U22516 (N_22516,N_22399,N_22227);
nor U22517 (N_22517,N_22333,N_22235);
nand U22518 (N_22518,N_22401,N_22236);
nand U22519 (N_22519,N_22216,N_22338);
nor U22520 (N_22520,N_22340,N_22259);
nor U22521 (N_22521,N_22467,N_22309);
nor U22522 (N_22522,N_22328,N_22346);
and U22523 (N_22523,N_22288,N_22432);
xnor U22524 (N_22524,N_22408,N_22348);
nor U22525 (N_22525,N_22206,N_22225);
xor U22526 (N_22526,N_22376,N_22491);
xnor U22527 (N_22527,N_22217,N_22224);
nor U22528 (N_22528,N_22411,N_22367);
xor U22529 (N_22529,N_22238,N_22226);
or U22530 (N_22530,N_22462,N_22294);
and U22531 (N_22531,N_22319,N_22359);
xor U22532 (N_22532,N_22285,N_22374);
and U22533 (N_22533,N_22499,N_22380);
nand U22534 (N_22534,N_22373,N_22347);
or U22535 (N_22535,N_22451,N_22444);
or U22536 (N_22536,N_22243,N_22422);
and U22537 (N_22537,N_22485,N_22395);
xor U22538 (N_22538,N_22272,N_22264);
and U22539 (N_22539,N_22415,N_22321);
or U22540 (N_22540,N_22282,N_22394);
xnor U22541 (N_22541,N_22381,N_22363);
nand U22542 (N_22542,N_22427,N_22476);
nand U22543 (N_22543,N_22247,N_22286);
or U22544 (N_22544,N_22495,N_22343);
or U22545 (N_22545,N_22426,N_22281);
and U22546 (N_22546,N_22336,N_22443);
nor U22547 (N_22547,N_22301,N_22267);
or U22548 (N_22548,N_22488,N_22290);
nand U22549 (N_22549,N_22213,N_22218);
and U22550 (N_22550,N_22482,N_22231);
xnor U22551 (N_22551,N_22389,N_22470);
nor U22552 (N_22552,N_22254,N_22484);
or U22553 (N_22553,N_22413,N_22450);
nor U22554 (N_22554,N_22240,N_22208);
or U22555 (N_22555,N_22246,N_22406);
and U22556 (N_22556,N_22445,N_22349);
and U22557 (N_22557,N_22404,N_22402);
nor U22558 (N_22558,N_22345,N_22420);
or U22559 (N_22559,N_22478,N_22361);
or U22560 (N_22560,N_22250,N_22255);
nor U22561 (N_22561,N_22365,N_22475);
and U22562 (N_22562,N_22452,N_22332);
xnor U22563 (N_22563,N_22397,N_22439);
xnor U22564 (N_22564,N_22364,N_22229);
xor U22565 (N_22565,N_22493,N_22291);
nor U22566 (N_22566,N_22486,N_22419);
or U22567 (N_22567,N_22350,N_22228);
xor U22568 (N_22568,N_22407,N_22339);
and U22569 (N_22569,N_22418,N_22400);
nor U22570 (N_22570,N_22266,N_22239);
nand U22571 (N_22571,N_22383,N_22352);
xnor U22572 (N_22572,N_22477,N_22385);
nand U22573 (N_22573,N_22269,N_22302);
xnor U22574 (N_22574,N_22351,N_22466);
or U22575 (N_22575,N_22341,N_22360);
nor U22576 (N_22576,N_22425,N_22318);
and U22577 (N_22577,N_22230,N_22468);
xor U22578 (N_22578,N_22417,N_22314);
or U22579 (N_22579,N_22457,N_22260);
or U22580 (N_22580,N_22342,N_22257);
nand U22581 (N_22581,N_22244,N_22201);
nor U22582 (N_22582,N_22271,N_22209);
nand U22583 (N_22583,N_22200,N_22496);
and U22584 (N_22584,N_22378,N_22211);
nor U22585 (N_22585,N_22423,N_22335);
and U22586 (N_22586,N_22440,N_22472);
nand U22587 (N_22587,N_22388,N_22289);
nor U22588 (N_22588,N_22303,N_22287);
and U22589 (N_22589,N_22366,N_22315);
and U22590 (N_22590,N_22438,N_22481);
nor U22591 (N_22591,N_22256,N_22306);
xnor U22592 (N_22592,N_22308,N_22249);
and U22593 (N_22593,N_22434,N_22494);
nand U22594 (N_22594,N_22448,N_22221);
and U22595 (N_22595,N_22435,N_22262);
nand U22596 (N_22596,N_22316,N_22391);
or U22597 (N_22597,N_22202,N_22312);
or U22598 (N_22598,N_22458,N_22324);
xor U22599 (N_22599,N_22483,N_22362);
nor U22600 (N_22600,N_22207,N_22277);
nand U22601 (N_22601,N_22398,N_22410);
and U22602 (N_22602,N_22377,N_22453);
and U22603 (N_22603,N_22283,N_22203);
nor U22604 (N_22604,N_22490,N_22325);
or U22605 (N_22605,N_22492,N_22384);
nand U22606 (N_22606,N_22223,N_22465);
or U22607 (N_22607,N_22274,N_22390);
nor U22608 (N_22608,N_22414,N_22446);
nor U22609 (N_22609,N_22253,N_22354);
xor U22610 (N_22610,N_22479,N_22480);
or U22611 (N_22611,N_22421,N_22442);
nor U22612 (N_22612,N_22412,N_22358);
nor U22613 (N_22613,N_22429,N_22428);
or U22614 (N_22614,N_22449,N_22299);
or U22615 (N_22615,N_22387,N_22386);
nand U22616 (N_22616,N_22326,N_22248);
xnor U22617 (N_22617,N_22469,N_22292);
xor U22618 (N_22618,N_22320,N_22245);
xnor U22619 (N_22619,N_22276,N_22455);
nand U22620 (N_22620,N_22437,N_22344);
xor U22621 (N_22621,N_22252,N_22392);
xnor U22622 (N_22622,N_22251,N_22278);
xnor U22623 (N_22623,N_22498,N_22237);
or U22624 (N_22624,N_22430,N_22219);
or U22625 (N_22625,N_22265,N_22305);
nor U22626 (N_22626,N_22357,N_22273);
xnor U22627 (N_22627,N_22270,N_22241);
or U22628 (N_22628,N_22375,N_22279);
nand U22629 (N_22629,N_22261,N_22497);
nor U22630 (N_22630,N_22436,N_22297);
or U22631 (N_22631,N_22337,N_22331);
xnor U22632 (N_22632,N_22215,N_22355);
or U22633 (N_22633,N_22307,N_22441);
nor U22634 (N_22634,N_22379,N_22464);
nor U22635 (N_22635,N_22473,N_22280);
and U22636 (N_22636,N_22327,N_22330);
or U22637 (N_22637,N_22431,N_22369);
and U22638 (N_22638,N_22295,N_22460);
nor U22639 (N_22639,N_22471,N_22304);
nor U22640 (N_22640,N_22284,N_22234);
xor U22641 (N_22641,N_22382,N_22454);
and U22642 (N_22642,N_22300,N_22372);
xnor U22643 (N_22643,N_22298,N_22405);
and U22644 (N_22644,N_22205,N_22393);
nor U22645 (N_22645,N_22242,N_22263);
xnor U22646 (N_22646,N_22268,N_22310);
nand U22647 (N_22647,N_22433,N_22214);
and U22648 (N_22648,N_22258,N_22296);
and U22649 (N_22649,N_22489,N_22210);
or U22650 (N_22650,N_22408,N_22236);
or U22651 (N_22651,N_22294,N_22240);
and U22652 (N_22652,N_22498,N_22252);
and U22653 (N_22653,N_22351,N_22291);
xnor U22654 (N_22654,N_22452,N_22348);
xnor U22655 (N_22655,N_22326,N_22222);
nand U22656 (N_22656,N_22260,N_22462);
and U22657 (N_22657,N_22377,N_22260);
and U22658 (N_22658,N_22347,N_22482);
and U22659 (N_22659,N_22223,N_22387);
xnor U22660 (N_22660,N_22329,N_22335);
nor U22661 (N_22661,N_22414,N_22307);
and U22662 (N_22662,N_22222,N_22394);
xnor U22663 (N_22663,N_22279,N_22453);
xor U22664 (N_22664,N_22210,N_22438);
and U22665 (N_22665,N_22397,N_22213);
xnor U22666 (N_22666,N_22207,N_22359);
nor U22667 (N_22667,N_22284,N_22375);
and U22668 (N_22668,N_22431,N_22303);
nand U22669 (N_22669,N_22416,N_22253);
and U22670 (N_22670,N_22484,N_22307);
xnor U22671 (N_22671,N_22449,N_22239);
and U22672 (N_22672,N_22218,N_22473);
nand U22673 (N_22673,N_22224,N_22399);
or U22674 (N_22674,N_22389,N_22479);
nor U22675 (N_22675,N_22321,N_22389);
nand U22676 (N_22676,N_22420,N_22452);
nand U22677 (N_22677,N_22410,N_22223);
or U22678 (N_22678,N_22317,N_22323);
or U22679 (N_22679,N_22300,N_22347);
nor U22680 (N_22680,N_22487,N_22461);
nor U22681 (N_22681,N_22422,N_22239);
nand U22682 (N_22682,N_22370,N_22419);
or U22683 (N_22683,N_22430,N_22334);
xnor U22684 (N_22684,N_22404,N_22215);
and U22685 (N_22685,N_22394,N_22228);
xor U22686 (N_22686,N_22361,N_22364);
nor U22687 (N_22687,N_22200,N_22288);
nor U22688 (N_22688,N_22236,N_22430);
and U22689 (N_22689,N_22209,N_22264);
and U22690 (N_22690,N_22488,N_22201);
nor U22691 (N_22691,N_22279,N_22442);
nand U22692 (N_22692,N_22459,N_22421);
nand U22693 (N_22693,N_22359,N_22345);
or U22694 (N_22694,N_22347,N_22292);
or U22695 (N_22695,N_22229,N_22248);
nand U22696 (N_22696,N_22362,N_22267);
xnor U22697 (N_22697,N_22313,N_22489);
nor U22698 (N_22698,N_22393,N_22467);
xor U22699 (N_22699,N_22244,N_22243);
xnor U22700 (N_22700,N_22255,N_22440);
nor U22701 (N_22701,N_22360,N_22244);
and U22702 (N_22702,N_22262,N_22463);
nand U22703 (N_22703,N_22305,N_22429);
nand U22704 (N_22704,N_22331,N_22225);
xnor U22705 (N_22705,N_22444,N_22203);
nor U22706 (N_22706,N_22250,N_22204);
nand U22707 (N_22707,N_22257,N_22447);
and U22708 (N_22708,N_22255,N_22287);
and U22709 (N_22709,N_22429,N_22348);
and U22710 (N_22710,N_22415,N_22472);
or U22711 (N_22711,N_22228,N_22300);
nand U22712 (N_22712,N_22405,N_22321);
xor U22713 (N_22713,N_22400,N_22300);
and U22714 (N_22714,N_22277,N_22468);
nor U22715 (N_22715,N_22243,N_22339);
nor U22716 (N_22716,N_22366,N_22261);
or U22717 (N_22717,N_22476,N_22245);
nand U22718 (N_22718,N_22352,N_22477);
nand U22719 (N_22719,N_22436,N_22211);
nand U22720 (N_22720,N_22452,N_22210);
and U22721 (N_22721,N_22229,N_22345);
nand U22722 (N_22722,N_22265,N_22237);
or U22723 (N_22723,N_22434,N_22265);
or U22724 (N_22724,N_22408,N_22221);
xor U22725 (N_22725,N_22219,N_22396);
or U22726 (N_22726,N_22371,N_22447);
nand U22727 (N_22727,N_22450,N_22404);
nor U22728 (N_22728,N_22291,N_22300);
xor U22729 (N_22729,N_22472,N_22346);
or U22730 (N_22730,N_22211,N_22306);
and U22731 (N_22731,N_22449,N_22448);
nand U22732 (N_22732,N_22444,N_22473);
xnor U22733 (N_22733,N_22477,N_22216);
nand U22734 (N_22734,N_22284,N_22313);
and U22735 (N_22735,N_22368,N_22461);
xor U22736 (N_22736,N_22335,N_22489);
xnor U22737 (N_22737,N_22498,N_22325);
and U22738 (N_22738,N_22414,N_22390);
nand U22739 (N_22739,N_22481,N_22231);
xnor U22740 (N_22740,N_22257,N_22292);
and U22741 (N_22741,N_22342,N_22434);
and U22742 (N_22742,N_22463,N_22406);
nand U22743 (N_22743,N_22476,N_22447);
nor U22744 (N_22744,N_22322,N_22270);
nor U22745 (N_22745,N_22213,N_22369);
nand U22746 (N_22746,N_22409,N_22302);
and U22747 (N_22747,N_22381,N_22255);
and U22748 (N_22748,N_22457,N_22286);
xor U22749 (N_22749,N_22283,N_22455);
nor U22750 (N_22750,N_22391,N_22215);
nor U22751 (N_22751,N_22362,N_22444);
nor U22752 (N_22752,N_22294,N_22392);
nand U22753 (N_22753,N_22378,N_22388);
and U22754 (N_22754,N_22382,N_22462);
or U22755 (N_22755,N_22262,N_22216);
nor U22756 (N_22756,N_22301,N_22403);
and U22757 (N_22757,N_22269,N_22230);
nand U22758 (N_22758,N_22242,N_22235);
nand U22759 (N_22759,N_22444,N_22478);
nand U22760 (N_22760,N_22329,N_22277);
and U22761 (N_22761,N_22461,N_22373);
and U22762 (N_22762,N_22246,N_22492);
and U22763 (N_22763,N_22397,N_22339);
nand U22764 (N_22764,N_22439,N_22235);
and U22765 (N_22765,N_22453,N_22396);
xor U22766 (N_22766,N_22203,N_22480);
or U22767 (N_22767,N_22258,N_22208);
nor U22768 (N_22768,N_22256,N_22281);
and U22769 (N_22769,N_22308,N_22342);
xor U22770 (N_22770,N_22350,N_22438);
or U22771 (N_22771,N_22411,N_22279);
nor U22772 (N_22772,N_22267,N_22282);
nand U22773 (N_22773,N_22463,N_22286);
nand U22774 (N_22774,N_22318,N_22495);
xnor U22775 (N_22775,N_22340,N_22339);
nand U22776 (N_22776,N_22299,N_22278);
or U22777 (N_22777,N_22288,N_22446);
and U22778 (N_22778,N_22350,N_22408);
nor U22779 (N_22779,N_22395,N_22324);
nand U22780 (N_22780,N_22243,N_22421);
nor U22781 (N_22781,N_22361,N_22495);
nand U22782 (N_22782,N_22309,N_22475);
nand U22783 (N_22783,N_22245,N_22238);
or U22784 (N_22784,N_22369,N_22222);
xor U22785 (N_22785,N_22338,N_22212);
and U22786 (N_22786,N_22340,N_22226);
xnor U22787 (N_22787,N_22231,N_22249);
nor U22788 (N_22788,N_22394,N_22486);
nor U22789 (N_22789,N_22213,N_22371);
nor U22790 (N_22790,N_22272,N_22422);
and U22791 (N_22791,N_22449,N_22335);
nor U22792 (N_22792,N_22445,N_22351);
or U22793 (N_22793,N_22229,N_22458);
xor U22794 (N_22794,N_22324,N_22427);
and U22795 (N_22795,N_22438,N_22201);
nor U22796 (N_22796,N_22271,N_22348);
nor U22797 (N_22797,N_22437,N_22476);
and U22798 (N_22798,N_22377,N_22462);
nand U22799 (N_22799,N_22403,N_22319);
xnor U22800 (N_22800,N_22558,N_22703);
nand U22801 (N_22801,N_22733,N_22764);
xor U22802 (N_22802,N_22680,N_22666);
or U22803 (N_22803,N_22785,N_22753);
or U22804 (N_22804,N_22645,N_22531);
xnor U22805 (N_22805,N_22561,N_22503);
nor U22806 (N_22806,N_22588,N_22735);
or U22807 (N_22807,N_22799,N_22501);
nor U22808 (N_22808,N_22623,N_22739);
and U22809 (N_22809,N_22508,N_22513);
xor U22810 (N_22810,N_22563,N_22571);
or U22811 (N_22811,N_22604,N_22796);
nand U22812 (N_22812,N_22759,N_22629);
or U22813 (N_22813,N_22639,N_22589);
nand U22814 (N_22814,N_22697,N_22579);
xnor U22815 (N_22815,N_22732,N_22590);
nand U22816 (N_22816,N_22632,N_22784);
and U22817 (N_22817,N_22675,N_22611);
or U22818 (N_22818,N_22706,N_22622);
xor U22819 (N_22819,N_22567,N_22650);
nor U22820 (N_22820,N_22520,N_22660);
nand U22821 (N_22821,N_22718,N_22711);
or U22822 (N_22822,N_22747,N_22748);
and U22823 (N_22823,N_22762,N_22528);
or U22824 (N_22824,N_22519,N_22720);
xor U22825 (N_22825,N_22782,N_22670);
nor U22826 (N_22826,N_22610,N_22510);
nor U22827 (N_22827,N_22730,N_22790);
or U22828 (N_22828,N_22668,N_22545);
nand U22829 (N_22829,N_22564,N_22701);
nand U22830 (N_22830,N_22712,N_22690);
or U22831 (N_22831,N_22793,N_22540);
and U22832 (N_22832,N_22797,N_22667);
nand U22833 (N_22833,N_22631,N_22500);
or U22834 (N_22834,N_22647,N_22757);
or U22835 (N_22835,N_22620,N_22769);
xnor U22836 (N_22836,N_22778,N_22634);
or U22837 (N_22837,N_22615,N_22582);
nor U22838 (N_22838,N_22694,N_22641);
and U22839 (N_22839,N_22532,N_22774);
nand U22840 (N_22840,N_22648,N_22717);
nor U22841 (N_22841,N_22673,N_22502);
or U22842 (N_22842,N_22614,N_22691);
xnor U22843 (N_22843,N_22552,N_22524);
nand U22844 (N_22844,N_22521,N_22750);
nand U22845 (N_22845,N_22550,N_22656);
nor U22846 (N_22846,N_22755,N_22683);
nand U22847 (N_22847,N_22578,N_22533);
nor U22848 (N_22848,N_22577,N_22781);
or U22849 (N_22849,N_22530,N_22773);
and U22850 (N_22850,N_22713,N_22637);
nor U22851 (N_22851,N_22547,N_22643);
xor U22852 (N_22852,N_22758,N_22704);
and U22853 (N_22853,N_22723,N_22583);
and U22854 (N_22854,N_22557,N_22601);
xnor U22855 (N_22855,N_22655,N_22761);
nand U22856 (N_22856,N_22738,N_22572);
and U22857 (N_22857,N_22657,N_22731);
nor U22858 (N_22858,N_22576,N_22736);
nand U22859 (N_22859,N_22776,N_22535);
nor U22860 (N_22860,N_22646,N_22662);
xnor U22861 (N_22861,N_22585,N_22798);
nand U22862 (N_22862,N_22708,N_22659);
nor U22863 (N_22863,N_22526,N_22630);
nor U22864 (N_22864,N_22682,N_22702);
or U22865 (N_22865,N_22743,N_22746);
xnor U22866 (N_22866,N_22763,N_22543);
nor U22867 (N_22867,N_22607,N_22672);
nand U22868 (N_22868,N_22676,N_22695);
xor U22869 (N_22869,N_22726,N_22688);
nor U22870 (N_22870,N_22555,N_22644);
nand U22871 (N_22871,N_22621,N_22551);
xor U22872 (N_22872,N_22581,N_22674);
and U22873 (N_22873,N_22664,N_22504);
or U22874 (N_22874,N_22569,N_22779);
xnor U22875 (N_22875,N_22618,N_22619);
xor U22876 (N_22876,N_22783,N_22651);
nor U22877 (N_22877,N_22721,N_22625);
xnor U22878 (N_22878,N_22517,N_22600);
and U22879 (N_22879,N_22705,N_22699);
or U22880 (N_22880,N_22693,N_22603);
nor U22881 (N_22881,N_22679,N_22587);
nand U22882 (N_22882,N_22516,N_22669);
and U22883 (N_22883,N_22624,N_22766);
nand U22884 (N_22884,N_22709,N_22678);
or U22885 (N_22885,N_22653,N_22649);
nor U22886 (N_22886,N_22792,N_22642);
or U22887 (N_22887,N_22608,N_22595);
xor U22888 (N_22888,N_22724,N_22715);
nor U22889 (N_22889,N_22770,N_22789);
nand U22890 (N_22890,N_22714,N_22627);
nor U22891 (N_22891,N_22698,N_22740);
or U22892 (N_22892,N_22514,N_22518);
and U22893 (N_22893,N_22525,N_22751);
or U22894 (N_22894,N_22719,N_22548);
and U22895 (N_22895,N_22538,N_22575);
xor U22896 (N_22896,N_22754,N_22775);
or U22897 (N_22897,N_22768,N_22628);
xor U22898 (N_22898,N_22729,N_22554);
nand U22899 (N_22899,N_22635,N_22786);
xor U22900 (N_22900,N_22559,N_22710);
xnor U22901 (N_22901,N_22725,N_22529);
and U22902 (N_22902,N_22599,N_22565);
nand U22903 (N_22903,N_22586,N_22606);
or U22904 (N_22904,N_22522,N_22507);
nor U22905 (N_22905,N_22686,N_22534);
xor U22906 (N_22906,N_22602,N_22546);
xnor U22907 (N_22907,N_22605,N_22593);
nand U22908 (N_22908,N_22560,N_22512);
nor U22909 (N_22909,N_22791,N_22638);
nand U22910 (N_22910,N_22787,N_22573);
and U22911 (N_22911,N_22661,N_22696);
and U22912 (N_22912,N_22592,N_22570);
nor U22913 (N_22913,N_22745,N_22542);
xor U22914 (N_22914,N_22752,N_22794);
xnor U22915 (N_22915,N_22511,N_22734);
xnor U22916 (N_22916,N_22741,N_22671);
or U22917 (N_22917,N_22568,N_22658);
or U22918 (N_22918,N_22566,N_22515);
or U22919 (N_22919,N_22767,N_22665);
xor U22920 (N_22920,N_22689,N_22765);
xnor U22921 (N_22921,N_22509,N_22539);
xnor U22922 (N_22922,N_22777,N_22609);
xor U22923 (N_22923,N_22737,N_22788);
nor U22924 (N_22924,N_22700,N_22596);
or U22925 (N_22925,N_22687,N_22684);
nand U22926 (N_22926,N_22584,N_22633);
and U22927 (N_22927,N_22640,N_22553);
nor U22928 (N_22928,N_22537,N_22574);
nand U22929 (N_22929,N_22780,N_22685);
and U22930 (N_22930,N_22727,N_22598);
or U22931 (N_22931,N_22742,N_22505);
nand U22932 (N_22932,N_22613,N_22652);
nand U22933 (N_22933,N_22771,N_22677);
or U22934 (N_22934,N_22692,N_22549);
or U22935 (N_22935,N_22728,N_22556);
nor U22936 (N_22936,N_22636,N_22707);
or U22937 (N_22937,N_22626,N_22744);
xnor U22938 (N_22938,N_22663,N_22591);
or U22939 (N_22939,N_22536,N_22594);
xnor U22940 (N_22940,N_22523,N_22795);
and U22941 (N_22941,N_22722,N_22617);
and U22942 (N_22942,N_22756,N_22681);
or U22943 (N_22943,N_22580,N_22597);
nand U22944 (N_22944,N_22544,N_22716);
and U22945 (N_22945,N_22506,N_22541);
nand U22946 (N_22946,N_22616,N_22749);
or U22947 (N_22947,N_22760,N_22654);
nand U22948 (N_22948,N_22772,N_22527);
xor U22949 (N_22949,N_22612,N_22562);
xnor U22950 (N_22950,N_22773,N_22719);
and U22951 (N_22951,N_22550,N_22707);
nor U22952 (N_22952,N_22632,N_22578);
nand U22953 (N_22953,N_22737,N_22557);
nor U22954 (N_22954,N_22593,N_22733);
nand U22955 (N_22955,N_22775,N_22611);
and U22956 (N_22956,N_22643,N_22629);
xnor U22957 (N_22957,N_22631,N_22506);
and U22958 (N_22958,N_22594,N_22743);
xor U22959 (N_22959,N_22774,N_22690);
nand U22960 (N_22960,N_22503,N_22649);
xnor U22961 (N_22961,N_22582,N_22630);
nor U22962 (N_22962,N_22753,N_22627);
or U22963 (N_22963,N_22672,N_22780);
nand U22964 (N_22964,N_22708,N_22562);
xnor U22965 (N_22965,N_22791,N_22795);
nor U22966 (N_22966,N_22621,N_22591);
and U22967 (N_22967,N_22771,N_22681);
nand U22968 (N_22968,N_22769,N_22505);
or U22969 (N_22969,N_22753,N_22759);
and U22970 (N_22970,N_22703,N_22746);
xnor U22971 (N_22971,N_22693,N_22721);
and U22972 (N_22972,N_22610,N_22640);
xor U22973 (N_22973,N_22623,N_22516);
xor U22974 (N_22974,N_22781,N_22788);
nand U22975 (N_22975,N_22598,N_22612);
nand U22976 (N_22976,N_22550,N_22686);
nand U22977 (N_22977,N_22770,N_22537);
nand U22978 (N_22978,N_22726,N_22603);
and U22979 (N_22979,N_22560,N_22692);
or U22980 (N_22980,N_22771,N_22647);
nor U22981 (N_22981,N_22593,N_22669);
nand U22982 (N_22982,N_22509,N_22734);
nor U22983 (N_22983,N_22702,N_22562);
or U22984 (N_22984,N_22683,N_22776);
xnor U22985 (N_22985,N_22611,N_22790);
nor U22986 (N_22986,N_22698,N_22500);
nor U22987 (N_22987,N_22550,N_22504);
xor U22988 (N_22988,N_22573,N_22758);
nor U22989 (N_22989,N_22575,N_22559);
nand U22990 (N_22990,N_22634,N_22594);
nand U22991 (N_22991,N_22530,N_22599);
nor U22992 (N_22992,N_22681,N_22509);
nor U22993 (N_22993,N_22631,N_22754);
and U22994 (N_22994,N_22700,N_22724);
xor U22995 (N_22995,N_22649,N_22715);
xnor U22996 (N_22996,N_22715,N_22521);
or U22997 (N_22997,N_22745,N_22671);
and U22998 (N_22998,N_22636,N_22510);
and U22999 (N_22999,N_22620,N_22625);
nor U23000 (N_23000,N_22768,N_22627);
nor U23001 (N_23001,N_22528,N_22542);
and U23002 (N_23002,N_22556,N_22523);
nand U23003 (N_23003,N_22763,N_22718);
nand U23004 (N_23004,N_22739,N_22525);
or U23005 (N_23005,N_22749,N_22507);
and U23006 (N_23006,N_22547,N_22667);
xnor U23007 (N_23007,N_22593,N_22646);
nand U23008 (N_23008,N_22517,N_22791);
xor U23009 (N_23009,N_22518,N_22597);
nor U23010 (N_23010,N_22738,N_22555);
and U23011 (N_23011,N_22604,N_22665);
nor U23012 (N_23012,N_22564,N_22726);
or U23013 (N_23013,N_22766,N_22705);
nand U23014 (N_23014,N_22719,N_22687);
nand U23015 (N_23015,N_22635,N_22610);
nor U23016 (N_23016,N_22699,N_22570);
xnor U23017 (N_23017,N_22539,N_22517);
xor U23018 (N_23018,N_22525,N_22600);
nand U23019 (N_23019,N_22576,N_22701);
xor U23020 (N_23020,N_22594,N_22674);
and U23021 (N_23021,N_22675,N_22561);
nor U23022 (N_23022,N_22697,N_22531);
nor U23023 (N_23023,N_22504,N_22542);
and U23024 (N_23024,N_22605,N_22747);
nor U23025 (N_23025,N_22596,N_22548);
nand U23026 (N_23026,N_22665,N_22753);
and U23027 (N_23027,N_22527,N_22790);
nor U23028 (N_23028,N_22513,N_22716);
and U23029 (N_23029,N_22584,N_22714);
nand U23030 (N_23030,N_22750,N_22653);
nor U23031 (N_23031,N_22673,N_22797);
xnor U23032 (N_23032,N_22579,N_22604);
nor U23033 (N_23033,N_22714,N_22683);
nor U23034 (N_23034,N_22656,N_22538);
nor U23035 (N_23035,N_22694,N_22647);
nor U23036 (N_23036,N_22684,N_22527);
xnor U23037 (N_23037,N_22767,N_22660);
xnor U23038 (N_23038,N_22615,N_22691);
and U23039 (N_23039,N_22727,N_22770);
or U23040 (N_23040,N_22767,N_22699);
xnor U23041 (N_23041,N_22740,N_22728);
xor U23042 (N_23042,N_22603,N_22757);
or U23043 (N_23043,N_22564,N_22713);
nand U23044 (N_23044,N_22527,N_22619);
and U23045 (N_23045,N_22727,N_22504);
nand U23046 (N_23046,N_22796,N_22542);
nand U23047 (N_23047,N_22751,N_22730);
or U23048 (N_23048,N_22713,N_22514);
and U23049 (N_23049,N_22658,N_22734);
or U23050 (N_23050,N_22546,N_22794);
or U23051 (N_23051,N_22738,N_22544);
nand U23052 (N_23052,N_22621,N_22614);
nand U23053 (N_23053,N_22730,N_22595);
nor U23054 (N_23054,N_22746,N_22708);
or U23055 (N_23055,N_22761,N_22630);
xnor U23056 (N_23056,N_22767,N_22531);
xnor U23057 (N_23057,N_22710,N_22675);
or U23058 (N_23058,N_22672,N_22633);
and U23059 (N_23059,N_22678,N_22748);
nand U23060 (N_23060,N_22617,N_22648);
xnor U23061 (N_23061,N_22518,N_22708);
and U23062 (N_23062,N_22652,N_22639);
or U23063 (N_23063,N_22794,N_22703);
and U23064 (N_23064,N_22627,N_22761);
and U23065 (N_23065,N_22610,N_22543);
nor U23066 (N_23066,N_22644,N_22707);
and U23067 (N_23067,N_22543,N_22667);
xor U23068 (N_23068,N_22545,N_22557);
nor U23069 (N_23069,N_22749,N_22758);
or U23070 (N_23070,N_22603,N_22700);
and U23071 (N_23071,N_22794,N_22671);
xnor U23072 (N_23072,N_22569,N_22533);
nand U23073 (N_23073,N_22566,N_22725);
xor U23074 (N_23074,N_22688,N_22755);
xor U23075 (N_23075,N_22643,N_22550);
xor U23076 (N_23076,N_22525,N_22591);
nand U23077 (N_23077,N_22648,N_22552);
and U23078 (N_23078,N_22562,N_22662);
nand U23079 (N_23079,N_22665,N_22662);
or U23080 (N_23080,N_22693,N_22513);
and U23081 (N_23081,N_22771,N_22673);
or U23082 (N_23082,N_22570,N_22775);
nor U23083 (N_23083,N_22737,N_22710);
or U23084 (N_23084,N_22508,N_22743);
nor U23085 (N_23085,N_22611,N_22799);
or U23086 (N_23086,N_22584,N_22705);
and U23087 (N_23087,N_22508,N_22589);
or U23088 (N_23088,N_22740,N_22673);
and U23089 (N_23089,N_22589,N_22623);
and U23090 (N_23090,N_22767,N_22562);
nor U23091 (N_23091,N_22784,N_22750);
or U23092 (N_23092,N_22615,N_22522);
xor U23093 (N_23093,N_22764,N_22606);
xor U23094 (N_23094,N_22773,N_22721);
or U23095 (N_23095,N_22641,N_22796);
xnor U23096 (N_23096,N_22544,N_22790);
or U23097 (N_23097,N_22529,N_22639);
or U23098 (N_23098,N_22761,N_22724);
nor U23099 (N_23099,N_22679,N_22729);
nand U23100 (N_23100,N_22907,N_22849);
nand U23101 (N_23101,N_22940,N_22846);
and U23102 (N_23102,N_22897,N_22876);
xor U23103 (N_23103,N_22821,N_22951);
nor U23104 (N_23104,N_22893,N_22898);
xor U23105 (N_23105,N_22874,N_22807);
or U23106 (N_23106,N_23035,N_23004);
nand U23107 (N_23107,N_23059,N_22931);
nand U23108 (N_23108,N_22946,N_23036);
nor U23109 (N_23109,N_22803,N_22922);
or U23110 (N_23110,N_22935,N_22861);
and U23111 (N_23111,N_22853,N_22947);
nor U23112 (N_23112,N_22965,N_22886);
nand U23113 (N_23113,N_23097,N_22912);
or U23114 (N_23114,N_22975,N_23039);
xor U23115 (N_23115,N_23010,N_22904);
nor U23116 (N_23116,N_22905,N_23012);
nor U23117 (N_23117,N_22958,N_22819);
nor U23118 (N_23118,N_22945,N_22890);
or U23119 (N_23119,N_22923,N_23021);
and U23120 (N_23120,N_22805,N_23098);
and U23121 (N_23121,N_22824,N_22987);
and U23122 (N_23122,N_23075,N_22869);
and U23123 (N_23123,N_22909,N_22857);
or U23124 (N_23124,N_22867,N_23083);
xnor U23125 (N_23125,N_23006,N_22955);
nand U23126 (N_23126,N_23040,N_22970);
and U23127 (N_23127,N_22942,N_22903);
and U23128 (N_23128,N_23063,N_23018);
or U23129 (N_23129,N_22833,N_22981);
nor U23130 (N_23130,N_23064,N_22982);
and U23131 (N_23131,N_22873,N_23081);
nor U23132 (N_23132,N_23053,N_22936);
nand U23133 (N_23133,N_23046,N_22915);
and U23134 (N_23134,N_22832,N_22875);
and U23135 (N_23135,N_22804,N_23090);
or U23136 (N_23136,N_22837,N_22968);
xor U23137 (N_23137,N_23099,N_23043);
nand U23138 (N_23138,N_22925,N_23034);
or U23139 (N_23139,N_23089,N_23091);
and U23140 (N_23140,N_23057,N_22825);
nand U23141 (N_23141,N_22924,N_22842);
nor U23142 (N_23142,N_22887,N_23054);
nand U23143 (N_23143,N_23001,N_22813);
nand U23144 (N_23144,N_22989,N_22995);
nand U23145 (N_23145,N_23029,N_22834);
xnor U23146 (N_23146,N_23068,N_23028);
nand U23147 (N_23147,N_23062,N_22892);
or U23148 (N_23148,N_22938,N_22812);
xnor U23149 (N_23149,N_23008,N_22950);
and U23150 (N_23150,N_22883,N_23072);
and U23151 (N_23151,N_22944,N_22964);
and U23152 (N_23152,N_22919,N_22838);
xor U23153 (N_23153,N_23024,N_23071);
xnor U23154 (N_23154,N_22872,N_23014);
xnor U23155 (N_23155,N_22854,N_23019);
and U23156 (N_23156,N_23041,N_22961);
nor U23157 (N_23157,N_23045,N_23076);
or U23158 (N_23158,N_23070,N_23074);
and U23159 (N_23159,N_22863,N_23047);
xor U23160 (N_23160,N_22865,N_23022);
nor U23161 (N_23161,N_22941,N_22934);
or U23162 (N_23162,N_22808,N_22843);
or U23163 (N_23163,N_22827,N_22848);
nand U23164 (N_23164,N_22847,N_22957);
nor U23165 (N_23165,N_22993,N_23007);
nand U23166 (N_23166,N_22976,N_22966);
xor U23167 (N_23167,N_22878,N_22962);
xnor U23168 (N_23168,N_22800,N_22841);
nor U23169 (N_23169,N_23017,N_22967);
xnor U23170 (N_23170,N_22990,N_23005);
nand U23171 (N_23171,N_22999,N_22918);
xnor U23172 (N_23172,N_23026,N_23082);
or U23173 (N_23173,N_22927,N_22933);
nand U23174 (N_23174,N_23000,N_22906);
and U23175 (N_23175,N_23052,N_22953);
nor U23176 (N_23176,N_22911,N_22879);
nor U23177 (N_23177,N_22992,N_23080);
nand U23178 (N_23178,N_22851,N_22984);
and U23179 (N_23179,N_22889,N_23092);
or U23180 (N_23180,N_22895,N_23042);
and U23181 (N_23181,N_22877,N_22835);
nand U23182 (N_23182,N_22963,N_22818);
nand U23183 (N_23183,N_22926,N_22985);
and U23184 (N_23184,N_22900,N_23079);
nor U23185 (N_23185,N_22928,N_22932);
and U23186 (N_23186,N_23031,N_22952);
or U23187 (N_23187,N_22994,N_22913);
and U23188 (N_23188,N_22917,N_23038);
xor U23189 (N_23189,N_23050,N_22814);
nor U23190 (N_23190,N_22839,N_22826);
or U23191 (N_23191,N_22974,N_22870);
and U23192 (N_23192,N_22823,N_22979);
nor U23193 (N_23193,N_22820,N_23049);
nand U23194 (N_23194,N_23066,N_22973);
or U23195 (N_23195,N_23065,N_22810);
or U23196 (N_23196,N_22891,N_22860);
nor U23197 (N_23197,N_22980,N_23093);
nand U23198 (N_23198,N_22996,N_22971);
and U23199 (N_23199,N_23055,N_22831);
nand U23200 (N_23200,N_22809,N_23061);
xor U23201 (N_23201,N_23073,N_22956);
xnor U23202 (N_23202,N_23044,N_22977);
or U23203 (N_23203,N_22850,N_22828);
nand U23204 (N_23204,N_22859,N_23048);
and U23205 (N_23205,N_22840,N_22845);
xnor U23206 (N_23206,N_22983,N_23032);
xor U23207 (N_23207,N_23051,N_22855);
and U23208 (N_23208,N_22930,N_22836);
and U23209 (N_23209,N_22988,N_22885);
nor U23210 (N_23210,N_22920,N_22829);
nand U23211 (N_23211,N_22868,N_22949);
nand U23212 (N_23212,N_23096,N_22908);
xor U23213 (N_23213,N_22902,N_22862);
and U23214 (N_23214,N_23056,N_22815);
nor U23215 (N_23215,N_22954,N_22806);
or U23216 (N_23216,N_22882,N_23033);
xnor U23217 (N_23217,N_22929,N_22884);
or U23218 (N_23218,N_23094,N_23002);
nand U23219 (N_23219,N_22960,N_22972);
nand U23220 (N_23220,N_22856,N_23058);
xnor U23221 (N_23221,N_22959,N_22852);
nor U23222 (N_23222,N_22830,N_22801);
nand U23223 (N_23223,N_23095,N_23016);
xnor U23224 (N_23224,N_22986,N_22866);
and U23225 (N_23225,N_22914,N_22943);
and U23226 (N_23226,N_23087,N_22948);
and U23227 (N_23227,N_22916,N_22858);
nor U23228 (N_23228,N_22997,N_22816);
nor U23229 (N_23229,N_22817,N_22888);
and U23230 (N_23230,N_22921,N_23084);
xnor U23231 (N_23231,N_23003,N_22871);
nor U23232 (N_23232,N_23030,N_22969);
or U23233 (N_23233,N_23015,N_22844);
nand U23234 (N_23234,N_23025,N_22910);
nand U23235 (N_23235,N_22978,N_23037);
nor U23236 (N_23236,N_23009,N_23013);
or U23237 (N_23237,N_23027,N_22864);
nand U23238 (N_23238,N_23020,N_22939);
nand U23239 (N_23239,N_23011,N_22937);
and U23240 (N_23240,N_23077,N_23086);
nor U23241 (N_23241,N_22896,N_22880);
nand U23242 (N_23242,N_22822,N_23069);
and U23243 (N_23243,N_23088,N_22901);
nor U23244 (N_23244,N_23085,N_23078);
or U23245 (N_23245,N_22881,N_22894);
xor U23246 (N_23246,N_23023,N_22991);
and U23247 (N_23247,N_22899,N_22811);
nor U23248 (N_23248,N_22998,N_23060);
and U23249 (N_23249,N_23067,N_22802);
xnor U23250 (N_23250,N_22861,N_23013);
nor U23251 (N_23251,N_22989,N_22870);
and U23252 (N_23252,N_23075,N_22984);
nor U23253 (N_23253,N_22929,N_23048);
xor U23254 (N_23254,N_23017,N_22976);
and U23255 (N_23255,N_22922,N_22827);
xnor U23256 (N_23256,N_23024,N_22877);
nor U23257 (N_23257,N_22862,N_22803);
or U23258 (N_23258,N_22903,N_22862);
nand U23259 (N_23259,N_22984,N_22918);
xnor U23260 (N_23260,N_22937,N_22896);
and U23261 (N_23261,N_23011,N_22909);
xor U23262 (N_23262,N_22821,N_23095);
xnor U23263 (N_23263,N_22815,N_22919);
or U23264 (N_23264,N_22862,N_23008);
nand U23265 (N_23265,N_22929,N_23032);
nand U23266 (N_23266,N_22816,N_23035);
and U23267 (N_23267,N_23029,N_23027);
or U23268 (N_23268,N_22905,N_22812);
nor U23269 (N_23269,N_23035,N_23016);
and U23270 (N_23270,N_22835,N_23049);
or U23271 (N_23271,N_23088,N_22958);
and U23272 (N_23272,N_22838,N_23075);
nand U23273 (N_23273,N_22857,N_22933);
or U23274 (N_23274,N_22824,N_22931);
or U23275 (N_23275,N_22910,N_22923);
nand U23276 (N_23276,N_22996,N_23040);
xnor U23277 (N_23277,N_23075,N_23018);
nand U23278 (N_23278,N_22950,N_22934);
and U23279 (N_23279,N_22987,N_22913);
and U23280 (N_23280,N_22957,N_22811);
nor U23281 (N_23281,N_22880,N_23066);
or U23282 (N_23282,N_23075,N_22902);
nand U23283 (N_23283,N_22874,N_23019);
or U23284 (N_23284,N_22973,N_22971);
xnor U23285 (N_23285,N_23020,N_23019);
nor U23286 (N_23286,N_22861,N_22991);
nand U23287 (N_23287,N_22818,N_22804);
and U23288 (N_23288,N_23047,N_23011);
nand U23289 (N_23289,N_22827,N_23099);
nand U23290 (N_23290,N_22839,N_22904);
nor U23291 (N_23291,N_22919,N_22932);
nand U23292 (N_23292,N_22870,N_22918);
and U23293 (N_23293,N_22858,N_23051);
xor U23294 (N_23294,N_22808,N_23082);
nor U23295 (N_23295,N_23077,N_23032);
nand U23296 (N_23296,N_23061,N_22991);
xnor U23297 (N_23297,N_23063,N_22936);
nor U23298 (N_23298,N_22889,N_22985);
or U23299 (N_23299,N_23016,N_22885);
or U23300 (N_23300,N_22984,N_22966);
and U23301 (N_23301,N_22821,N_22841);
nand U23302 (N_23302,N_22819,N_22817);
and U23303 (N_23303,N_22811,N_23085);
and U23304 (N_23304,N_23055,N_22893);
and U23305 (N_23305,N_23058,N_22976);
or U23306 (N_23306,N_22833,N_22818);
nand U23307 (N_23307,N_22959,N_23052);
nand U23308 (N_23308,N_22800,N_23066);
and U23309 (N_23309,N_22818,N_22889);
nor U23310 (N_23310,N_23055,N_22947);
and U23311 (N_23311,N_23021,N_22955);
nor U23312 (N_23312,N_23020,N_22977);
nor U23313 (N_23313,N_22807,N_23087);
nand U23314 (N_23314,N_22914,N_22863);
or U23315 (N_23315,N_22904,N_22957);
nand U23316 (N_23316,N_23065,N_22816);
or U23317 (N_23317,N_22962,N_22921);
xnor U23318 (N_23318,N_22805,N_23088);
and U23319 (N_23319,N_23038,N_22817);
xor U23320 (N_23320,N_23032,N_22998);
nand U23321 (N_23321,N_22940,N_22871);
nor U23322 (N_23322,N_22904,N_23048);
or U23323 (N_23323,N_23052,N_22971);
nand U23324 (N_23324,N_23056,N_22999);
and U23325 (N_23325,N_22822,N_23018);
xnor U23326 (N_23326,N_22954,N_22953);
nand U23327 (N_23327,N_22880,N_22988);
nand U23328 (N_23328,N_23015,N_23085);
nor U23329 (N_23329,N_22895,N_22901);
xnor U23330 (N_23330,N_23059,N_22942);
xnor U23331 (N_23331,N_23049,N_22890);
nor U23332 (N_23332,N_23036,N_22969);
or U23333 (N_23333,N_23062,N_23072);
nand U23334 (N_23334,N_22921,N_23059);
and U23335 (N_23335,N_22892,N_22803);
nand U23336 (N_23336,N_23005,N_22838);
xor U23337 (N_23337,N_22902,N_22828);
and U23338 (N_23338,N_22983,N_22827);
nor U23339 (N_23339,N_22845,N_23054);
nand U23340 (N_23340,N_22923,N_23032);
or U23341 (N_23341,N_23049,N_23097);
nor U23342 (N_23342,N_23073,N_23066);
and U23343 (N_23343,N_22933,N_22920);
or U23344 (N_23344,N_22966,N_23034);
or U23345 (N_23345,N_23020,N_23038);
and U23346 (N_23346,N_23072,N_22925);
nor U23347 (N_23347,N_22873,N_22998);
xor U23348 (N_23348,N_23000,N_23029);
xnor U23349 (N_23349,N_23074,N_23006);
or U23350 (N_23350,N_22817,N_23035);
or U23351 (N_23351,N_22944,N_22826);
nand U23352 (N_23352,N_22888,N_22983);
or U23353 (N_23353,N_22863,N_22842);
or U23354 (N_23354,N_22851,N_23017);
xnor U23355 (N_23355,N_22889,N_22951);
and U23356 (N_23356,N_22825,N_22850);
and U23357 (N_23357,N_22943,N_22966);
xor U23358 (N_23358,N_22922,N_22943);
or U23359 (N_23359,N_23015,N_23060);
nor U23360 (N_23360,N_22937,N_23043);
and U23361 (N_23361,N_22969,N_23009);
or U23362 (N_23362,N_22875,N_23093);
or U23363 (N_23363,N_22881,N_22860);
or U23364 (N_23364,N_22848,N_23056);
and U23365 (N_23365,N_22902,N_22941);
xor U23366 (N_23366,N_22996,N_22885);
and U23367 (N_23367,N_23009,N_23089);
nand U23368 (N_23368,N_22962,N_23045);
and U23369 (N_23369,N_22971,N_22801);
and U23370 (N_23370,N_22882,N_23088);
nor U23371 (N_23371,N_23079,N_22844);
nand U23372 (N_23372,N_22986,N_23019);
nand U23373 (N_23373,N_22882,N_22986);
or U23374 (N_23374,N_22832,N_23045);
xor U23375 (N_23375,N_22984,N_23077);
or U23376 (N_23376,N_22963,N_22875);
or U23377 (N_23377,N_23047,N_22929);
nand U23378 (N_23378,N_23078,N_22910);
and U23379 (N_23379,N_22841,N_22902);
nor U23380 (N_23380,N_23087,N_22932);
and U23381 (N_23381,N_22986,N_22822);
nor U23382 (N_23382,N_23025,N_22979);
nand U23383 (N_23383,N_23060,N_22881);
nand U23384 (N_23384,N_23035,N_23067);
or U23385 (N_23385,N_22886,N_22890);
nand U23386 (N_23386,N_22922,N_22807);
or U23387 (N_23387,N_22847,N_22828);
xor U23388 (N_23388,N_23049,N_22806);
or U23389 (N_23389,N_22895,N_22950);
nor U23390 (N_23390,N_22832,N_22840);
xor U23391 (N_23391,N_22966,N_23082);
nor U23392 (N_23392,N_22954,N_22906);
xnor U23393 (N_23393,N_23048,N_22989);
nor U23394 (N_23394,N_23036,N_23078);
and U23395 (N_23395,N_22801,N_23016);
nand U23396 (N_23396,N_22889,N_22918);
and U23397 (N_23397,N_23009,N_22880);
nand U23398 (N_23398,N_22943,N_23083);
or U23399 (N_23399,N_23010,N_22824);
nand U23400 (N_23400,N_23258,N_23121);
or U23401 (N_23401,N_23145,N_23376);
nor U23402 (N_23402,N_23396,N_23227);
nand U23403 (N_23403,N_23374,N_23228);
and U23404 (N_23404,N_23154,N_23256);
xnor U23405 (N_23405,N_23365,N_23157);
xnor U23406 (N_23406,N_23229,N_23272);
nor U23407 (N_23407,N_23250,N_23137);
nor U23408 (N_23408,N_23142,N_23378);
xor U23409 (N_23409,N_23398,N_23202);
and U23410 (N_23410,N_23138,N_23291);
nor U23411 (N_23411,N_23271,N_23148);
nor U23412 (N_23412,N_23348,N_23215);
nor U23413 (N_23413,N_23355,N_23340);
xor U23414 (N_23414,N_23139,N_23356);
or U23415 (N_23415,N_23130,N_23373);
and U23416 (N_23416,N_23399,N_23395);
xnor U23417 (N_23417,N_23380,N_23204);
and U23418 (N_23418,N_23205,N_23175);
or U23419 (N_23419,N_23113,N_23331);
nand U23420 (N_23420,N_23252,N_23102);
and U23421 (N_23421,N_23296,N_23264);
or U23422 (N_23422,N_23387,N_23134);
nor U23423 (N_23423,N_23289,N_23276);
xor U23424 (N_23424,N_23372,N_23176);
nor U23425 (N_23425,N_23318,N_23159);
nor U23426 (N_23426,N_23201,N_23337);
nor U23427 (N_23427,N_23251,N_23320);
xor U23428 (N_23428,N_23287,N_23300);
and U23429 (N_23429,N_23120,N_23327);
nor U23430 (N_23430,N_23246,N_23254);
xor U23431 (N_23431,N_23126,N_23194);
and U23432 (N_23432,N_23129,N_23248);
and U23433 (N_23433,N_23312,N_23325);
nor U23434 (N_23434,N_23141,N_23110);
xor U23435 (N_23435,N_23104,N_23219);
xnor U23436 (N_23436,N_23156,N_23132);
nand U23437 (N_23437,N_23239,N_23161);
or U23438 (N_23438,N_23107,N_23283);
and U23439 (N_23439,N_23238,N_23209);
nor U23440 (N_23440,N_23343,N_23332);
xnor U23441 (N_23441,N_23358,N_23370);
nor U23442 (N_23442,N_23278,N_23269);
nand U23443 (N_23443,N_23203,N_23393);
or U23444 (N_23444,N_23367,N_23218);
nand U23445 (N_23445,N_23379,N_23207);
nand U23446 (N_23446,N_23108,N_23324);
nand U23447 (N_23447,N_23143,N_23124);
nor U23448 (N_23448,N_23242,N_23191);
nand U23449 (N_23449,N_23232,N_23273);
nor U23450 (N_23450,N_23210,N_23304);
and U23451 (N_23451,N_23371,N_23383);
xor U23452 (N_23452,N_23182,N_23294);
nor U23453 (N_23453,N_23266,N_23341);
xor U23454 (N_23454,N_23275,N_23106);
or U23455 (N_23455,N_23316,N_23184);
xnor U23456 (N_23456,N_23185,N_23263);
or U23457 (N_23457,N_23359,N_23150);
xnor U23458 (N_23458,N_23149,N_23153);
or U23459 (N_23459,N_23206,N_23174);
nand U23460 (N_23460,N_23315,N_23101);
and U23461 (N_23461,N_23155,N_23178);
xnor U23462 (N_23462,N_23310,N_23303);
or U23463 (N_23463,N_23330,N_23375);
nor U23464 (N_23464,N_23190,N_23173);
xor U23465 (N_23465,N_23119,N_23249);
xor U23466 (N_23466,N_23127,N_23196);
xor U23467 (N_23467,N_23165,N_23241);
nand U23468 (N_23468,N_23200,N_23195);
nor U23469 (N_23469,N_23240,N_23347);
xnor U23470 (N_23470,N_23122,N_23117);
nand U23471 (N_23471,N_23225,N_23255);
nor U23472 (N_23472,N_23169,N_23322);
nor U23473 (N_23473,N_23279,N_23236);
xnor U23474 (N_23474,N_23197,N_23319);
nor U23475 (N_23475,N_23345,N_23354);
nor U23476 (N_23476,N_23147,N_23268);
or U23477 (N_23477,N_23260,N_23166);
or U23478 (N_23478,N_23285,N_23144);
nand U23479 (N_23479,N_23362,N_23351);
nor U23480 (N_23480,N_23237,N_23188);
nand U23481 (N_23481,N_23234,N_23336);
and U23482 (N_23482,N_23381,N_23140);
or U23483 (N_23483,N_23257,N_23288);
and U23484 (N_23484,N_23103,N_23160);
nor U23485 (N_23485,N_23286,N_23189);
nand U23486 (N_23486,N_23226,N_23180);
or U23487 (N_23487,N_23244,N_23222);
nand U23488 (N_23488,N_23172,N_23163);
xnor U23489 (N_23489,N_23211,N_23323);
and U23490 (N_23490,N_23193,N_23298);
and U23491 (N_23491,N_23162,N_23235);
and U23492 (N_23492,N_23259,N_23183);
nand U23493 (N_23493,N_23302,N_23192);
and U23494 (N_23494,N_23357,N_23293);
nor U23495 (N_23495,N_23146,N_23136);
nand U23496 (N_23496,N_23301,N_23133);
or U23497 (N_23497,N_23350,N_23353);
nand U23498 (N_23498,N_23306,N_23295);
nand U23499 (N_23499,N_23168,N_23392);
nor U23500 (N_23500,N_23212,N_23181);
and U23501 (N_23501,N_23281,N_23167);
or U23502 (N_23502,N_23164,N_23224);
and U23503 (N_23503,N_23282,N_23280);
nor U23504 (N_23504,N_23368,N_23313);
nand U23505 (N_23505,N_23217,N_23290);
xnor U23506 (N_23506,N_23261,N_23344);
or U23507 (N_23507,N_23369,N_23389);
and U23508 (N_23508,N_23270,N_23352);
xnor U23509 (N_23509,N_23307,N_23216);
nand U23510 (N_23510,N_23297,N_23333);
nor U23511 (N_23511,N_23314,N_23223);
nor U23512 (N_23512,N_23360,N_23221);
nand U23513 (N_23513,N_23179,N_23123);
and U23514 (N_23514,N_23233,N_23186);
nand U23515 (N_23515,N_23317,N_23334);
xor U23516 (N_23516,N_23309,N_23247);
xnor U23517 (N_23517,N_23265,N_23231);
xnor U23518 (N_23518,N_23349,N_23118);
nor U23519 (N_23519,N_23171,N_23384);
nor U23520 (N_23520,N_23151,N_23397);
nor U23521 (N_23521,N_23245,N_23363);
and U23522 (N_23522,N_23335,N_23338);
and U23523 (N_23523,N_23326,N_23388);
nor U23524 (N_23524,N_23220,N_23274);
and U23525 (N_23525,N_23131,N_23329);
nor U23526 (N_23526,N_23115,N_23152);
and U23527 (N_23527,N_23299,N_23214);
nand U23528 (N_23528,N_23385,N_23361);
nor U23529 (N_23529,N_23377,N_23390);
nand U23530 (N_23530,N_23328,N_23177);
xor U23531 (N_23531,N_23230,N_23109);
xnor U23532 (N_23532,N_23199,N_23125);
and U23533 (N_23533,N_23284,N_23277);
nand U23534 (N_23534,N_23111,N_23346);
nor U23535 (N_23535,N_23170,N_23135);
nand U23536 (N_23536,N_23100,N_23311);
nor U23537 (N_23537,N_23342,N_23116);
or U23538 (N_23538,N_23243,N_23292);
nor U23539 (N_23539,N_23253,N_23386);
and U23540 (N_23540,N_23308,N_23187);
and U23541 (N_23541,N_23198,N_23208);
or U23542 (N_23542,N_23158,N_23366);
nand U23543 (N_23543,N_23305,N_23114);
and U23544 (N_23544,N_23267,N_23391);
nand U23545 (N_23545,N_23262,N_23394);
xnor U23546 (N_23546,N_23105,N_23112);
nand U23547 (N_23547,N_23321,N_23213);
and U23548 (N_23548,N_23364,N_23128);
and U23549 (N_23549,N_23382,N_23339);
nor U23550 (N_23550,N_23177,N_23311);
nor U23551 (N_23551,N_23302,N_23201);
or U23552 (N_23552,N_23103,N_23398);
nor U23553 (N_23553,N_23298,N_23396);
xor U23554 (N_23554,N_23205,N_23133);
and U23555 (N_23555,N_23117,N_23281);
nor U23556 (N_23556,N_23286,N_23298);
nor U23557 (N_23557,N_23136,N_23211);
nand U23558 (N_23558,N_23392,N_23380);
nand U23559 (N_23559,N_23319,N_23215);
and U23560 (N_23560,N_23169,N_23265);
or U23561 (N_23561,N_23141,N_23281);
xor U23562 (N_23562,N_23287,N_23137);
nor U23563 (N_23563,N_23279,N_23250);
nand U23564 (N_23564,N_23276,N_23284);
and U23565 (N_23565,N_23391,N_23146);
nor U23566 (N_23566,N_23374,N_23147);
xor U23567 (N_23567,N_23204,N_23111);
and U23568 (N_23568,N_23319,N_23395);
and U23569 (N_23569,N_23350,N_23329);
nor U23570 (N_23570,N_23263,N_23368);
or U23571 (N_23571,N_23322,N_23376);
and U23572 (N_23572,N_23143,N_23139);
xnor U23573 (N_23573,N_23232,N_23190);
nor U23574 (N_23574,N_23119,N_23262);
nor U23575 (N_23575,N_23178,N_23247);
or U23576 (N_23576,N_23363,N_23103);
xor U23577 (N_23577,N_23213,N_23124);
xor U23578 (N_23578,N_23370,N_23253);
nor U23579 (N_23579,N_23147,N_23378);
or U23580 (N_23580,N_23121,N_23389);
xnor U23581 (N_23581,N_23186,N_23242);
nand U23582 (N_23582,N_23292,N_23106);
nor U23583 (N_23583,N_23122,N_23174);
or U23584 (N_23584,N_23376,N_23281);
xnor U23585 (N_23585,N_23187,N_23246);
or U23586 (N_23586,N_23277,N_23352);
nand U23587 (N_23587,N_23383,N_23376);
nor U23588 (N_23588,N_23379,N_23351);
nor U23589 (N_23589,N_23101,N_23213);
xor U23590 (N_23590,N_23207,N_23163);
and U23591 (N_23591,N_23128,N_23233);
and U23592 (N_23592,N_23382,N_23146);
nand U23593 (N_23593,N_23330,N_23382);
xor U23594 (N_23594,N_23324,N_23200);
nand U23595 (N_23595,N_23210,N_23363);
and U23596 (N_23596,N_23340,N_23106);
nor U23597 (N_23597,N_23365,N_23192);
and U23598 (N_23598,N_23284,N_23282);
xnor U23599 (N_23599,N_23332,N_23369);
and U23600 (N_23600,N_23130,N_23325);
nand U23601 (N_23601,N_23209,N_23316);
and U23602 (N_23602,N_23399,N_23248);
and U23603 (N_23603,N_23252,N_23135);
xor U23604 (N_23604,N_23328,N_23301);
nor U23605 (N_23605,N_23348,N_23163);
nor U23606 (N_23606,N_23181,N_23148);
and U23607 (N_23607,N_23344,N_23248);
or U23608 (N_23608,N_23321,N_23123);
nor U23609 (N_23609,N_23395,N_23176);
and U23610 (N_23610,N_23155,N_23337);
and U23611 (N_23611,N_23378,N_23213);
and U23612 (N_23612,N_23250,N_23213);
or U23613 (N_23613,N_23289,N_23341);
and U23614 (N_23614,N_23122,N_23389);
xor U23615 (N_23615,N_23228,N_23348);
and U23616 (N_23616,N_23304,N_23331);
nor U23617 (N_23617,N_23231,N_23250);
or U23618 (N_23618,N_23182,N_23201);
and U23619 (N_23619,N_23374,N_23341);
nand U23620 (N_23620,N_23163,N_23139);
or U23621 (N_23621,N_23301,N_23371);
or U23622 (N_23622,N_23179,N_23261);
nor U23623 (N_23623,N_23271,N_23206);
nand U23624 (N_23624,N_23163,N_23166);
and U23625 (N_23625,N_23281,N_23187);
or U23626 (N_23626,N_23331,N_23147);
xor U23627 (N_23627,N_23378,N_23129);
nand U23628 (N_23628,N_23140,N_23289);
and U23629 (N_23629,N_23149,N_23366);
nand U23630 (N_23630,N_23347,N_23260);
xor U23631 (N_23631,N_23109,N_23334);
xnor U23632 (N_23632,N_23275,N_23291);
and U23633 (N_23633,N_23136,N_23366);
or U23634 (N_23634,N_23185,N_23115);
nor U23635 (N_23635,N_23366,N_23221);
xor U23636 (N_23636,N_23382,N_23356);
xnor U23637 (N_23637,N_23108,N_23116);
nand U23638 (N_23638,N_23260,N_23389);
xor U23639 (N_23639,N_23302,N_23233);
xnor U23640 (N_23640,N_23352,N_23283);
nor U23641 (N_23641,N_23166,N_23127);
and U23642 (N_23642,N_23239,N_23219);
nor U23643 (N_23643,N_23222,N_23169);
or U23644 (N_23644,N_23117,N_23227);
xnor U23645 (N_23645,N_23360,N_23225);
xnor U23646 (N_23646,N_23101,N_23189);
nand U23647 (N_23647,N_23241,N_23166);
nor U23648 (N_23648,N_23246,N_23382);
or U23649 (N_23649,N_23246,N_23148);
xnor U23650 (N_23650,N_23341,N_23182);
xnor U23651 (N_23651,N_23296,N_23305);
nor U23652 (N_23652,N_23358,N_23107);
and U23653 (N_23653,N_23117,N_23353);
and U23654 (N_23654,N_23326,N_23186);
nand U23655 (N_23655,N_23250,N_23264);
and U23656 (N_23656,N_23236,N_23296);
nand U23657 (N_23657,N_23326,N_23245);
nor U23658 (N_23658,N_23397,N_23194);
nand U23659 (N_23659,N_23268,N_23200);
or U23660 (N_23660,N_23169,N_23388);
and U23661 (N_23661,N_23324,N_23136);
xnor U23662 (N_23662,N_23362,N_23318);
and U23663 (N_23663,N_23249,N_23283);
nor U23664 (N_23664,N_23174,N_23230);
nand U23665 (N_23665,N_23259,N_23295);
or U23666 (N_23666,N_23300,N_23360);
nor U23667 (N_23667,N_23102,N_23147);
xor U23668 (N_23668,N_23394,N_23320);
and U23669 (N_23669,N_23243,N_23112);
nor U23670 (N_23670,N_23183,N_23263);
nor U23671 (N_23671,N_23294,N_23210);
nand U23672 (N_23672,N_23373,N_23186);
xnor U23673 (N_23673,N_23235,N_23379);
xor U23674 (N_23674,N_23185,N_23330);
xnor U23675 (N_23675,N_23232,N_23107);
xnor U23676 (N_23676,N_23171,N_23272);
nand U23677 (N_23677,N_23356,N_23372);
xor U23678 (N_23678,N_23101,N_23269);
nand U23679 (N_23679,N_23276,N_23222);
nor U23680 (N_23680,N_23183,N_23349);
xor U23681 (N_23681,N_23384,N_23213);
and U23682 (N_23682,N_23287,N_23322);
or U23683 (N_23683,N_23219,N_23361);
or U23684 (N_23684,N_23211,N_23226);
and U23685 (N_23685,N_23183,N_23300);
and U23686 (N_23686,N_23233,N_23348);
nand U23687 (N_23687,N_23251,N_23156);
and U23688 (N_23688,N_23298,N_23381);
nor U23689 (N_23689,N_23149,N_23377);
nand U23690 (N_23690,N_23261,N_23120);
nor U23691 (N_23691,N_23378,N_23319);
nor U23692 (N_23692,N_23280,N_23299);
or U23693 (N_23693,N_23209,N_23307);
xnor U23694 (N_23694,N_23333,N_23374);
nor U23695 (N_23695,N_23123,N_23188);
nand U23696 (N_23696,N_23331,N_23111);
nand U23697 (N_23697,N_23212,N_23253);
nor U23698 (N_23698,N_23322,N_23258);
nor U23699 (N_23699,N_23220,N_23265);
nor U23700 (N_23700,N_23483,N_23575);
nand U23701 (N_23701,N_23657,N_23426);
xor U23702 (N_23702,N_23526,N_23452);
xor U23703 (N_23703,N_23470,N_23551);
xnor U23704 (N_23704,N_23446,N_23695);
and U23705 (N_23705,N_23460,N_23607);
nor U23706 (N_23706,N_23417,N_23490);
or U23707 (N_23707,N_23493,N_23419);
nor U23708 (N_23708,N_23683,N_23504);
or U23709 (N_23709,N_23475,N_23599);
nor U23710 (N_23710,N_23651,N_23619);
or U23711 (N_23711,N_23616,N_23652);
and U23712 (N_23712,N_23517,N_23543);
or U23713 (N_23713,N_23447,N_23502);
nor U23714 (N_23714,N_23429,N_23583);
or U23715 (N_23715,N_23612,N_23615);
xnor U23716 (N_23716,N_23596,N_23643);
nor U23717 (N_23717,N_23510,N_23527);
nand U23718 (N_23718,N_23680,N_23423);
nand U23719 (N_23719,N_23554,N_23529);
nand U23720 (N_23720,N_23610,N_23591);
nor U23721 (N_23721,N_23542,N_23671);
and U23722 (N_23722,N_23560,N_23598);
nor U23723 (N_23723,N_23676,N_23416);
nor U23724 (N_23724,N_23590,N_23477);
and U23725 (N_23725,N_23432,N_23669);
nor U23726 (N_23726,N_23618,N_23660);
nand U23727 (N_23727,N_23459,N_23686);
and U23728 (N_23728,N_23541,N_23521);
or U23729 (N_23729,N_23530,N_23584);
nand U23730 (N_23730,N_23533,N_23454);
xnor U23731 (N_23731,N_23581,N_23649);
nor U23732 (N_23732,N_23573,N_23414);
nor U23733 (N_23733,N_23518,N_23558);
nand U23734 (N_23734,N_23613,N_23571);
nand U23735 (N_23735,N_23539,N_23552);
and U23736 (N_23736,N_23611,N_23609);
xnor U23737 (N_23737,N_23614,N_23544);
and U23738 (N_23738,N_23620,N_23699);
and U23739 (N_23739,N_23630,N_23507);
or U23740 (N_23740,N_23656,N_23640);
nor U23741 (N_23741,N_23650,N_23677);
nand U23742 (N_23742,N_23582,N_23546);
and U23743 (N_23743,N_23678,N_23561);
nor U23744 (N_23744,N_23471,N_23629);
or U23745 (N_23745,N_23566,N_23421);
or U23746 (N_23746,N_23668,N_23628);
or U23747 (N_23747,N_23500,N_23427);
nand U23748 (N_23748,N_23468,N_23523);
nand U23749 (N_23749,N_23684,N_23666);
and U23750 (N_23750,N_23570,N_23675);
and U23751 (N_23751,N_23531,N_23667);
nand U23752 (N_23752,N_23645,N_23519);
nor U23753 (N_23753,N_23633,N_23644);
and U23754 (N_23754,N_23453,N_23430);
nor U23755 (N_23755,N_23679,N_23617);
or U23756 (N_23756,N_23594,N_23457);
nor U23757 (N_23757,N_23685,N_23580);
nor U23758 (N_23758,N_23512,N_23435);
nand U23759 (N_23759,N_23437,N_23442);
or U23760 (N_23760,N_23497,N_23661);
and U23761 (N_23761,N_23511,N_23402);
and U23762 (N_23762,N_23673,N_23444);
or U23763 (N_23763,N_23403,N_23592);
nand U23764 (N_23764,N_23503,N_23588);
xor U23765 (N_23765,N_23597,N_23694);
nor U23766 (N_23766,N_23602,N_23494);
nor U23767 (N_23767,N_23639,N_23476);
xor U23768 (N_23768,N_23627,N_23664);
and U23769 (N_23769,N_23479,N_23522);
nand U23770 (N_23770,N_23491,N_23622);
and U23771 (N_23771,N_23687,N_23557);
xnor U23772 (N_23772,N_23422,N_23410);
and U23773 (N_23773,N_23455,N_23698);
xnor U23774 (N_23774,N_23451,N_23670);
or U23775 (N_23775,N_23545,N_23434);
xor U23776 (N_23776,N_23458,N_23537);
xor U23777 (N_23777,N_23681,N_23450);
and U23778 (N_23778,N_23572,N_23485);
xnor U23779 (N_23779,N_23568,N_23593);
or U23780 (N_23780,N_23654,N_23555);
or U23781 (N_23781,N_23495,N_23632);
nand U23782 (N_23782,N_23589,N_23549);
or U23783 (N_23783,N_23408,N_23578);
and U23784 (N_23784,N_23516,N_23492);
nand U23785 (N_23785,N_23642,N_23534);
nand U23786 (N_23786,N_23436,N_23641);
nand U23787 (N_23787,N_23449,N_23431);
or U23788 (N_23788,N_23506,N_23462);
nand U23789 (N_23789,N_23469,N_23621);
or U23790 (N_23790,N_23562,N_23556);
xor U23791 (N_23791,N_23400,N_23662);
and U23792 (N_23792,N_23484,N_23606);
or U23793 (N_23793,N_23532,N_23463);
nor U23794 (N_23794,N_23472,N_23601);
and U23795 (N_23795,N_23428,N_23579);
xor U23796 (N_23796,N_23646,N_23538);
nand U23797 (N_23797,N_23653,N_23623);
xnor U23798 (N_23798,N_23631,N_23540);
and U23799 (N_23799,N_23647,N_23440);
or U23800 (N_23800,N_23488,N_23505);
nor U23801 (N_23801,N_23663,N_23443);
nand U23802 (N_23802,N_23420,N_23689);
and U23803 (N_23803,N_23515,N_23466);
nand U23804 (N_23804,N_23691,N_23585);
or U23805 (N_23805,N_23567,N_23473);
or U23806 (N_23806,N_23625,N_23425);
nor U23807 (N_23807,N_23482,N_23674);
or U23808 (N_23808,N_23513,N_23587);
and U23809 (N_23809,N_23659,N_23520);
or U23810 (N_23810,N_23595,N_23411);
xor U23811 (N_23811,N_23550,N_23577);
or U23812 (N_23812,N_23547,N_23603);
and U23813 (N_23813,N_23486,N_23478);
xor U23814 (N_23814,N_23480,N_23418);
nand U23815 (N_23815,N_23439,N_23481);
xnor U23816 (N_23816,N_23461,N_23487);
and U23817 (N_23817,N_23524,N_23682);
and U23818 (N_23818,N_23424,N_23665);
xor U23819 (N_23819,N_23658,N_23648);
xnor U23820 (N_23820,N_23514,N_23692);
and U23821 (N_23821,N_23604,N_23636);
or U23822 (N_23822,N_23401,N_23413);
or U23823 (N_23823,N_23407,N_23672);
and U23824 (N_23824,N_23456,N_23489);
xnor U23825 (N_23825,N_23535,N_23528);
and U23826 (N_23826,N_23501,N_23564);
xor U23827 (N_23827,N_23499,N_23608);
or U23828 (N_23828,N_23404,N_23509);
nand U23829 (N_23829,N_23445,N_23496);
xnor U23830 (N_23830,N_23574,N_23525);
xnor U23831 (N_23831,N_23536,N_23576);
and U23832 (N_23832,N_23563,N_23600);
or U23833 (N_23833,N_23548,N_23559);
nor U23834 (N_23834,N_23412,N_23624);
nand U23835 (N_23835,N_23690,N_23438);
xnor U23836 (N_23836,N_23465,N_23474);
nand U23837 (N_23837,N_23441,N_23467);
nor U23838 (N_23838,N_23688,N_23638);
nor U23839 (N_23839,N_23405,N_23565);
xor U23840 (N_23840,N_23569,N_23693);
and U23841 (N_23841,N_23448,N_23655);
or U23842 (N_23842,N_23553,N_23409);
xnor U23843 (N_23843,N_23635,N_23498);
xnor U23844 (N_23844,N_23605,N_23637);
or U23845 (N_23845,N_23433,N_23586);
nor U23846 (N_23846,N_23696,N_23508);
or U23847 (N_23847,N_23415,N_23464);
nor U23848 (N_23848,N_23406,N_23626);
xnor U23849 (N_23849,N_23634,N_23697);
xnor U23850 (N_23850,N_23504,N_23567);
nor U23851 (N_23851,N_23632,N_23536);
and U23852 (N_23852,N_23627,N_23614);
nand U23853 (N_23853,N_23465,N_23660);
nor U23854 (N_23854,N_23473,N_23502);
nor U23855 (N_23855,N_23405,N_23661);
or U23856 (N_23856,N_23589,N_23442);
nand U23857 (N_23857,N_23588,N_23441);
nor U23858 (N_23858,N_23524,N_23564);
nor U23859 (N_23859,N_23549,N_23461);
or U23860 (N_23860,N_23443,N_23581);
nand U23861 (N_23861,N_23519,N_23688);
and U23862 (N_23862,N_23442,N_23401);
or U23863 (N_23863,N_23442,N_23674);
nand U23864 (N_23864,N_23627,N_23484);
nor U23865 (N_23865,N_23441,N_23454);
or U23866 (N_23866,N_23690,N_23409);
or U23867 (N_23867,N_23476,N_23541);
and U23868 (N_23868,N_23576,N_23595);
and U23869 (N_23869,N_23592,N_23446);
or U23870 (N_23870,N_23553,N_23599);
and U23871 (N_23871,N_23572,N_23495);
or U23872 (N_23872,N_23442,N_23634);
xor U23873 (N_23873,N_23494,N_23439);
nand U23874 (N_23874,N_23613,N_23675);
xnor U23875 (N_23875,N_23423,N_23618);
and U23876 (N_23876,N_23667,N_23538);
and U23877 (N_23877,N_23617,N_23511);
xor U23878 (N_23878,N_23427,N_23608);
and U23879 (N_23879,N_23645,N_23683);
or U23880 (N_23880,N_23569,N_23670);
and U23881 (N_23881,N_23516,N_23642);
xor U23882 (N_23882,N_23687,N_23431);
and U23883 (N_23883,N_23486,N_23501);
nand U23884 (N_23884,N_23542,N_23651);
xor U23885 (N_23885,N_23579,N_23612);
nand U23886 (N_23886,N_23607,N_23601);
or U23887 (N_23887,N_23618,N_23506);
and U23888 (N_23888,N_23557,N_23675);
and U23889 (N_23889,N_23668,N_23442);
and U23890 (N_23890,N_23696,N_23472);
nor U23891 (N_23891,N_23661,N_23606);
nand U23892 (N_23892,N_23615,N_23681);
or U23893 (N_23893,N_23555,N_23690);
nand U23894 (N_23894,N_23617,N_23561);
and U23895 (N_23895,N_23456,N_23691);
xor U23896 (N_23896,N_23591,N_23666);
xnor U23897 (N_23897,N_23631,N_23643);
and U23898 (N_23898,N_23596,N_23546);
or U23899 (N_23899,N_23572,N_23539);
or U23900 (N_23900,N_23522,N_23580);
nor U23901 (N_23901,N_23551,N_23456);
and U23902 (N_23902,N_23523,N_23579);
or U23903 (N_23903,N_23455,N_23424);
nand U23904 (N_23904,N_23618,N_23491);
nor U23905 (N_23905,N_23690,N_23596);
or U23906 (N_23906,N_23616,N_23452);
xnor U23907 (N_23907,N_23534,N_23632);
xor U23908 (N_23908,N_23692,N_23472);
nand U23909 (N_23909,N_23537,N_23533);
and U23910 (N_23910,N_23587,N_23585);
nand U23911 (N_23911,N_23620,N_23615);
xor U23912 (N_23912,N_23630,N_23528);
and U23913 (N_23913,N_23559,N_23411);
or U23914 (N_23914,N_23597,N_23490);
nand U23915 (N_23915,N_23612,N_23537);
or U23916 (N_23916,N_23661,N_23434);
or U23917 (N_23917,N_23684,N_23596);
nand U23918 (N_23918,N_23404,N_23624);
and U23919 (N_23919,N_23540,N_23459);
nor U23920 (N_23920,N_23676,N_23630);
and U23921 (N_23921,N_23432,N_23666);
and U23922 (N_23922,N_23637,N_23650);
xnor U23923 (N_23923,N_23563,N_23566);
nor U23924 (N_23924,N_23693,N_23512);
nor U23925 (N_23925,N_23663,N_23575);
and U23926 (N_23926,N_23530,N_23467);
nor U23927 (N_23927,N_23492,N_23439);
or U23928 (N_23928,N_23607,N_23430);
and U23929 (N_23929,N_23500,N_23663);
nand U23930 (N_23930,N_23519,N_23446);
and U23931 (N_23931,N_23618,N_23480);
nand U23932 (N_23932,N_23650,N_23402);
or U23933 (N_23933,N_23696,N_23409);
nor U23934 (N_23934,N_23548,N_23438);
and U23935 (N_23935,N_23413,N_23591);
or U23936 (N_23936,N_23492,N_23628);
nor U23937 (N_23937,N_23426,N_23402);
nor U23938 (N_23938,N_23697,N_23463);
xor U23939 (N_23939,N_23457,N_23513);
and U23940 (N_23940,N_23508,N_23428);
or U23941 (N_23941,N_23464,N_23585);
nand U23942 (N_23942,N_23666,N_23621);
xnor U23943 (N_23943,N_23615,N_23430);
and U23944 (N_23944,N_23602,N_23643);
and U23945 (N_23945,N_23546,N_23424);
or U23946 (N_23946,N_23512,N_23578);
nand U23947 (N_23947,N_23559,N_23524);
or U23948 (N_23948,N_23419,N_23607);
nor U23949 (N_23949,N_23497,N_23653);
or U23950 (N_23950,N_23590,N_23427);
and U23951 (N_23951,N_23568,N_23645);
xor U23952 (N_23952,N_23681,N_23519);
nor U23953 (N_23953,N_23687,N_23420);
xor U23954 (N_23954,N_23470,N_23676);
nand U23955 (N_23955,N_23532,N_23660);
xnor U23956 (N_23956,N_23595,N_23654);
xor U23957 (N_23957,N_23595,N_23566);
xor U23958 (N_23958,N_23578,N_23524);
and U23959 (N_23959,N_23422,N_23678);
nand U23960 (N_23960,N_23602,N_23479);
xor U23961 (N_23961,N_23578,N_23525);
and U23962 (N_23962,N_23657,N_23678);
nor U23963 (N_23963,N_23674,N_23509);
nand U23964 (N_23964,N_23585,N_23589);
nand U23965 (N_23965,N_23512,N_23604);
and U23966 (N_23966,N_23461,N_23612);
xor U23967 (N_23967,N_23456,N_23515);
nand U23968 (N_23968,N_23544,N_23402);
and U23969 (N_23969,N_23547,N_23496);
or U23970 (N_23970,N_23601,N_23677);
nor U23971 (N_23971,N_23441,N_23552);
or U23972 (N_23972,N_23530,N_23677);
nand U23973 (N_23973,N_23516,N_23447);
nor U23974 (N_23974,N_23558,N_23463);
nand U23975 (N_23975,N_23597,N_23616);
and U23976 (N_23976,N_23687,N_23664);
xor U23977 (N_23977,N_23546,N_23695);
and U23978 (N_23978,N_23485,N_23595);
nand U23979 (N_23979,N_23606,N_23607);
or U23980 (N_23980,N_23455,N_23688);
xor U23981 (N_23981,N_23630,N_23561);
nand U23982 (N_23982,N_23542,N_23648);
nand U23983 (N_23983,N_23553,N_23592);
nor U23984 (N_23984,N_23527,N_23676);
xnor U23985 (N_23985,N_23686,N_23650);
and U23986 (N_23986,N_23512,N_23673);
or U23987 (N_23987,N_23558,N_23414);
nand U23988 (N_23988,N_23452,N_23435);
or U23989 (N_23989,N_23654,N_23402);
xor U23990 (N_23990,N_23676,N_23668);
and U23991 (N_23991,N_23410,N_23608);
and U23992 (N_23992,N_23673,N_23621);
xnor U23993 (N_23993,N_23471,N_23676);
and U23994 (N_23994,N_23672,N_23637);
nand U23995 (N_23995,N_23412,N_23625);
nor U23996 (N_23996,N_23474,N_23508);
nand U23997 (N_23997,N_23591,N_23654);
xor U23998 (N_23998,N_23641,N_23655);
nand U23999 (N_23999,N_23696,N_23493);
nand U24000 (N_24000,N_23833,N_23761);
nand U24001 (N_24001,N_23746,N_23965);
nand U24002 (N_24002,N_23997,N_23843);
and U24003 (N_24003,N_23947,N_23803);
nand U24004 (N_24004,N_23981,N_23788);
or U24005 (N_24005,N_23739,N_23767);
xor U24006 (N_24006,N_23921,N_23934);
nor U24007 (N_24007,N_23868,N_23734);
xnor U24008 (N_24008,N_23926,N_23955);
and U24009 (N_24009,N_23718,N_23757);
xor U24010 (N_24010,N_23889,N_23996);
xor U24011 (N_24011,N_23736,N_23800);
nand U24012 (N_24012,N_23875,N_23970);
or U24013 (N_24013,N_23842,N_23922);
and U24014 (N_24014,N_23887,N_23933);
nand U24015 (N_24015,N_23978,N_23785);
or U24016 (N_24016,N_23975,N_23766);
nand U24017 (N_24017,N_23902,N_23863);
nor U24018 (N_24018,N_23764,N_23799);
or U24019 (N_24019,N_23704,N_23879);
or U24020 (N_24020,N_23993,N_23849);
or U24021 (N_24021,N_23814,N_23769);
xnor U24022 (N_24022,N_23885,N_23852);
nor U24023 (N_24023,N_23771,N_23848);
and U24024 (N_24024,N_23983,N_23949);
nand U24025 (N_24025,N_23756,N_23869);
and U24026 (N_24026,N_23721,N_23827);
nor U24027 (N_24027,N_23758,N_23811);
xnor U24028 (N_24028,N_23991,N_23824);
nand U24029 (N_24029,N_23893,N_23715);
or U24030 (N_24030,N_23895,N_23999);
xnor U24031 (N_24031,N_23805,N_23751);
nand U24032 (N_24032,N_23722,N_23915);
and U24033 (N_24033,N_23948,N_23728);
xnor U24034 (N_24034,N_23775,N_23702);
xor U24035 (N_24035,N_23919,N_23851);
xor U24036 (N_24036,N_23931,N_23857);
nor U24037 (N_24037,N_23829,N_23910);
nor U24038 (N_24038,N_23930,N_23813);
nor U24039 (N_24039,N_23765,N_23936);
and U24040 (N_24040,N_23914,N_23943);
nand U24041 (N_24041,N_23841,N_23801);
and U24042 (N_24042,N_23817,N_23872);
xnor U24043 (N_24043,N_23807,N_23752);
nand U24044 (N_24044,N_23952,N_23859);
and U24045 (N_24045,N_23747,N_23742);
or U24046 (N_24046,N_23714,N_23945);
nor U24047 (N_24047,N_23762,N_23760);
nor U24048 (N_24048,N_23867,N_23950);
or U24049 (N_24049,N_23938,N_23759);
nor U24050 (N_24050,N_23809,N_23784);
xnor U24051 (N_24051,N_23990,N_23740);
or U24052 (N_24052,N_23946,N_23802);
or U24053 (N_24053,N_23719,N_23836);
xor U24054 (N_24054,N_23907,N_23964);
nand U24055 (N_24055,N_23711,N_23880);
xor U24056 (N_24056,N_23973,N_23847);
xnor U24057 (N_24057,N_23717,N_23846);
nand U24058 (N_24058,N_23707,N_23753);
and U24059 (N_24059,N_23731,N_23748);
xnor U24060 (N_24060,N_23866,N_23986);
nand U24061 (N_24061,N_23783,N_23725);
xnor U24062 (N_24062,N_23710,N_23873);
nand U24063 (N_24063,N_23845,N_23806);
or U24064 (N_24064,N_23966,N_23708);
or U24065 (N_24065,N_23723,N_23793);
or U24066 (N_24066,N_23994,N_23897);
nand U24067 (N_24067,N_23960,N_23898);
xor U24068 (N_24068,N_23831,N_23888);
nand U24069 (N_24069,N_23703,N_23939);
or U24070 (N_24070,N_23858,N_23726);
or U24071 (N_24071,N_23834,N_23822);
nor U24072 (N_24072,N_23720,N_23860);
and U24073 (N_24073,N_23980,N_23917);
nor U24074 (N_24074,N_23787,N_23716);
xor U24075 (N_24075,N_23944,N_23730);
and U24076 (N_24076,N_23871,N_23923);
nor U24077 (N_24077,N_23808,N_23878);
xor U24078 (N_24078,N_23804,N_23972);
nor U24079 (N_24079,N_23743,N_23796);
nand U24080 (N_24080,N_23810,N_23925);
nand U24081 (N_24081,N_23777,N_23957);
or U24082 (N_24082,N_23838,N_23882);
nor U24083 (N_24083,N_23985,N_23969);
and U24084 (N_24084,N_23844,N_23729);
or U24085 (N_24085,N_23874,N_23790);
nand U24086 (N_24086,N_23837,N_23828);
and U24087 (N_24087,N_23744,N_23968);
xnor U24088 (N_24088,N_23735,N_23750);
nor U24089 (N_24089,N_23977,N_23942);
nor U24090 (N_24090,N_23826,N_23789);
xnor U24091 (N_24091,N_23961,N_23892);
xor U24092 (N_24092,N_23916,N_23782);
and U24093 (N_24093,N_23755,N_23974);
nor U24094 (N_24094,N_23855,N_23899);
and U24095 (N_24095,N_23770,N_23749);
nand U24096 (N_24096,N_23901,N_23786);
or U24097 (N_24097,N_23954,N_23896);
and U24098 (N_24098,N_23900,N_23705);
nand U24099 (N_24099,N_23905,N_23741);
nand U24100 (N_24100,N_23832,N_23876);
xor U24101 (N_24101,N_23976,N_23854);
and U24102 (N_24102,N_23881,N_23924);
xnor U24103 (N_24103,N_23825,N_23861);
and U24104 (N_24104,N_23894,N_23862);
nor U24105 (N_24105,N_23780,N_23940);
nand U24106 (N_24106,N_23956,N_23912);
nor U24107 (N_24107,N_23904,N_23913);
xor U24108 (N_24108,N_23724,N_23818);
or U24109 (N_24109,N_23886,N_23870);
nand U24110 (N_24110,N_23958,N_23962);
nor U24111 (N_24111,N_23737,N_23941);
nand U24112 (N_24112,N_23982,N_23989);
or U24113 (N_24113,N_23795,N_23745);
xor U24114 (N_24114,N_23918,N_23920);
xnor U24115 (N_24115,N_23891,N_23988);
nor U24116 (N_24116,N_23821,N_23823);
nand U24117 (N_24117,N_23778,N_23850);
nand U24118 (N_24118,N_23911,N_23701);
xnor U24119 (N_24119,N_23967,N_23700);
and U24120 (N_24120,N_23738,N_23733);
nor U24121 (N_24121,N_23935,N_23856);
or U24122 (N_24122,N_23779,N_23979);
nor U24123 (N_24123,N_23998,N_23992);
nand U24124 (N_24124,N_23706,N_23835);
or U24125 (N_24125,N_23963,N_23773);
nor U24126 (N_24126,N_23727,N_23929);
nor U24127 (N_24127,N_23971,N_23864);
nand U24128 (N_24128,N_23953,N_23839);
or U24129 (N_24129,N_23776,N_23732);
nand U24130 (N_24130,N_23791,N_23794);
or U24131 (N_24131,N_23987,N_23903);
and U24132 (N_24132,N_23840,N_23774);
nand U24133 (N_24133,N_23713,N_23781);
and U24134 (N_24134,N_23984,N_23877);
nor U24135 (N_24135,N_23909,N_23890);
and U24136 (N_24136,N_23927,N_23995);
and U24137 (N_24137,N_23772,N_23797);
and U24138 (N_24138,N_23883,N_23884);
and U24139 (N_24139,N_23820,N_23768);
nand U24140 (N_24140,N_23906,N_23951);
nand U24141 (N_24141,N_23830,N_23959);
or U24142 (N_24142,N_23792,N_23937);
or U24143 (N_24143,N_23816,N_23709);
nor U24144 (N_24144,N_23798,N_23908);
and U24145 (N_24145,N_23865,N_23712);
xnor U24146 (N_24146,N_23815,N_23928);
xor U24147 (N_24147,N_23812,N_23754);
xor U24148 (N_24148,N_23932,N_23853);
xor U24149 (N_24149,N_23819,N_23763);
and U24150 (N_24150,N_23969,N_23942);
nor U24151 (N_24151,N_23935,N_23764);
nand U24152 (N_24152,N_23705,N_23997);
and U24153 (N_24153,N_23988,N_23733);
nand U24154 (N_24154,N_23892,N_23753);
xnor U24155 (N_24155,N_23937,N_23832);
or U24156 (N_24156,N_23864,N_23947);
nor U24157 (N_24157,N_23876,N_23751);
nand U24158 (N_24158,N_23922,N_23823);
xnor U24159 (N_24159,N_23714,N_23724);
or U24160 (N_24160,N_23990,N_23753);
and U24161 (N_24161,N_23846,N_23809);
xnor U24162 (N_24162,N_23962,N_23978);
and U24163 (N_24163,N_23848,N_23926);
or U24164 (N_24164,N_23777,N_23734);
or U24165 (N_24165,N_23998,N_23847);
and U24166 (N_24166,N_23817,N_23827);
or U24167 (N_24167,N_23881,N_23928);
nor U24168 (N_24168,N_23964,N_23889);
xnor U24169 (N_24169,N_23888,N_23936);
and U24170 (N_24170,N_23765,N_23810);
xnor U24171 (N_24171,N_23872,N_23929);
xor U24172 (N_24172,N_23910,N_23767);
nand U24173 (N_24173,N_23810,N_23829);
and U24174 (N_24174,N_23904,N_23962);
nor U24175 (N_24175,N_23851,N_23803);
xor U24176 (N_24176,N_23764,N_23735);
and U24177 (N_24177,N_23881,N_23979);
or U24178 (N_24178,N_23702,N_23725);
nor U24179 (N_24179,N_23893,N_23967);
nand U24180 (N_24180,N_23701,N_23764);
nand U24181 (N_24181,N_23903,N_23921);
xor U24182 (N_24182,N_23773,N_23843);
nor U24183 (N_24183,N_23894,N_23992);
or U24184 (N_24184,N_23833,N_23780);
or U24185 (N_24185,N_23865,N_23756);
nor U24186 (N_24186,N_23926,N_23794);
xnor U24187 (N_24187,N_23723,N_23808);
nand U24188 (N_24188,N_23986,N_23969);
and U24189 (N_24189,N_23855,N_23719);
or U24190 (N_24190,N_23835,N_23981);
or U24191 (N_24191,N_23973,N_23784);
or U24192 (N_24192,N_23835,N_23902);
nor U24193 (N_24193,N_23782,N_23724);
and U24194 (N_24194,N_23820,N_23723);
and U24195 (N_24195,N_23935,N_23866);
or U24196 (N_24196,N_23868,N_23796);
and U24197 (N_24197,N_23937,N_23897);
nor U24198 (N_24198,N_23804,N_23763);
nor U24199 (N_24199,N_23719,N_23903);
xnor U24200 (N_24200,N_23918,N_23992);
nor U24201 (N_24201,N_23767,N_23799);
and U24202 (N_24202,N_23951,N_23734);
nor U24203 (N_24203,N_23799,N_23975);
nor U24204 (N_24204,N_23773,N_23789);
xnor U24205 (N_24205,N_23722,N_23788);
nor U24206 (N_24206,N_23794,N_23978);
nor U24207 (N_24207,N_23944,N_23964);
or U24208 (N_24208,N_23835,N_23787);
nand U24209 (N_24209,N_23751,N_23740);
xor U24210 (N_24210,N_23812,N_23743);
or U24211 (N_24211,N_23931,N_23933);
or U24212 (N_24212,N_23827,N_23749);
nand U24213 (N_24213,N_23807,N_23780);
nor U24214 (N_24214,N_23891,N_23894);
xor U24215 (N_24215,N_23743,N_23929);
xnor U24216 (N_24216,N_23746,N_23964);
and U24217 (N_24217,N_23956,N_23982);
and U24218 (N_24218,N_23876,N_23975);
or U24219 (N_24219,N_23765,N_23701);
nor U24220 (N_24220,N_23899,N_23726);
nor U24221 (N_24221,N_23886,N_23895);
nand U24222 (N_24222,N_23908,N_23881);
or U24223 (N_24223,N_23817,N_23857);
nand U24224 (N_24224,N_23746,N_23872);
nand U24225 (N_24225,N_23715,N_23785);
xnor U24226 (N_24226,N_23839,N_23890);
nand U24227 (N_24227,N_23718,N_23809);
and U24228 (N_24228,N_23735,N_23881);
and U24229 (N_24229,N_23790,N_23727);
xnor U24230 (N_24230,N_23947,N_23928);
nor U24231 (N_24231,N_23702,N_23827);
xnor U24232 (N_24232,N_23749,N_23958);
or U24233 (N_24233,N_23748,N_23713);
nand U24234 (N_24234,N_23714,N_23708);
or U24235 (N_24235,N_23780,N_23777);
or U24236 (N_24236,N_23899,N_23918);
or U24237 (N_24237,N_23991,N_23958);
nor U24238 (N_24238,N_23920,N_23702);
nand U24239 (N_24239,N_23988,N_23983);
nor U24240 (N_24240,N_23877,N_23822);
nor U24241 (N_24241,N_23824,N_23803);
and U24242 (N_24242,N_23766,N_23889);
and U24243 (N_24243,N_23726,N_23990);
xor U24244 (N_24244,N_23961,N_23927);
or U24245 (N_24245,N_23894,N_23913);
or U24246 (N_24246,N_23774,N_23975);
nand U24247 (N_24247,N_23958,N_23712);
nor U24248 (N_24248,N_23792,N_23848);
nand U24249 (N_24249,N_23737,N_23972);
and U24250 (N_24250,N_23709,N_23839);
nor U24251 (N_24251,N_23846,N_23730);
nand U24252 (N_24252,N_23882,N_23887);
and U24253 (N_24253,N_23727,N_23930);
nand U24254 (N_24254,N_23728,N_23853);
and U24255 (N_24255,N_23952,N_23891);
nand U24256 (N_24256,N_23789,N_23745);
xor U24257 (N_24257,N_23743,N_23872);
xnor U24258 (N_24258,N_23966,N_23913);
nor U24259 (N_24259,N_23767,N_23878);
nor U24260 (N_24260,N_23924,N_23741);
xor U24261 (N_24261,N_23787,N_23794);
xor U24262 (N_24262,N_23717,N_23748);
xor U24263 (N_24263,N_23926,N_23819);
nor U24264 (N_24264,N_23941,N_23928);
xnor U24265 (N_24265,N_23880,N_23723);
or U24266 (N_24266,N_23873,N_23946);
nand U24267 (N_24267,N_23987,N_23765);
nand U24268 (N_24268,N_23883,N_23784);
xor U24269 (N_24269,N_23752,N_23932);
or U24270 (N_24270,N_23982,N_23765);
nor U24271 (N_24271,N_23988,N_23869);
nor U24272 (N_24272,N_23838,N_23941);
or U24273 (N_24273,N_23814,N_23932);
or U24274 (N_24274,N_23973,N_23841);
xor U24275 (N_24275,N_23917,N_23861);
or U24276 (N_24276,N_23999,N_23872);
and U24277 (N_24277,N_23856,N_23990);
nand U24278 (N_24278,N_23956,N_23771);
xnor U24279 (N_24279,N_23749,N_23934);
nor U24280 (N_24280,N_23794,N_23703);
nand U24281 (N_24281,N_23998,N_23997);
nand U24282 (N_24282,N_23741,N_23910);
nor U24283 (N_24283,N_23905,N_23721);
or U24284 (N_24284,N_23865,N_23799);
nor U24285 (N_24285,N_23903,N_23923);
nand U24286 (N_24286,N_23805,N_23709);
nand U24287 (N_24287,N_23918,N_23975);
nand U24288 (N_24288,N_23919,N_23790);
or U24289 (N_24289,N_23785,N_23767);
and U24290 (N_24290,N_23792,N_23705);
or U24291 (N_24291,N_23814,N_23885);
and U24292 (N_24292,N_23877,N_23789);
nor U24293 (N_24293,N_23960,N_23882);
nor U24294 (N_24294,N_23926,N_23885);
or U24295 (N_24295,N_23887,N_23776);
xnor U24296 (N_24296,N_23891,N_23950);
nor U24297 (N_24297,N_23956,N_23746);
nand U24298 (N_24298,N_23928,N_23983);
xor U24299 (N_24299,N_23966,N_23826);
or U24300 (N_24300,N_24230,N_24157);
nand U24301 (N_24301,N_24147,N_24148);
and U24302 (N_24302,N_24040,N_24134);
or U24303 (N_24303,N_24237,N_24196);
or U24304 (N_24304,N_24140,N_24082);
xnor U24305 (N_24305,N_24116,N_24167);
nand U24306 (N_24306,N_24276,N_24264);
nor U24307 (N_24307,N_24011,N_24117);
nand U24308 (N_24308,N_24164,N_24259);
nand U24309 (N_24309,N_24071,N_24168);
and U24310 (N_24310,N_24240,N_24008);
and U24311 (N_24311,N_24278,N_24097);
and U24312 (N_24312,N_24246,N_24266);
and U24313 (N_24313,N_24154,N_24214);
and U24314 (N_24314,N_24221,N_24138);
and U24315 (N_24315,N_24195,N_24085);
nand U24316 (N_24316,N_24223,N_24174);
nor U24317 (N_24317,N_24067,N_24075);
and U24318 (N_24318,N_24247,N_24204);
nor U24319 (N_24319,N_24038,N_24182);
nand U24320 (N_24320,N_24050,N_24072);
xnor U24321 (N_24321,N_24288,N_24025);
nand U24322 (N_24322,N_24143,N_24163);
nor U24323 (N_24323,N_24131,N_24216);
or U24324 (N_24324,N_24233,N_24091);
nor U24325 (N_24325,N_24009,N_24136);
nor U24326 (N_24326,N_24094,N_24274);
xor U24327 (N_24327,N_24291,N_24110);
nor U24328 (N_24328,N_24027,N_24229);
nand U24329 (N_24329,N_24088,N_24206);
or U24330 (N_24330,N_24173,N_24296);
and U24331 (N_24331,N_24107,N_24203);
xnor U24332 (N_24332,N_24297,N_24236);
nor U24333 (N_24333,N_24102,N_24007);
nor U24334 (N_24334,N_24292,N_24033);
nand U24335 (N_24335,N_24244,N_24101);
xnor U24336 (N_24336,N_24257,N_24044);
nor U24337 (N_24337,N_24049,N_24179);
nor U24338 (N_24338,N_24061,N_24153);
nor U24339 (N_24339,N_24202,N_24031);
or U24340 (N_24340,N_24210,N_24087);
nor U24341 (N_24341,N_24205,N_24121);
nor U24342 (N_24342,N_24208,N_24172);
xor U24343 (N_24343,N_24299,N_24263);
or U24344 (N_24344,N_24286,N_24289);
and U24345 (N_24345,N_24238,N_24281);
nor U24346 (N_24346,N_24287,N_24074);
and U24347 (N_24347,N_24267,N_24060);
and U24348 (N_24348,N_24224,N_24066);
nand U24349 (N_24349,N_24184,N_24165);
or U24350 (N_24350,N_24036,N_24218);
and U24351 (N_24351,N_24133,N_24022);
nand U24352 (N_24352,N_24290,N_24078);
nand U24353 (N_24353,N_24190,N_24100);
nand U24354 (N_24354,N_24089,N_24251);
or U24355 (N_24355,N_24029,N_24241);
nand U24356 (N_24356,N_24012,N_24188);
nor U24357 (N_24357,N_24004,N_24255);
nor U24358 (N_24358,N_24169,N_24130);
xnor U24359 (N_24359,N_24144,N_24252);
xnor U24360 (N_24360,N_24059,N_24199);
nand U24361 (N_24361,N_24201,N_24146);
nor U24362 (N_24362,N_24181,N_24096);
and U24363 (N_24363,N_24162,N_24063);
nor U24364 (N_24364,N_24024,N_24177);
nor U24365 (N_24365,N_24000,N_24090);
and U24366 (N_24366,N_24248,N_24084);
nor U24367 (N_24367,N_24242,N_24231);
or U24368 (N_24368,N_24023,N_24217);
nor U24369 (N_24369,N_24282,N_24200);
and U24370 (N_24370,N_24080,N_24285);
nor U24371 (N_24371,N_24209,N_24260);
nand U24372 (N_24372,N_24211,N_24037);
or U24373 (N_24373,N_24152,N_24120);
and U24374 (N_24374,N_24207,N_24086);
nor U24375 (N_24375,N_24149,N_24034);
nand U24376 (N_24376,N_24175,N_24032);
or U24377 (N_24377,N_24064,N_24092);
or U24378 (N_24378,N_24010,N_24056);
nor U24379 (N_24379,N_24076,N_24052);
nor U24380 (N_24380,N_24258,N_24113);
nand U24381 (N_24381,N_24161,N_24159);
nand U24382 (N_24382,N_24176,N_24283);
or U24383 (N_24383,N_24171,N_24020);
nand U24384 (N_24384,N_24268,N_24180);
or U24385 (N_24385,N_24099,N_24279);
xor U24386 (N_24386,N_24127,N_24243);
and U24387 (N_24387,N_24095,N_24077);
xnor U24388 (N_24388,N_24232,N_24235);
or U24389 (N_24389,N_24277,N_24017);
or U24390 (N_24390,N_24272,N_24114);
and U24391 (N_24391,N_24122,N_24189);
nor U24392 (N_24392,N_24119,N_24270);
xor U24393 (N_24393,N_24129,N_24055);
or U24394 (N_24394,N_24013,N_24108);
nand U24395 (N_24395,N_24105,N_24228);
or U24396 (N_24396,N_24141,N_24135);
nor U24397 (N_24397,N_24225,N_24170);
nand U24398 (N_24398,N_24058,N_24001);
or U24399 (N_24399,N_24193,N_24028);
nand U24400 (N_24400,N_24098,N_24271);
nor U24401 (N_24401,N_24021,N_24178);
nand U24402 (N_24402,N_24018,N_24226);
nand U24403 (N_24403,N_24045,N_24003);
nor U24404 (N_24404,N_24262,N_24043);
nand U24405 (N_24405,N_24115,N_24124);
xnor U24406 (N_24406,N_24106,N_24126);
or U24407 (N_24407,N_24123,N_24273);
nand U24408 (N_24408,N_24215,N_24269);
xnor U24409 (N_24409,N_24185,N_24132);
nor U24410 (N_24410,N_24249,N_24068);
and U24411 (N_24411,N_24198,N_24142);
xnor U24412 (N_24412,N_24245,N_24042);
xnor U24413 (N_24413,N_24053,N_24227);
or U24414 (N_24414,N_24019,N_24139);
nor U24415 (N_24415,N_24051,N_24026);
nor U24416 (N_24416,N_24006,N_24057);
and U24417 (N_24417,N_24111,N_24093);
nand U24418 (N_24418,N_24239,N_24030);
nand U24419 (N_24419,N_24158,N_24222);
nand U24420 (N_24420,N_24219,N_24081);
nand U24421 (N_24421,N_24253,N_24234);
nand U24422 (N_24422,N_24194,N_24039);
and U24423 (N_24423,N_24160,N_24294);
xor U24424 (N_24424,N_24212,N_24250);
or U24425 (N_24425,N_24014,N_24293);
nand U24426 (N_24426,N_24070,N_24083);
nand U24427 (N_24427,N_24284,N_24192);
or U24428 (N_24428,N_24150,N_24275);
nor U24429 (N_24429,N_24002,N_24104);
nor U24430 (N_24430,N_24261,N_24295);
and U24431 (N_24431,N_24073,N_24186);
or U24432 (N_24432,N_24128,N_24191);
and U24433 (N_24433,N_24125,N_24145);
or U24434 (N_24434,N_24015,N_24155);
or U24435 (N_24435,N_24156,N_24137);
xor U24436 (N_24436,N_24265,N_24118);
nor U24437 (N_24437,N_24035,N_24079);
or U24438 (N_24438,N_24220,N_24048);
nand U24439 (N_24439,N_24254,N_24183);
and U24440 (N_24440,N_24112,N_24047);
nor U24441 (N_24441,N_24280,N_24062);
nor U24442 (N_24442,N_24016,N_24256);
or U24443 (N_24443,N_24103,N_24069);
nor U24444 (N_24444,N_24197,N_24041);
or U24445 (N_24445,N_24046,N_24151);
xor U24446 (N_24446,N_24213,N_24166);
and U24447 (N_24447,N_24187,N_24065);
nor U24448 (N_24448,N_24054,N_24109);
nor U24449 (N_24449,N_24298,N_24005);
or U24450 (N_24450,N_24041,N_24182);
nor U24451 (N_24451,N_24287,N_24195);
and U24452 (N_24452,N_24273,N_24260);
nand U24453 (N_24453,N_24016,N_24125);
nand U24454 (N_24454,N_24119,N_24006);
and U24455 (N_24455,N_24280,N_24132);
nor U24456 (N_24456,N_24162,N_24098);
or U24457 (N_24457,N_24176,N_24023);
or U24458 (N_24458,N_24012,N_24278);
and U24459 (N_24459,N_24211,N_24227);
nand U24460 (N_24460,N_24131,N_24237);
or U24461 (N_24461,N_24216,N_24165);
and U24462 (N_24462,N_24160,N_24186);
nand U24463 (N_24463,N_24084,N_24028);
xor U24464 (N_24464,N_24102,N_24107);
xnor U24465 (N_24465,N_24027,N_24179);
xor U24466 (N_24466,N_24015,N_24147);
xnor U24467 (N_24467,N_24240,N_24253);
or U24468 (N_24468,N_24017,N_24269);
or U24469 (N_24469,N_24290,N_24083);
nor U24470 (N_24470,N_24092,N_24009);
xor U24471 (N_24471,N_24110,N_24028);
and U24472 (N_24472,N_24203,N_24082);
nand U24473 (N_24473,N_24233,N_24128);
or U24474 (N_24474,N_24206,N_24131);
or U24475 (N_24475,N_24132,N_24114);
xnor U24476 (N_24476,N_24040,N_24154);
xor U24477 (N_24477,N_24008,N_24022);
nand U24478 (N_24478,N_24290,N_24151);
or U24479 (N_24479,N_24133,N_24171);
nand U24480 (N_24480,N_24096,N_24139);
nor U24481 (N_24481,N_24098,N_24042);
or U24482 (N_24482,N_24147,N_24277);
xor U24483 (N_24483,N_24274,N_24247);
nor U24484 (N_24484,N_24084,N_24227);
xnor U24485 (N_24485,N_24079,N_24046);
or U24486 (N_24486,N_24178,N_24181);
xnor U24487 (N_24487,N_24189,N_24229);
or U24488 (N_24488,N_24174,N_24010);
and U24489 (N_24489,N_24068,N_24145);
and U24490 (N_24490,N_24161,N_24147);
and U24491 (N_24491,N_24040,N_24228);
nor U24492 (N_24492,N_24148,N_24265);
and U24493 (N_24493,N_24274,N_24144);
and U24494 (N_24494,N_24083,N_24221);
and U24495 (N_24495,N_24136,N_24192);
or U24496 (N_24496,N_24263,N_24208);
or U24497 (N_24497,N_24138,N_24249);
nand U24498 (N_24498,N_24009,N_24299);
nand U24499 (N_24499,N_24062,N_24244);
or U24500 (N_24500,N_24066,N_24293);
and U24501 (N_24501,N_24239,N_24167);
xor U24502 (N_24502,N_24006,N_24090);
xor U24503 (N_24503,N_24133,N_24044);
nor U24504 (N_24504,N_24029,N_24231);
nand U24505 (N_24505,N_24234,N_24146);
xor U24506 (N_24506,N_24215,N_24091);
and U24507 (N_24507,N_24002,N_24132);
and U24508 (N_24508,N_24052,N_24110);
or U24509 (N_24509,N_24294,N_24159);
and U24510 (N_24510,N_24174,N_24290);
nand U24511 (N_24511,N_24284,N_24020);
nand U24512 (N_24512,N_24238,N_24198);
and U24513 (N_24513,N_24152,N_24073);
or U24514 (N_24514,N_24226,N_24295);
and U24515 (N_24515,N_24236,N_24086);
or U24516 (N_24516,N_24155,N_24028);
and U24517 (N_24517,N_24151,N_24007);
nor U24518 (N_24518,N_24054,N_24237);
xor U24519 (N_24519,N_24147,N_24149);
xnor U24520 (N_24520,N_24228,N_24084);
nor U24521 (N_24521,N_24220,N_24181);
nand U24522 (N_24522,N_24169,N_24193);
nand U24523 (N_24523,N_24134,N_24280);
nor U24524 (N_24524,N_24121,N_24152);
nor U24525 (N_24525,N_24105,N_24124);
or U24526 (N_24526,N_24247,N_24152);
and U24527 (N_24527,N_24081,N_24075);
nor U24528 (N_24528,N_24078,N_24021);
xnor U24529 (N_24529,N_24258,N_24181);
and U24530 (N_24530,N_24190,N_24137);
nand U24531 (N_24531,N_24133,N_24024);
nand U24532 (N_24532,N_24038,N_24007);
xor U24533 (N_24533,N_24002,N_24226);
and U24534 (N_24534,N_24220,N_24208);
nor U24535 (N_24535,N_24188,N_24174);
and U24536 (N_24536,N_24269,N_24271);
nand U24537 (N_24537,N_24023,N_24265);
nor U24538 (N_24538,N_24075,N_24145);
and U24539 (N_24539,N_24069,N_24062);
nor U24540 (N_24540,N_24180,N_24239);
xor U24541 (N_24541,N_24125,N_24037);
and U24542 (N_24542,N_24179,N_24232);
nand U24543 (N_24543,N_24168,N_24155);
xnor U24544 (N_24544,N_24213,N_24251);
xor U24545 (N_24545,N_24101,N_24248);
nand U24546 (N_24546,N_24181,N_24249);
or U24547 (N_24547,N_24097,N_24275);
or U24548 (N_24548,N_24057,N_24068);
and U24549 (N_24549,N_24120,N_24258);
or U24550 (N_24550,N_24116,N_24141);
nor U24551 (N_24551,N_24012,N_24054);
nor U24552 (N_24552,N_24234,N_24144);
nor U24553 (N_24553,N_24036,N_24048);
and U24554 (N_24554,N_24024,N_24119);
nor U24555 (N_24555,N_24000,N_24159);
nor U24556 (N_24556,N_24173,N_24198);
and U24557 (N_24557,N_24195,N_24116);
nand U24558 (N_24558,N_24095,N_24122);
or U24559 (N_24559,N_24087,N_24024);
nand U24560 (N_24560,N_24119,N_24054);
and U24561 (N_24561,N_24175,N_24271);
and U24562 (N_24562,N_24070,N_24249);
xnor U24563 (N_24563,N_24198,N_24208);
and U24564 (N_24564,N_24296,N_24225);
and U24565 (N_24565,N_24278,N_24212);
and U24566 (N_24566,N_24270,N_24002);
nor U24567 (N_24567,N_24242,N_24085);
nor U24568 (N_24568,N_24024,N_24279);
and U24569 (N_24569,N_24210,N_24102);
nand U24570 (N_24570,N_24233,N_24287);
nor U24571 (N_24571,N_24263,N_24191);
or U24572 (N_24572,N_24143,N_24215);
and U24573 (N_24573,N_24296,N_24171);
nor U24574 (N_24574,N_24179,N_24001);
and U24575 (N_24575,N_24136,N_24061);
and U24576 (N_24576,N_24277,N_24215);
nor U24577 (N_24577,N_24189,N_24277);
xnor U24578 (N_24578,N_24061,N_24194);
xor U24579 (N_24579,N_24052,N_24163);
nand U24580 (N_24580,N_24264,N_24088);
and U24581 (N_24581,N_24173,N_24069);
nor U24582 (N_24582,N_24256,N_24182);
and U24583 (N_24583,N_24167,N_24080);
nand U24584 (N_24584,N_24283,N_24109);
xor U24585 (N_24585,N_24211,N_24162);
xnor U24586 (N_24586,N_24207,N_24214);
xnor U24587 (N_24587,N_24182,N_24258);
xnor U24588 (N_24588,N_24054,N_24268);
and U24589 (N_24589,N_24103,N_24296);
nor U24590 (N_24590,N_24102,N_24173);
nand U24591 (N_24591,N_24263,N_24200);
xnor U24592 (N_24592,N_24257,N_24299);
nand U24593 (N_24593,N_24143,N_24066);
or U24594 (N_24594,N_24159,N_24066);
or U24595 (N_24595,N_24259,N_24071);
or U24596 (N_24596,N_24219,N_24232);
nand U24597 (N_24597,N_24242,N_24022);
or U24598 (N_24598,N_24247,N_24196);
nand U24599 (N_24599,N_24094,N_24195);
nand U24600 (N_24600,N_24509,N_24331);
and U24601 (N_24601,N_24465,N_24404);
and U24602 (N_24602,N_24420,N_24400);
or U24603 (N_24603,N_24410,N_24334);
or U24604 (N_24604,N_24387,N_24514);
and U24605 (N_24605,N_24542,N_24344);
and U24606 (N_24606,N_24586,N_24375);
and U24607 (N_24607,N_24392,N_24581);
or U24608 (N_24608,N_24524,N_24516);
xnor U24609 (N_24609,N_24498,N_24385);
or U24610 (N_24610,N_24541,N_24356);
and U24611 (N_24611,N_24429,N_24533);
or U24612 (N_24612,N_24565,N_24376);
nor U24613 (N_24613,N_24560,N_24348);
xnor U24614 (N_24614,N_24557,N_24324);
nor U24615 (N_24615,N_24545,N_24361);
and U24616 (N_24616,N_24489,N_24415);
nor U24617 (N_24617,N_24412,N_24580);
nor U24618 (N_24618,N_24468,N_24578);
nand U24619 (N_24619,N_24366,N_24561);
nand U24620 (N_24620,N_24590,N_24474);
and U24621 (N_24621,N_24496,N_24443);
xnor U24622 (N_24622,N_24493,N_24364);
or U24623 (N_24623,N_24574,N_24510);
nand U24624 (N_24624,N_24491,N_24372);
nand U24625 (N_24625,N_24359,N_24351);
nand U24626 (N_24626,N_24582,N_24502);
xor U24627 (N_24627,N_24454,N_24480);
xor U24628 (N_24628,N_24587,N_24492);
nor U24629 (N_24629,N_24529,N_24437);
xnor U24630 (N_24630,N_24520,N_24576);
xnor U24631 (N_24631,N_24579,N_24540);
xor U24632 (N_24632,N_24483,N_24471);
nand U24633 (N_24633,N_24575,N_24534);
and U24634 (N_24634,N_24414,N_24456);
and U24635 (N_24635,N_24511,N_24597);
xor U24636 (N_24636,N_24304,N_24409);
or U24637 (N_24637,N_24390,N_24365);
nor U24638 (N_24638,N_24428,N_24399);
or U24639 (N_24639,N_24380,N_24316);
nor U24640 (N_24640,N_24452,N_24338);
and U24641 (N_24641,N_24459,N_24401);
nor U24642 (N_24642,N_24558,N_24537);
nor U24643 (N_24643,N_24431,N_24320);
nand U24644 (N_24644,N_24595,N_24333);
nand U24645 (N_24645,N_24583,N_24307);
or U24646 (N_24646,N_24588,N_24360);
and U24647 (N_24647,N_24310,N_24425);
nor U24648 (N_24648,N_24355,N_24473);
or U24649 (N_24649,N_24552,N_24463);
nand U24650 (N_24650,N_24345,N_24423);
or U24651 (N_24651,N_24330,N_24599);
xnor U24652 (N_24652,N_24556,N_24469);
and U24653 (N_24653,N_24317,N_24354);
xor U24654 (N_24654,N_24477,N_24551);
xor U24655 (N_24655,N_24306,N_24593);
nor U24656 (N_24656,N_24417,N_24538);
nand U24657 (N_24657,N_24536,N_24357);
nor U24658 (N_24658,N_24455,N_24315);
or U24659 (N_24659,N_24403,N_24508);
and U24660 (N_24660,N_24384,N_24460);
and U24661 (N_24661,N_24475,N_24362);
xor U24662 (N_24662,N_24346,N_24393);
or U24663 (N_24663,N_24594,N_24373);
xor U24664 (N_24664,N_24577,N_24523);
nor U24665 (N_24665,N_24497,N_24458);
xor U24666 (N_24666,N_24518,N_24381);
nor U24667 (N_24667,N_24548,N_24563);
nor U24668 (N_24668,N_24323,N_24451);
nand U24669 (N_24669,N_24522,N_24379);
nor U24670 (N_24670,N_24457,N_24433);
nand U24671 (N_24671,N_24314,N_24539);
nand U24672 (N_24672,N_24371,N_24300);
or U24673 (N_24673,N_24513,N_24466);
or U24674 (N_24674,N_24564,N_24391);
or U24675 (N_24675,N_24569,N_24506);
or U24676 (N_24676,N_24439,N_24305);
and U24677 (N_24677,N_24573,N_24419);
xor U24678 (N_24678,N_24313,N_24377);
and U24679 (N_24679,N_24318,N_24369);
xor U24680 (N_24680,N_24341,N_24544);
nor U24681 (N_24681,N_24440,N_24407);
and U24682 (N_24682,N_24535,N_24405);
xnor U24683 (N_24683,N_24462,N_24447);
xor U24684 (N_24684,N_24589,N_24461);
or U24685 (N_24685,N_24470,N_24505);
xor U24686 (N_24686,N_24389,N_24309);
and U24687 (N_24687,N_24430,N_24519);
nor U24688 (N_24688,N_24490,N_24485);
xor U24689 (N_24689,N_24350,N_24528);
xor U24690 (N_24690,N_24402,N_24396);
nand U24691 (N_24691,N_24435,N_24571);
nor U24692 (N_24692,N_24453,N_24386);
xor U24693 (N_24693,N_24352,N_24449);
nand U24694 (N_24694,N_24500,N_24559);
or U24695 (N_24695,N_24398,N_24358);
xor U24696 (N_24696,N_24416,N_24367);
nor U24697 (N_24697,N_24501,N_24343);
nand U24698 (N_24698,N_24445,N_24572);
nand U24699 (N_24699,N_24312,N_24424);
and U24700 (N_24700,N_24411,N_24598);
or U24701 (N_24701,N_24486,N_24566);
nor U24702 (N_24702,N_24383,N_24467);
and U24703 (N_24703,N_24421,N_24302);
and U24704 (N_24704,N_24531,N_24363);
xnor U24705 (N_24705,N_24340,N_24442);
or U24706 (N_24706,N_24584,N_24327);
nand U24707 (N_24707,N_24394,N_24448);
and U24708 (N_24708,N_24438,N_24413);
nand U24709 (N_24709,N_24503,N_24526);
nor U24710 (N_24710,N_24374,N_24335);
xor U24711 (N_24711,N_24530,N_24408);
or U24712 (N_24712,N_24353,N_24336);
or U24713 (N_24713,N_24507,N_24546);
nand U24714 (N_24714,N_24322,N_24512);
and U24715 (N_24715,N_24476,N_24555);
nor U24716 (N_24716,N_24499,N_24481);
nor U24717 (N_24717,N_24326,N_24418);
nand U24718 (N_24718,N_24446,N_24567);
nor U24719 (N_24719,N_24308,N_24434);
nor U24720 (N_24720,N_24570,N_24311);
xnor U24721 (N_24721,N_24487,N_24432);
xor U24722 (N_24722,N_24479,N_24549);
xor U24723 (N_24723,N_24388,N_24397);
or U24724 (N_24724,N_24321,N_24596);
nor U24725 (N_24725,N_24592,N_24444);
nor U24726 (N_24726,N_24301,N_24543);
and U24727 (N_24727,N_24568,N_24426);
xor U24728 (N_24728,N_24521,N_24337);
nor U24729 (N_24729,N_24378,N_24441);
xor U24730 (N_24730,N_24553,N_24472);
and U24731 (N_24731,N_24550,N_24562);
nor U24732 (N_24732,N_24328,N_24339);
and U24733 (N_24733,N_24585,N_24342);
xnor U24734 (N_24734,N_24464,N_24515);
nor U24735 (N_24735,N_24347,N_24450);
and U24736 (N_24736,N_24303,N_24422);
nor U24737 (N_24737,N_24547,N_24478);
nand U24738 (N_24738,N_24325,N_24332);
nand U24739 (N_24739,N_24484,N_24488);
and U24740 (N_24740,N_24525,N_24517);
nand U24741 (N_24741,N_24495,N_24329);
and U24742 (N_24742,N_24591,N_24504);
or U24743 (N_24743,N_24370,N_24406);
nor U24744 (N_24744,N_24436,N_24427);
or U24745 (N_24745,N_24368,N_24532);
and U24746 (N_24746,N_24382,N_24319);
or U24747 (N_24747,N_24395,N_24527);
and U24748 (N_24748,N_24554,N_24494);
nand U24749 (N_24749,N_24482,N_24349);
xnor U24750 (N_24750,N_24593,N_24314);
xnor U24751 (N_24751,N_24436,N_24339);
or U24752 (N_24752,N_24462,N_24382);
and U24753 (N_24753,N_24597,N_24499);
or U24754 (N_24754,N_24446,N_24388);
and U24755 (N_24755,N_24356,N_24526);
xnor U24756 (N_24756,N_24406,N_24300);
xnor U24757 (N_24757,N_24555,N_24508);
nor U24758 (N_24758,N_24384,N_24323);
xnor U24759 (N_24759,N_24450,N_24513);
nand U24760 (N_24760,N_24328,N_24518);
xor U24761 (N_24761,N_24327,N_24347);
nor U24762 (N_24762,N_24364,N_24434);
and U24763 (N_24763,N_24420,N_24384);
xor U24764 (N_24764,N_24419,N_24393);
nor U24765 (N_24765,N_24355,N_24352);
nor U24766 (N_24766,N_24483,N_24347);
or U24767 (N_24767,N_24597,N_24483);
nand U24768 (N_24768,N_24325,N_24503);
nand U24769 (N_24769,N_24591,N_24345);
and U24770 (N_24770,N_24500,N_24365);
nor U24771 (N_24771,N_24403,N_24518);
and U24772 (N_24772,N_24516,N_24520);
nor U24773 (N_24773,N_24567,N_24580);
nor U24774 (N_24774,N_24514,N_24332);
nand U24775 (N_24775,N_24367,N_24435);
nor U24776 (N_24776,N_24351,N_24418);
nand U24777 (N_24777,N_24325,N_24349);
and U24778 (N_24778,N_24348,N_24539);
and U24779 (N_24779,N_24329,N_24490);
and U24780 (N_24780,N_24325,N_24591);
and U24781 (N_24781,N_24585,N_24557);
nand U24782 (N_24782,N_24340,N_24577);
and U24783 (N_24783,N_24322,N_24367);
or U24784 (N_24784,N_24555,N_24377);
xnor U24785 (N_24785,N_24510,N_24412);
xnor U24786 (N_24786,N_24544,N_24325);
nor U24787 (N_24787,N_24467,N_24566);
or U24788 (N_24788,N_24444,N_24376);
or U24789 (N_24789,N_24441,N_24424);
xnor U24790 (N_24790,N_24556,N_24536);
xnor U24791 (N_24791,N_24529,N_24459);
and U24792 (N_24792,N_24310,N_24309);
and U24793 (N_24793,N_24390,N_24479);
and U24794 (N_24794,N_24359,N_24440);
nor U24795 (N_24795,N_24543,N_24417);
or U24796 (N_24796,N_24499,N_24437);
and U24797 (N_24797,N_24500,N_24513);
nand U24798 (N_24798,N_24508,N_24433);
nor U24799 (N_24799,N_24569,N_24489);
and U24800 (N_24800,N_24509,N_24546);
xnor U24801 (N_24801,N_24449,N_24341);
or U24802 (N_24802,N_24442,N_24528);
nor U24803 (N_24803,N_24339,N_24538);
xnor U24804 (N_24804,N_24431,N_24460);
and U24805 (N_24805,N_24396,N_24302);
xor U24806 (N_24806,N_24340,N_24595);
nor U24807 (N_24807,N_24531,N_24352);
nand U24808 (N_24808,N_24596,N_24341);
nor U24809 (N_24809,N_24370,N_24340);
nor U24810 (N_24810,N_24339,N_24341);
nor U24811 (N_24811,N_24483,N_24449);
and U24812 (N_24812,N_24482,N_24414);
and U24813 (N_24813,N_24362,N_24531);
nor U24814 (N_24814,N_24592,N_24359);
nor U24815 (N_24815,N_24377,N_24322);
nand U24816 (N_24816,N_24333,N_24374);
nand U24817 (N_24817,N_24332,N_24421);
nor U24818 (N_24818,N_24372,N_24574);
or U24819 (N_24819,N_24573,N_24332);
nor U24820 (N_24820,N_24458,N_24541);
xnor U24821 (N_24821,N_24347,N_24383);
xnor U24822 (N_24822,N_24400,N_24344);
nand U24823 (N_24823,N_24568,N_24531);
nand U24824 (N_24824,N_24338,N_24591);
and U24825 (N_24825,N_24432,N_24414);
and U24826 (N_24826,N_24313,N_24385);
xor U24827 (N_24827,N_24322,N_24541);
and U24828 (N_24828,N_24412,N_24332);
xor U24829 (N_24829,N_24395,N_24502);
and U24830 (N_24830,N_24344,N_24555);
xnor U24831 (N_24831,N_24407,N_24477);
nor U24832 (N_24832,N_24449,N_24441);
nor U24833 (N_24833,N_24527,N_24564);
nor U24834 (N_24834,N_24368,N_24569);
xor U24835 (N_24835,N_24478,N_24390);
nor U24836 (N_24836,N_24412,N_24516);
xnor U24837 (N_24837,N_24541,N_24457);
and U24838 (N_24838,N_24554,N_24532);
nor U24839 (N_24839,N_24406,N_24598);
xnor U24840 (N_24840,N_24381,N_24488);
nand U24841 (N_24841,N_24447,N_24371);
nor U24842 (N_24842,N_24414,N_24576);
or U24843 (N_24843,N_24308,N_24366);
nand U24844 (N_24844,N_24338,N_24387);
xor U24845 (N_24845,N_24460,N_24314);
nand U24846 (N_24846,N_24539,N_24344);
xor U24847 (N_24847,N_24424,N_24498);
and U24848 (N_24848,N_24326,N_24371);
nor U24849 (N_24849,N_24318,N_24360);
and U24850 (N_24850,N_24416,N_24374);
xor U24851 (N_24851,N_24552,N_24435);
nand U24852 (N_24852,N_24352,N_24442);
nor U24853 (N_24853,N_24379,N_24418);
nor U24854 (N_24854,N_24319,N_24494);
or U24855 (N_24855,N_24503,N_24369);
or U24856 (N_24856,N_24555,N_24568);
nor U24857 (N_24857,N_24549,N_24323);
xor U24858 (N_24858,N_24501,N_24317);
nand U24859 (N_24859,N_24491,N_24439);
nor U24860 (N_24860,N_24324,N_24351);
xor U24861 (N_24861,N_24459,N_24429);
nand U24862 (N_24862,N_24351,N_24568);
nand U24863 (N_24863,N_24559,N_24561);
xnor U24864 (N_24864,N_24485,N_24321);
nor U24865 (N_24865,N_24306,N_24562);
nor U24866 (N_24866,N_24402,N_24433);
nand U24867 (N_24867,N_24568,N_24427);
nor U24868 (N_24868,N_24390,N_24581);
xor U24869 (N_24869,N_24579,N_24336);
xor U24870 (N_24870,N_24410,N_24512);
or U24871 (N_24871,N_24327,N_24428);
and U24872 (N_24872,N_24462,N_24356);
nor U24873 (N_24873,N_24590,N_24399);
nor U24874 (N_24874,N_24549,N_24424);
xnor U24875 (N_24875,N_24524,N_24451);
nor U24876 (N_24876,N_24488,N_24456);
xnor U24877 (N_24877,N_24584,N_24451);
nand U24878 (N_24878,N_24547,N_24300);
xnor U24879 (N_24879,N_24344,N_24327);
nor U24880 (N_24880,N_24581,N_24498);
nor U24881 (N_24881,N_24358,N_24490);
and U24882 (N_24882,N_24372,N_24427);
xnor U24883 (N_24883,N_24511,N_24313);
and U24884 (N_24884,N_24357,N_24506);
or U24885 (N_24885,N_24365,N_24576);
nor U24886 (N_24886,N_24497,N_24447);
nand U24887 (N_24887,N_24349,N_24305);
and U24888 (N_24888,N_24463,N_24389);
and U24889 (N_24889,N_24573,N_24593);
nor U24890 (N_24890,N_24537,N_24587);
nor U24891 (N_24891,N_24397,N_24540);
or U24892 (N_24892,N_24335,N_24551);
and U24893 (N_24893,N_24497,N_24304);
nor U24894 (N_24894,N_24433,N_24571);
nor U24895 (N_24895,N_24467,N_24319);
nand U24896 (N_24896,N_24427,N_24539);
nand U24897 (N_24897,N_24478,N_24387);
nor U24898 (N_24898,N_24443,N_24465);
xor U24899 (N_24899,N_24431,N_24567);
or U24900 (N_24900,N_24637,N_24839);
nand U24901 (N_24901,N_24765,N_24885);
or U24902 (N_24902,N_24808,N_24797);
nor U24903 (N_24903,N_24620,N_24721);
xor U24904 (N_24904,N_24604,N_24848);
and U24905 (N_24905,N_24898,N_24829);
or U24906 (N_24906,N_24825,N_24840);
xnor U24907 (N_24907,N_24841,N_24695);
nand U24908 (N_24908,N_24785,N_24767);
xor U24909 (N_24909,N_24664,N_24766);
xor U24910 (N_24910,N_24716,N_24856);
xor U24911 (N_24911,N_24728,N_24826);
nand U24912 (N_24912,N_24777,N_24718);
xnor U24913 (N_24913,N_24884,N_24867);
xnor U24914 (N_24914,N_24820,N_24675);
nor U24915 (N_24915,N_24621,N_24630);
or U24916 (N_24916,N_24617,N_24786);
nand U24917 (N_24917,N_24656,N_24871);
nor U24918 (N_24918,N_24883,N_24875);
nand U24919 (N_24919,N_24782,N_24753);
and U24920 (N_24920,N_24763,N_24689);
xor U24921 (N_24921,N_24613,N_24749);
or U24922 (N_24922,N_24691,N_24746);
or U24923 (N_24923,N_24878,N_24877);
nor U24924 (N_24924,N_24838,N_24778);
xnor U24925 (N_24925,N_24636,N_24819);
and U24926 (N_24926,N_24869,N_24633);
nor U24927 (N_24927,N_24654,N_24816);
and U24928 (N_24928,N_24834,N_24876);
xor U24929 (N_24929,N_24639,N_24605);
and U24930 (N_24930,N_24872,N_24791);
and U24931 (N_24931,N_24655,N_24892);
and U24932 (N_24932,N_24804,N_24762);
and U24933 (N_24933,N_24806,N_24852);
or U24934 (N_24934,N_24851,N_24625);
and U24935 (N_24935,N_24739,N_24824);
xor U24936 (N_24936,N_24775,N_24814);
and U24937 (N_24937,N_24607,N_24756);
or U24938 (N_24938,N_24711,N_24671);
nor U24939 (N_24939,N_24652,N_24653);
nor U24940 (N_24940,N_24635,N_24812);
xnor U24941 (N_24941,N_24809,N_24729);
xnor U24942 (N_24942,N_24678,N_24703);
xnor U24943 (N_24943,N_24609,N_24815);
and U24944 (N_24944,N_24614,N_24865);
xnor U24945 (N_24945,N_24895,N_24685);
nand U24946 (N_24946,N_24744,N_24626);
nand U24947 (N_24947,N_24798,N_24833);
xnor U24948 (N_24948,N_24686,N_24890);
nand U24949 (N_24949,N_24725,N_24684);
or U24950 (N_24950,N_24880,N_24759);
nand U24951 (N_24951,N_24602,N_24757);
and U24952 (N_24952,N_24855,N_24616);
or U24953 (N_24953,N_24781,N_24672);
nor U24954 (N_24954,N_24611,N_24835);
nand U24955 (N_24955,N_24854,N_24697);
xor U24956 (N_24956,N_24836,N_24717);
nand U24957 (N_24957,N_24669,N_24667);
xnor U24958 (N_24958,N_24747,N_24692);
nand U24959 (N_24959,N_24722,N_24640);
nand U24960 (N_24960,N_24790,N_24683);
nor U24961 (N_24961,N_24748,N_24649);
nand U24962 (N_24962,N_24868,N_24849);
xnor U24963 (N_24963,N_24770,N_24817);
and U24964 (N_24964,N_24774,N_24870);
xor U24965 (N_24965,N_24874,N_24634);
xnor U24966 (N_24966,N_24641,N_24643);
and U24967 (N_24967,N_24623,N_24818);
or U24968 (N_24968,N_24795,N_24730);
nand U24969 (N_24969,N_24807,N_24644);
xnor U24970 (N_24970,N_24688,N_24881);
xnor U24971 (N_24971,N_24862,N_24801);
nor U24972 (N_24972,N_24680,N_24648);
xor U24973 (N_24973,N_24891,N_24896);
nor U24974 (N_24974,N_24708,N_24600);
nor U24975 (N_24975,N_24886,N_24732);
nor U24976 (N_24976,N_24823,N_24647);
or U24977 (N_24977,N_24779,N_24745);
nor U24978 (N_24978,N_24857,N_24670);
nand U24979 (N_24979,N_24610,N_24735);
and U24980 (N_24980,N_24666,N_24789);
and U24981 (N_24981,N_24603,N_24741);
xor U24982 (N_24982,N_24776,N_24661);
and U24983 (N_24983,N_24632,N_24631);
nand U24984 (N_24984,N_24679,N_24887);
or U24985 (N_24985,N_24743,N_24690);
and U24986 (N_24986,N_24780,N_24837);
xnor U24987 (N_24987,N_24805,N_24752);
nand U24988 (N_24988,N_24698,N_24799);
xnor U24989 (N_24989,N_24802,N_24897);
nor U24990 (N_24990,N_24737,N_24783);
or U24991 (N_24991,N_24657,N_24699);
or U24992 (N_24992,N_24662,N_24676);
xnor U24993 (N_24993,N_24750,N_24832);
xnor U24994 (N_24994,N_24642,N_24638);
nor U24995 (N_24995,N_24701,N_24754);
xor U24996 (N_24996,N_24810,N_24793);
or U24997 (N_24997,N_24788,N_24758);
nand U24998 (N_24998,N_24707,N_24850);
nor U24999 (N_24999,N_24822,N_24608);
nor U25000 (N_25000,N_24612,N_24659);
nor U25001 (N_25001,N_24860,N_24742);
nand U25002 (N_25002,N_24682,N_24894);
xor U25003 (N_25003,N_24687,N_24696);
or U25004 (N_25004,N_24700,N_24606);
nand U25005 (N_25005,N_24693,N_24723);
nor U25006 (N_25006,N_24719,N_24845);
or U25007 (N_25007,N_24681,N_24853);
nand U25008 (N_25008,N_24624,N_24858);
nor U25009 (N_25009,N_24764,N_24866);
or U25010 (N_25010,N_24846,N_24601);
and U25011 (N_25011,N_24771,N_24800);
and U25012 (N_25012,N_24727,N_24665);
or U25013 (N_25013,N_24736,N_24787);
nand U25014 (N_25014,N_24899,N_24627);
or U25015 (N_25015,N_24773,N_24645);
and U25016 (N_25016,N_24709,N_24828);
xor U25017 (N_25017,N_24619,N_24755);
nand U25018 (N_25018,N_24615,N_24831);
nand U25019 (N_25019,N_24734,N_24618);
or U25020 (N_25020,N_24768,N_24879);
xnor U25021 (N_25021,N_24769,N_24760);
nand U25022 (N_25022,N_24704,N_24677);
nand U25023 (N_25023,N_24674,N_24650);
xnor U25024 (N_25024,N_24873,N_24842);
xor U25025 (N_25025,N_24893,N_24827);
and U25026 (N_25026,N_24794,N_24651);
or U25027 (N_25027,N_24713,N_24622);
nand U25028 (N_25028,N_24830,N_24811);
xor U25029 (N_25029,N_24705,N_24673);
nor U25030 (N_25030,N_24726,N_24844);
or U25031 (N_25031,N_24740,N_24702);
xnor U25032 (N_25032,N_24712,N_24738);
nand U25033 (N_25033,N_24843,N_24813);
nor U25034 (N_25034,N_24888,N_24706);
xor U25035 (N_25035,N_24821,N_24658);
nand U25036 (N_25036,N_24715,N_24720);
and U25037 (N_25037,N_24714,N_24710);
or U25038 (N_25038,N_24663,N_24772);
nor U25039 (N_25039,N_24660,N_24863);
or U25040 (N_25040,N_24792,N_24668);
xor U25041 (N_25041,N_24864,N_24733);
xnor U25042 (N_25042,N_24731,N_24628);
or U25043 (N_25043,N_24882,N_24784);
xor U25044 (N_25044,N_24889,N_24847);
or U25045 (N_25045,N_24761,N_24629);
and U25046 (N_25046,N_24694,N_24751);
xnor U25047 (N_25047,N_24724,N_24859);
xor U25048 (N_25048,N_24796,N_24646);
xor U25049 (N_25049,N_24803,N_24861);
nand U25050 (N_25050,N_24675,N_24846);
nand U25051 (N_25051,N_24849,N_24768);
xor U25052 (N_25052,N_24757,N_24781);
nand U25053 (N_25053,N_24840,N_24843);
or U25054 (N_25054,N_24658,N_24717);
nor U25055 (N_25055,N_24790,N_24782);
nor U25056 (N_25056,N_24664,N_24812);
or U25057 (N_25057,N_24875,N_24735);
nor U25058 (N_25058,N_24645,N_24842);
or U25059 (N_25059,N_24891,N_24700);
and U25060 (N_25060,N_24608,N_24659);
and U25061 (N_25061,N_24883,N_24708);
xor U25062 (N_25062,N_24668,N_24750);
nor U25063 (N_25063,N_24736,N_24826);
nor U25064 (N_25064,N_24879,N_24737);
nor U25065 (N_25065,N_24864,N_24788);
and U25066 (N_25066,N_24845,N_24898);
or U25067 (N_25067,N_24653,N_24717);
and U25068 (N_25068,N_24852,N_24712);
or U25069 (N_25069,N_24608,N_24706);
nand U25070 (N_25070,N_24838,N_24773);
nand U25071 (N_25071,N_24864,N_24690);
or U25072 (N_25072,N_24761,N_24860);
xor U25073 (N_25073,N_24875,N_24747);
nor U25074 (N_25074,N_24667,N_24700);
nand U25075 (N_25075,N_24894,N_24727);
or U25076 (N_25076,N_24881,N_24830);
and U25077 (N_25077,N_24864,N_24803);
or U25078 (N_25078,N_24639,N_24653);
xor U25079 (N_25079,N_24651,N_24734);
and U25080 (N_25080,N_24852,N_24632);
and U25081 (N_25081,N_24882,N_24761);
and U25082 (N_25082,N_24741,N_24670);
and U25083 (N_25083,N_24696,N_24887);
nor U25084 (N_25084,N_24766,N_24821);
and U25085 (N_25085,N_24742,N_24710);
or U25086 (N_25086,N_24736,N_24854);
or U25087 (N_25087,N_24718,N_24893);
and U25088 (N_25088,N_24646,N_24879);
nand U25089 (N_25089,N_24875,N_24793);
and U25090 (N_25090,N_24751,N_24818);
and U25091 (N_25091,N_24624,N_24781);
or U25092 (N_25092,N_24869,N_24809);
nor U25093 (N_25093,N_24879,N_24704);
xnor U25094 (N_25094,N_24686,N_24786);
or U25095 (N_25095,N_24639,N_24657);
xor U25096 (N_25096,N_24889,N_24864);
or U25097 (N_25097,N_24632,N_24600);
or U25098 (N_25098,N_24758,N_24813);
nand U25099 (N_25099,N_24830,N_24784);
nor U25100 (N_25100,N_24685,N_24731);
nand U25101 (N_25101,N_24710,N_24871);
nand U25102 (N_25102,N_24700,N_24896);
nor U25103 (N_25103,N_24823,N_24793);
nand U25104 (N_25104,N_24878,N_24862);
and U25105 (N_25105,N_24620,N_24845);
nand U25106 (N_25106,N_24786,N_24671);
and U25107 (N_25107,N_24634,N_24762);
nand U25108 (N_25108,N_24675,N_24646);
and U25109 (N_25109,N_24736,N_24883);
nor U25110 (N_25110,N_24778,N_24642);
or U25111 (N_25111,N_24767,N_24602);
xor U25112 (N_25112,N_24808,N_24725);
nand U25113 (N_25113,N_24865,N_24756);
or U25114 (N_25114,N_24887,N_24759);
nor U25115 (N_25115,N_24859,N_24775);
nor U25116 (N_25116,N_24864,N_24867);
nand U25117 (N_25117,N_24890,N_24693);
nand U25118 (N_25118,N_24814,N_24641);
nor U25119 (N_25119,N_24678,N_24890);
nor U25120 (N_25120,N_24621,N_24618);
xnor U25121 (N_25121,N_24612,N_24822);
nor U25122 (N_25122,N_24609,N_24846);
nand U25123 (N_25123,N_24820,N_24696);
nor U25124 (N_25124,N_24774,N_24734);
nor U25125 (N_25125,N_24880,N_24703);
or U25126 (N_25126,N_24895,N_24711);
and U25127 (N_25127,N_24884,N_24737);
nand U25128 (N_25128,N_24645,N_24849);
and U25129 (N_25129,N_24758,N_24757);
xor U25130 (N_25130,N_24687,N_24809);
nor U25131 (N_25131,N_24603,N_24725);
nand U25132 (N_25132,N_24811,N_24665);
xnor U25133 (N_25133,N_24758,N_24645);
and U25134 (N_25134,N_24752,N_24869);
nand U25135 (N_25135,N_24882,N_24602);
nand U25136 (N_25136,N_24867,N_24661);
or U25137 (N_25137,N_24898,N_24689);
or U25138 (N_25138,N_24799,N_24665);
or U25139 (N_25139,N_24812,N_24621);
or U25140 (N_25140,N_24769,N_24772);
and U25141 (N_25141,N_24699,N_24852);
nand U25142 (N_25142,N_24741,N_24685);
nor U25143 (N_25143,N_24849,N_24617);
and U25144 (N_25144,N_24840,N_24763);
xnor U25145 (N_25145,N_24739,N_24711);
nor U25146 (N_25146,N_24891,N_24798);
nand U25147 (N_25147,N_24885,N_24829);
nor U25148 (N_25148,N_24876,N_24602);
or U25149 (N_25149,N_24789,N_24664);
nand U25150 (N_25150,N_24626,N_24804);
and U25151 (N_25151,N_24642,N_24665);
nor U25152 (N_25152,N_24794,N_24620);
nand U25153 (N_25153,N_24746,N_24807);
or U25154 (N_25154,N_24880,N_24638);
and U25155 (N_25155,N_24800,N_24814);
nand U25156 (N_25156,N_24645,N_24627);
nor U25157 (N_25157,N_24748,N_24800);
nand U25158 (N_25158,N_24867,N_24819);
nand U25159 (N_25159,N_24713,N_24780);
xor U25160 (N_25160,N_24617,N_24654);
or U25161 (N_25161,N_24724,N_24852);
or U25162 (N_25162,N_24725,N_24670);
or U25163 (N_25163,N_24690,N_24850);
xor U25164 (N_25164,N_24876,N_24707);
xnor U25165 (N_25165,N_24879,N_24647);
and U25166 (N_25166,N_24817,N_24806);
or U25167 (N_25167,N_24663,N_24758);
or U25168 (N_25168,N_24781,N_24634);
xor U25169 (N_25169,N_24730,N_24749);
or U25170 (N_25170,N_24635,N_24636);
and U25171 (N_25171,N_24603,N_24617);
or U25172 (N_25172,N_24667,N_24785);
or U25173 (N_25173,N_24620,N_24731);
nor U25174 (N_25174,N_24608,N_24796);
or U25175 (N_25175,N_24730,N_24703);
and U25176 (N_25176,N_24850,N_24712);
and U25177 (N_25177,N_24668,N_24838);
or U25178 (N_25178,N_24891,N_24767);
nor U25179 (N_25179,N_24739,N_24722);
xor U25180 (N_25180,N_24861,N_24839);
and U25181 (N_25181,N_24705,N_24600);
xor U25182 (N_25182,N_24812,N_24828);
xor U25183 (N_25183,N_24641,N_24881);
nand U25184 (N_25184,N_24664,N_24753);
or U25185 (N_25185,N_24768,N_24884);
and U25186 (N_25186,N_24852,N_24640);
nor U25187 (N_25187,N_24713,N_24876);
nand U25188 (N_25188,N_24725,N_24840);
and U25189 (N_25189,N_24846,N_24859);
and U25190 (N_25190,N_24657,N_24744);
nor U25191 (N_25191,N_24693,N_24633);
and U25192 (N_25192,N_24691,N_24725);
nand U25193 (N_25193,N_24658,N_24630);
and U25194 (N_25194,N_24885,N_24807);
xor U25195 (N_25195,N_24896,N_24756);
xor U25196 (N_25196,N_24808,N_24692);
or U25197 (N_25197,N_24797,N_24852);
or U25198 (N_25198,N_24784,N_24703);
xnor U25199 (N_25199,N_24666,N_24844);
nor U25200 (N_25200,N_25011,N_24904);
xnor U25201 (N_25201,N_25124,N_25141);
and U25202 (N_25202,N_25000,N_25114);
xor U25203 (N_25203,N_24942,N_24975);
nor U25204 (N_25204,N_25165,N_25123);
nand U25205 (N_25205,N_24932,N_24933);
nor U25206 (N_25206,N_24912,N_25089);
or U25207 (N_25207,N_25031,N_25079);
and U25208 (N_25208,N_25145,N_25016);
or U25209 (N_25209,N_25061,N_25147);
xnor U25210 (N_25210,N_25179,N_25197);
nor U25211 (N_25211,N_25178,N_24999);
or U25212 (N_25212,N_24907,N_25053);
xor U25213 (N_25213,N_25130,N_25188);
nand U25214 (N_25214,N_25126,N_25146);
nor U25215 (N_25215,N_25163,N_24987);
xor U25216 (N_25216,N_25043,N_25054);
or U25217 (N_25217,N_25175,N_24977);
and U25218 (N_25218,N_24952,N_25160);
nor U25219 (N_25219,N_25193,N_24921);
and U25220 (N_25220,N_25148,N_25095);
or U25221 (N_25221,N_25022,N_25083);
nor U25222 (N_25222,N_25009,N_25024);
xnor U25223 (N_25223,N_25021,N_25006);
or U25224 (N_25224,N_25131,N_25030);
nor U25225 (N_25225,N_24973,N_25167);
nor U25226 (N_25226,N_24971,N_25029);
nand U25227 (N_25227,N_24905,N_25045);
xor U25228 (N_25228,N_25080,N_25191);
nand U25229 (N_25229,N_25039,N_25049);
or U25230 (N_25230,N_24949,N_24974);
nand U25231 (N_25231,N_25180,N_25138);
and U25232 (N_25232,N_25102,N_24939);
nand U25233 (N_25233,N_25159,N_24992);
nor U25234 (N_25234,N_25104,N_24919);
and U25235 (N_25235,N_25196,N_25189);
xor U25236 (N_25236,N_24941,N_24981);
nand U25237 (N_25237,N_25065,N_25047);
xor U25238 (N_25238,N_24923,N_25170);
xnor U25239 (N_25239,N_25135,N_24958);
nand U25240 (N_25240,N_25062,N_25055);
xnor U25241 (N_25241,N_24968,N_25040);
and U25242 (N_25242,N_24994,N_25121);
nand U25243 (N_25243,N_24926,N_25142);
and U25244 (N_25244,N_25119,N_24929);
nand U25245 (N_25245,N_24931,N_25044);
nor U25246 (N_25246,N_25017,N_25073);
nand U25247 (N_25247,N_25183,N_25052);
xnor U25248 (N_25248,N_25105,N_24947);
nor U25249 (N_25249,N_24908,N_25036);
or U25250 (N_25250,N_24979,N_24950);
nand U25251 (N_25251,N_25046,N_25115);
and U25252 (N_25252,N_24946,N_25032);
nor U25253 (N_25253,N_25100,N_25087);
or U25254 (N_25254,N_24944,N_25139);
nand U25255 (N_25255,N_24997,N_25056);
nand U25256 (N_25256,N_25051,N_25068);
xnor U25257 (N_25257,N_25075,N_24988);
nor U25258 (N_25258,N_24938,N_24901);
or U25259 (N_25259,N_24995,N_24991);
xor U25260 (N_25260,N_24927,N_25008);
or U25261 (N_25261,N_24903,N_24959);
and U25262 (N_25262,N_24928,N_24996);
xnor U25263 (N_25263,N_24960,N_25005);
and U25264 (N_25264,N_25158,N_24961);
nor U25265 (N_25265,N_25195,N_25125);
nand U25266 (N_25266,N_25199,N_25077);
and U25267 (N_25267,N_25185,N_25157);
nand U25268 (N_25268,N_25042,N_25085);
and U25269 (N_25269,N_25001,N_25111);
or U25270 (N_25270,N_25136,N_25113);
nor U25271 (N_25271,N_24980,N_25152);
nor U25272 (N_25272,N_24955,N_24915);
and U25273 (N_25273,N_24918,N_24993);
and U25274 (N_25274,N_25133,N_24906);
nand U25275 (N_25275,N_25103,N_24948);
nand U25276 (N_25276,N_25174,N_24940);
nor U25277 (N_25277,N_24910,N_24983);
or U25278 (N_25278,N_24976,N_25122);
nand U25279 (N_25279,N_24900,N_25164);
nand U25280 (N_25280,N_25025,N_24925);
or U25281 (N_25281,N_25020,N_25093);
nand U25282 (N_25282,N_25059,N_25086);
nor U25283 (N_25283,N_25186,N_24913);
and U25284 (N_25284,N_25023,N_24902);
and U25285 (N_25285,N_24962,N_24916);
and U25286 (N_25286,N_24922,N_25074);
nand U25287 (N_25287,N_25067,N_24937);
nor U25288 (N_25288,N_24943,N_25127);
nand U25289 (N_25289,N_25019,N_25190);
nand U25290 (N_25290,N_25162,N_24989);
nor U25291 (N_25291,N_25140,N_25137);
xor U25292 (N_25292,N_24954,N_25066);
and U25293 (N_25293,N_24970,N_24911);
and U25294 (N_25294,N_25110,N_24951);
or U25295 (N_25295,N_25014,N_25128);
nand U25296 (N_25296,N_25120,N_24909);
or U25297 (N_25297,N_25144,N_25117);
nor U25298 (N_25298,N_24936,N_25172);
nand U25299 (N_25299,N_25028,N_25081);
or U25300 (N_25300,N_25088,N_25098);
nand U25301 (N_25301,N_25058,N_25091);
xnor U25302 (N_25302,N_25150,N_24945);
nor U25303 (N_25303,N_24953,N_25057);
and U25304 (N_25304,N_24956,N_25177);
nand U25305 (N_25305,N_24967,N_25154);
nor U25306 (N_25306,N_25048,N_24985);
nor U25307 (N_25307,N_25004,N_24998);
nor U25308 (N_25308,N_25050,N_25026);
or U25309 (N_25309,N_25129,N_25101);
and U25310 (N_25310,N_25033,N_25099);
xnor U25311 (N_25311,N_25176,N_24924);
xnor U25312 (N_25312,N_25096,N_25108);
or U25313 (N_25313,N_25038,N_24969);
nand U25314 (N_25314,N_25156,N_24964);
and U25315 (N_25315,N_25082,N_25034);
and U25316 (N_25316,N_24978,N_25076);
and U25317 (N_25317,N_25002,N_24914);
nand U25318 (N_25318,N_25007,N_24965);
nand U25319 (N_25319,N_25060,N_25112);
or U25320 (N_25320,N_25041,N_25192);
and U25321 (N_25321,N_25181,N_24920);
nor U25322 (N_25322,N_24966,N_25143);
nand U25323 (N_25323,N_24972,N_25035);
xnor U25324 (N_25324,N_24986,N_25169);
xor U25325 (N_25325,N_25187,N_24934);
xor U25326 (N_25326,N_25090,N_25171);
or U25327 (N_25327,N_25149,N_25027);
and U25328 (N_25328,N_25153,N_25010);
and U25329 (N_25329,N_24917,N_25018);
nor U25330 (N_25330,N_25109,N_25168);
nor U25331 (N_25331,N_25078,N_25012);
or U25332 (N_25332,N_25184,N_25069);
xnor U25333 (N_25333,N_25092,N_24984);
nor U25334 (N_25334,N_25015,N_25118);
xor U25335 (N_25335,N_25070,N_25084);
or U25336 (N_25336,N_25072,N_24957);
nand U25337 (N_25337,N_25161,N_24963);
or U25338 (N_25338,N_25063,N_25198);
or U25339 (N_25339,N_25107,N_24982);
nor U25340 (N_25340,N_25037,N_25071);
or U25341 (N_25341,N_24990,N_25013);
nor U25342 (N_25342,N_24935,N_24930);
nand U25343 (N_25343,N_25064,N_25116);
xnor U25344 (N_25344,N_25182,N_25097);
nand U25345 (N_25345,N_25155,N_25134);
nor U25346 (N_25346,N_25166,N_25094);
or U25347 (N_25347,N_25151,N_25132);
nand U25348 (N_25348,N_25003,N_25173);
nor U25349 (N_25349,N_25106,N_25194);
and U25350 (N_25350,N_25159,N_25026);
xnor U25351 (N_25351,N_24968,N_25055);
and U25352 (N_25352,N_25152,N_24968);
nor U25353 (N_25353,N_24984,N_25114);
and U25354 (N_25354,N_24946,N_25005);
and U25355 (N_25355,N_25069,N_25077);
or U25356 (N_25356,N_24970,N_25047);
xor U25357 (N_25357,N_24968,N_25091);
nand U25358 (N_25358,N_25047,N_24916);
xor U25359 (N_25359,N_24911,N_25023);
xnor U25360 (N_25360,N_24999,N_25025);
xnor U25361 (N_25361,N_24968,N_25124);
nor U25362 (N_25362,N_24989,N_25085);
or U25363 (N_25363,N_25006,N_24975);
and U25364 (N_25364,N_24922,N_24908);
or U25365 (N_25365,N_25176,N_25119);
and U25366 (N_25366,N_24965,N_25105);
xor U25367 (N_25367,N_25088,N_25130);
or U25368 (N_25368,N_25081,N_25063);
nand U25369 (N_25369,N_25109,N_25173);
and U25370 (N_25370,N_25072,N_24975);
xnor U25371 (N_25371,N_25118,N_25031);
xnor U25372 (N_25372,N_25061,N_25024);
nor U25373 (N_25373,N_24981,N_25075);
and U25374 (N_25374,N_25179,N_25091);
xnor U25375 (N_25375,N_24948,N_25166);
xor U25376 (N_25376,N_25011,N_25131);
nor U25377 (N_25377,N_25038,N_24970);
or U25378 (N_25378,N_25049,N_24962);
xnor U25379 (N_25379,N_25049,N_24915);
or U25380 (N_25380,N_25015,N_25040);
xor U25381 (N_25381,N_24982,N_24991);
nand U25382 (N_25382,N_25199,N_25031);
nor U25383 (N_25383,N_25104,N_25193);
xnor U25384 (N_25384,N_25131,N_25084);
nor U25385 (N_25385,N_25149,N_25141);
xnor U25386 (N_25386,N_24915,N_24920);
or U25387 (N_25387,N_25142,N_25131);
xnor U25388 (N_25388,N_24949,N_25093);
nand U25389 (N_25389,N_25095,N_25018);
xor U25390 (N_25390,N_25107,N_25119);
and U25391 (N_25391,N_25163,N_25021);
or U25392 (N_25392,N_25127,N_25068);
or U25393 (N_25393,N_24984,N_25167);
nor U25394 (N_25394,N_24965,N_25069);
xnor U25395 (N_25395,N_25015,N_25045);
and U25396 (N_25396,N_25176,N_25099);
and U25397 (N_25397,N_25102,N_25005);
and U25398 (N_25398,N_24945,N_24979);
or U25399 (N_25399,N_24996,N_24969);
nor U25400 (N_25400,N_25132,N_24907);
or U25401 (N_25401,N_25199,N_25009);
nor U25402 (N_25402,N_25199,N_24952);
and U25403 (N_25403,N_25133,N_25058);
or U25404 (N_25404,N_25037,N_25074);
and U25405 (N_25405,N_25183,N_25175);
nand U25406 (N_25406,N_25097,N_24943);
xor U25407 (N_25407,N_25042,N_24900);
nand U25408 (N_25408,N_25041,N_25055);
nor U25409 (N_25409,N_25177,N_25181);
and U25410 (N_25410,N_25097,N_25130);
nor U25411 (N_25411,N_24940,N_25021);
or U25412 (N_25412,N_24963,N_25024);
or U25413 (N_25413,N_24935,N_25176);
nor U25414 (N_25414,N_25071,N_24928);
nand U25415 (N_25415,N_25142,N_25174);
nor U25416 (N_25416,N_24944,N_25049);
nor U25417 (N_25417,N_25017,N_24903);
xnor U25418 (N_25418,N_24901,N_24956);
and U25419 (N_25419,N_25037,N_25164);
xnor U25420 (N_25420,N_25188,N_25156);
xnor U25421 (N_25421,N_25196,N_24992);
nor U25422 (N_25422,N_24950,N_25199);
nor U25423 (N_25423,N_24946,N_24934);
nand U25424 (N_25424,N_24924,N_25143);
nor U25425 (N_25425,N_24939,N_24969);
xor U25426 (N_25426,N_25166,N_24941);
nand U25427 (N_25427,N_24970,N_24999);
or U25428 (N_25428,N_25064,N_25102);
nand U25429 (N_25429,N_25084,N_24985);
and U25430 (N_25430,N_25097,N_24997);
xor U25431 (N_25431,N_24935,N_24970);
or U25432 (N_25432,N_25036,N_25093);
nor U25433 (N_25433,N_24910,N_25022);
nor U25434 (N_25434,N_25184,N_25049);
xor U25435 (N_25435,N_25123,N_25035);
nor U25436 (N_25436,N_25140,N_25116);
xor U25437 (N_25437,N_25044,N_25177);
or U25438 (N_25438,N_25008,N_25153);
nor U25439 (N_25439,N_24962,N_25121);
xor U25440 (N_25440,N_24910,N_25197);
or U25441 (N_25441,N_25041,N_25163);
nand U25442 (N_25442,N_25127,N_25064);
xor U25443 (N_25443,N_24941,N_25012);
or U25444 (N_25444,N_25041,N_25190);
nand U25445 (N_25445,N_25181,N_24998);
nand U25446 (N_25446,N_24913,N_25143);
or U25447 (N_25447,N_24932,N_25010);
or U25448 (N_25448,N_25159,N_24944);
and U25449 (N_25449,N_25107,N_24964);
or U25450 (N_25450,N_24945,N_25039);
xnor U25451 (N_25451,N_24974,N_25181);
and U25452 (N_25452,N_25124,N_25068);
xor U25453 (N_25453,N_24923,N_25186);
nand U25454 (N_25454,N_24952,N_24949);
and U25455 (N_25455,N_25169,N_24913);
and U25456 (N_25456,N_24999,N_25075);
nand U25457 (N_25457,N_24905,N_24935);
or U25458 (N_25458,N_24938,N_25109);
or U25459 (N_25459,N_25030,N_25129);
nand U25460 (N_25460,N_24916,N_25122);
and U25461 (N_25461,N_25001,N_25005);
nand U25462 (N_25462,N_25071,N_25018);
and U25463 (N_25463,N_24961,N_24946);
xnor U25464 (N_25464,N_24904,N_24973);
xnor U25465 (N_25465,N_25154,N_25184);
and U25466 (N_25466,N_25128,N_25040);
xnor U25467 (N_25467,N_25045,N_25111);
xnor U25468 (N_25468,N_25161,N_24986);
nand U25469 (N_25469,N_25080,N_25156);
and U25470 (N_25470,N_24991,N_24924);
nor U25471 (N_25471,N_24948,N_25122);
and U25472 (N_25472,N_25180,N_24993);
xor U25473 (N_25473,N_25083,N_25177);
xnor U25474 (N_25474,N_25050,N_24900);
nand U25475 (N_25475,N_25185,N_24997);
nor U25476 (N_25476,N_24981,N_24962);
and U25477 (N_25477,N_25080,N_25195);
nand U25478 (N_25478,N_25011,N_25023);
or U25479 (N_25479,N_25026,N_25196);
or U25480 (N_25480,N_25004,N_25123);
and U25481 (N_25481,N_24968,N_25199);
and U25482 (N_25482,N_25041,N_25177);
or U25483 (N_25483,N_24996,N_25028);
nor U25484 (N_25484,N_24916,N_24998);
nor U25485 (N_25485,N_25175,N_25061);
or U25486 (N_25486,N_25113,N_25174);
nor U25487 (N_25487,N_25074,N_25039);
nor U25488 (N_25488,N_25087,N_25052);
nor U25489 (N_25489,N_25098,N_25159);
nand U25490 (N_25490,N_25192,N_24985);
nand U25491 (N_25491,N_25032,N_25118);
nor U25492 (N_25492,N_25052,N_24934);
or U25493 (N_25493,N_25132,N_25050);
or U25494 (N_25494,N_25039,N_25146);
or U25495 (N_25495,N_25185,N_24965);
xnor U25496 (N_25496,N_25069,N_25109);
nand U25497 (N_25497,N_25018,N_25023);
nor U25498 (N_25498,N_25188,N_25133);
or U25499 (N_25499,N_25069,N_25002);
xnor U25500 (N_25500,N_25390,N_25484);
xor U25501 (N_25501,N_25316,N_25346);
or U25502 (N_25502,N_25419,N_25460);
nand U25503 (N_25503,N_25291,N_25481);
and U25504 (N_25504,N_25221,N_25278);
nand U25505 (N_25505,N_25360,N_25332);
and U25506 (N_25506,N_25434,N_25226);
and U25507 (N_25507,N_25229,N_25435);
nand U25508 (N_25508,N_25334,N_25279);
nor U25509 (N_25509,N_25374,N_25282);
nor U25510 (N_25510,N_25391,N_25202);
nor U25511 (N_25511,N_25248,N_25305);
or U25512 (N_25512,N_25265,N_25285);
nor U25513 (N_25513,N_25459,N_25491);
nand U25514 (N_25514,N_25228,N_25274);
or U25515 (N_25515,N_25362,N_25350);
nand U25516 (N_25516,N_25313,N_25338);
and U25517 (N_25517,N_25284,N_25406);
nor U25518 (N_25518,N_25424,N_25372);
or U25519 (N_25519,N_25428,N_25335);
and U25520 (N_25520,N_25266,N_25247);
nand U25521 (N_25521,N_25482,N_25369);
and U25522 (N_25522,N_25306,N_25377);
xor U25523 (N_25523,N_25402,N_25487);
nand U25524 (N_25524,N_25272,N_25463);
nor U25525 (N_25525,N_25280,N_25364);
xnor U25526 (N_25526,N_25498,N_25336);
nor U25527 (N_25527,N_25398,N_25296);
nand U25528 (N_25528,N_25474,N_25301);
and U25529 (N_25529,N_25339,N_25210);
nor U25530 (N_25530,N_25351,N_25212);
nand U25531 (N_25531,N_25224,N_25251);
or U25532 (N_25532,N_25277,N_25241);
nor U25533 (N_25533,N_25456,N_25206);
xnor U25534 (N_25534,N_25380,N_25401);
and U25535 (N_25535,N_25250,N_25264);
nand U25536 (N_25536,N_25384,N_25227);
nor U25537 (N_25537,N_25348,N_25497);
nor U25538 (N_25538,N_25433,N_25394);
and U25539 (N_25539,N_25446,N_25381);
nand U25540 (N_25540,N_25458,N_25337);
xor U25541 (N_25541,N_25492,N_25326);
or U25542 (N_25542,N_25449,N_25344);
and U25543 (N_25543,N_25421,N_25440);
or U25544 (N_25544,N_25499,N_25445);
and U25545 (N_25545,N_25429,N_25235);
xnor U25546 (N_25546,N_25341,N_25475);
xor U25547 (N_25547,N_25464,N_25246);
and U25548 (N_25548,N_25415,N_25454);
and U25549 (N_25549,N_25476,N_25447);
xor U25550 (N_25550,N_25437,N_25414);
and U25551 (N_25551,N_25349,N_25207);
and U25552 (N_25552,N_25363,N_25438);
and U25553 (N_25553,N_25310,N_25411);
or U25554 (N_25554,N_25366,N_25315);
and U25555 (N_25555,N_25451,N_25404);
and U25556 (N_25556,N_25288,N_25397);
and U25557 (N_25557,N_25214,N_25238);
nand U25558 (N_25558,N_25443,N_25312);
nand U25559 (N_25559,N_25358,N_25269);
nand U25560 (N_25560,N_25483,N_25489);
xor U25561 (N_25561,N_25299,N_25478);
or U25562 (N_25562,N_25289,N_25300);
nor U25563 (N_25563,N_25262,N_25263);
or U25564 (N_25564,N_25455,N_25383);
or U25565 (N_25565,N_25409,N_25314);
or U25566 (N_25566,N_25450,N_25457);
nand U25567 (N_25567,N_25392,N_25473);
or U25568 (N_25568,N_25201,N_25468);
xor U25569 (N_25569,N_25254,N_25295);
and U25570 (N_25570,N_25209,N_25425);
nand U25571 (N_25571,N_25304,N_25432);
or U25572 (N_25572,N_25410,N_25245);
nand U25573 (N_25573,N_25333,N_25215);
nand U25574 (N_25574,N_25239,N_25452);
xnor U25575 (N_25575,N_25240,N_25340);
xnor U25576 (N_25576,N_25396,N_25387);
nand U25577 (N_25577,N_25298,N_25273);
xor U25578 (N_25578,N_25386,N_25426);
or U25579 (N_25579,N_25236,N_25343);
or U25580 (N_25580,N_25393,N_25242);
or U25581 (N_25581,N_25311,N_25399);
xnor U25582 (N_25582,N_25423,N_25328);
and U25583 (N_25583,N_25308,N_25297);
nand U25584 (N_25584,N_25294,N_25268);
or U25585 (N_25585,N_25234,N_25453);
and U25586 (N_25586,N_25418,N_25237);
nand U25587 (N_25587,N_25490,N_25361);
and U25588 (N_25588,N_25325,N_25462);
or U25589 (N_25589,N_25309,N_25261);
nor U25590 (N_25590,N_25353,N_25480);
or U25591 (N_25591,N_25318,N_25412);
xor U25592 (N_25592,N_25253,N_25370);
or U25593 (N_25593,N_25467,N_25417);
nor U25594 (N_25594,N_25292,N_25407);
nand U25595 (N_25595,N_25231,N_25448);
nand U25596 (N_25596,N_25494,N_25485);
and U25597 (N_25597,N_25439,N_25472);
nor U25598 (N_25598,N_25222,N_25400);
and U25599 (N_25599,N_25465,N_25267);
xnor U25600 (N_25600,N_25357,N_25243);
or U25601 (N_25601,N_25217,N_25287);
xnor U25602 (N_25602,N_25249,N_25389);
nor U25603 (N_25603,N_25302,N_25225);
or U25604 (N_25604,N_25200,N_25368);
nand U25605 (N_25605,N_25211,N_25469);
or U25606 (N_25606,N_25470,N_25359);
and U25607 (N_25607,N_25271,N_25365);
or U25608 (N_25608,N_25307,N_25208);
xor U25609 (N_25609,N_25422,N_25255);
nand U25610 (N_25610,N_25233,N_25218);
nand U25611 (N_25611,N_25371,N_25223);
or U25612 (N_25612,N_25408,N_25388);
xnor U25613 (N_25613,N_25260,N_25431);
and U25614 (N_25614,N_25303,N_25352);
nor U25615 (N_25615,N_25427,N_25347);
and U25616 (N_25616,N_25354,N_25382);
nor U25617 (N_25617,N_25441,N_25493);
nor U25618 (N_25618,N_25376,N_25430);
and U25619 (N_25619,N_25461,N_25342);
nor U25620 (N_25620,N_25356,N_25436);
or U25621 (N_25621,N_25495,N_25275);
and U25622 (N_25622,N_25259,N_25252);
xnor U25623 (N_25623,N_25444,N_25323);
and U25624 (N_25624,N_25216,N_25324);
or U25625 (N_25625,N_25220,N_25230);
nor U25626 (N_25626,N_25442,N_25276);
xnor U25627 (N_25627,N_25317,N_25355);
nand U25628 (N_25628,N_25258,N_25403);
and U25629 (N_25629,N_25379,N_25319);
nor U25630 (N_25630,N_25486,N_25256);
xor U25631 (N_25631,N_25488,N_25203);
nand U25632 (N_25632,N_25321,N_25345);
nand U25633 (N_25633,N_25283,N_25244);
or U25634 (N_25634,N_25479,N_25331);
nand U25635 (N_25635,N_25413,N_25322);
nand U25636 (N_25636,N_25213,N_25373);
and U25637 (N_25637,N_25320,N_25385);
and U25638 (N_25638,N_25205,N_25466);
and U25639 (N_25639,N_25293,N_25286);
xnor U25640 (N_25640,N_25416,N_25270);
and U25641 (N_25641,N_25330,N_25375);
or U25642 (N_25642,N_25204,N_25378);
or U25643 (N_25643,N_25290,N_25329);
and U25644 (N_25644,N_25281,N_25496);
and U25645 (N_25645,N_25232,N_25367);
xor U25646 (N_25646,N_25327,N_25420);
and U25647 (N_25647,N_25257,N_25219);
xnor U25648 (N_25648,N_25471,N_25405);
or U25649 (N_25649,N_25395,N_25477);
and U25650 (N_25650,N_25266,N_25496);
or U25651 (N_25651,N_25218,N_25202);
nor U25652 (N_25652,N_25267,N_25358);
xor U25653 (N_25653,N_25434,N_25265);
or U25654 (N_25654,N_25434,N_25243);
or U25655 (N_25655,N_25451,N_25237);
and U25656 (N_25656,N_25452,N_25409);
nand U25657 (N_25657,N_25444,N_25358);
and U25658 (N_25658,N_25343,N_25452);
and U25659 (N_25659,N_25324,N_25450);
and U25660 (N_25660,N_25410,N_25431);
xnor U25661 (N_25661,N_25395,N_25497);
or U25662 (N_25662,N_25319,N_25307);
nor U25663 (N_25663,N_25274,N_25324);
nor U25664 (N_25664,N_25238,N_25233);
nand U25665 (N_25665,N_25448,N_25243);
xor U25666 (N_25666,N_25488,N_25439);
and U25667 (N_25667,N_25304,N_25228);
or U25668 (N_25668,N_25386,N_25318);
xor U25669 (N_25669,N_25201,N_25297);
nor U25670 (N_25670,N_25384,N_25228);
or U25671 (N_25671,N_25456,N_25409);
or U25672 (N_25672,N_25328,N_25480);
xnor U25673 (N_25673,N_25300,N_25299);
nor U25674 (N_25674,N_25390,N_25480);
nand U25675 (N_25675,N_25366,N_25392);
and U25676 (N_25676,N_25408,N_25346);
or U25677 (N_25677,N_25375,N_25349);
nand U25678 (N_25678,N_25389,N_25395);
xor U25679 (N_25679,N_25448,N_25245);
nor U25680 (N_25680,N_25478,N_25348);
xnor U25681 (N_25681,N_25255,N_25315);
xnor U25682 (N_25682,N_25495,N_25201);
nand U25683 (N_25683,N_25378,N_25247);
nand U25684 (N_25684,N_25397,N_25269);
and U25685 (N_25685,N_25394,N_25344);
nor U25686 (N_25686,N_25469,N_25414);
or U25687 (N_25687,N_25275,N_25259);
and U25688 (N_25688,N_25467,N_25392);
xnor U25689 (N_25689,N_25311,N_25428);
xnor U25690 (N_25690,N_25243,N_25298);
and U25691 (N_25691,N_25223,N_25328);
nand U25692 (N_25692,N_25423,N_25333);
xnor U25693 (N_25693,N_25426,N_25337);
or U25694 (N_25694,N_25255,N_25440);
xor U25695 (N_25695,N_25303,N_25479);
or U25696 (N_25696,N_25319,N_25399);
nand U25697 (N_25697,N_25406,N_25340);
nand U25698 (N_25698,N_25236,N_25238);
nand U25699 (N_25699,N_25363,N_25462);
and U25700 (N_25700,N_25447,N_25462);
nand U25701 (N_25701,N_25201,N_25444);
xor U25702 (N_25702,N_25280,N_25415);
nor U25703 (N_25703,N_25482,N_25320);
nand U25704 (N_25704,N_25442,N_25391);
and U25705 (N_25705,N_25258,N_25431);
nand U25706 (N_25706,N_25253,N_25367);
xor U25707 (N_25707,N_25438,N_25263);
and U25708 (N_25708,N_25408,N_25321);
and U25709 (N_25709,N_25252,N_25490);
nand U25710 (N_25710,N_25271,N_25230);
nand U25711 (N_25711,N_25358,N_25370);
or U25712 (N_25712,N_25410,N_25393);
nand U25713 (N_25713,N_25292,N_25397);
xnor U25714 (N_25714,N_25457,N_25403);
nor U25715 (N_25715,N_25402,N_25202);
or U25716 (N_25716,N_25473,N_25432);
nand U25717 (N_25717,N_25395,N_25415);
xor U25718 (N_25718,N_25338,N_25230);
or U25719 (N_25719,N_25223,N_25489);
and U25720 (N_25720,N_25343,N_25495);
nor U25721 (N_25721,N_25221,N_25304);
nor U25722 (N_25722,N_25315,N_25378);
xnor U25723 (N_25723,N_25492,N_25231);
or U25724 (N_25724,N_25232,N_25227);
xor U25725 (N_25725,N_25465,N_25264);
and U25726 (N_25726,N_25286,N_25371);
xor U25727 (N_25727,N_25314,N_25365);
nor U25728 (N_25728,N_25272,N_25273);
nor U25729 (N_25729,N_25253,N_25493);
xor U25730 (N_25730,N_25490,N_25311);
nand U25731 (N_25731,N_25470,N_25246);
and U25732 (N_25732,N_25467,N_25361);
and U25733 (N_25733,N_25440,N_25446);
or U25734 (N_25734,N_25227,N_25238);
or U25735 (N_25735,N_25244,N_25437);
nand U25736 (N_25736,N_25233,N_25258);
and U25737 (N_25737,N_25250,N_25303);
and U25738 (N_25738,N_25447,N_25458);
nand U25739 (N_25739,N_25448,N_25204);
and U25740 (N_25740,N_25417,N_25380);
or U25741 (N_25741,N_25373,N_25252);
and U25742 (N_25742,N_25222,N_25381);
nor U25743 (N_25743,N_25335,N_25208);
nor U25744 (N_25744,N_25250,N_25419);
nand U25745 (N_25745,N_25388,N_25317);
xnor U25746 (N_25746,N_25317,N_25365);
nand U25747 (N_25747,N_25308,N_25338);
or U25748 (N_25748,N_25439,N_25204);
nor U25749 (N_25749,N_25347,N_25373);
and U25750 (N_25750,N_25456,N_25298);
nand U25751 (N_25751,N_25229,N_25426);
and U25752 (N_25752,N_25468,N_25358);
and U25753 (N_25753,N_25236,N_25248);
or U25754 (N_25754,N_25331,N_25402);
nand U25755 (N_25755,N_25441,N_25431);
or U25756 (N_25756,N_25201,N_25342);
nand U25757 (N_25757,N_25487,N_25282);
or U25758 (N_25758,N_25393,N_25459);
xnor U25759 (N_25759,N_25341,N_25226);
or U25760 (N_25760,N_25403,N_25312);
nor U25761 (N_25761,N_25252,N_25265);
and U25762 (N_25762,N_25277,N_25254);
or U25763 (N_25763,N_25439,N_25272);
nand U25764 (N_25764,N_25262,N_25479);
xor U25765 (N_25765,N_25426,N_25334);
and U25766 (N_25766,N_25435,N_25406);
nor U25767 (N_25767,N_25458,N_25339);
or U25768 (N_25768,N_25356,N_25393);
or U25769 (N_25769,N_25451,N_25481);
or U25770 (N_25770,N_25215,N_25453);
or U25771 (N_25771,N_25474,N_25257);
nand U25772 (N_25772,N_25383,N_25484);
nor U25773 (N_25773,N_25496,N_25291);
nand U25774 (N_25774,N_25347,N_25489);
xor U25775 (N_25775,N_25367,N_25252);
nor U25776 (N_25776,N_25403,N_25293);
and U25777 (N_25777,N_25424,N_25359);
nand U25778 (N_25778,N_25245,N_25300);
or U25779 (N_25779,N_25465,N_25263);
xnor U25780 (N_25780,N_25406,N_25261);
and U25781 (N_25781,N_25291,N_25323);
xor U25782 (N_25782,N_25246,N_25298);
and U25783 (N_25783,N_25342,N_25480);
xor U25784 (N_25784,N_25383,N_25354);
and U25785 (N_25785,N_25438,N_25471);
and U25786 (N_25786,N_25297,N_25341);
nand U25787 (N_25787,N_25231,N_25365);
nor U25788 (N_25788,N_25392,N_25406);
and U25789 (N_25789,N_25349,N_25422);
xnor U25790 (N_25790,N_25380,N_25416);
and U25791 (N_25791,N_25346,N_25402);
nand U25792 (N_25792,N_25444,N_25411);
and U25793 (N_25793,N_25383,N_25288);
and U25794 (N_25794,N_25304,N_25435);
and U25795 (N_25795,N_25472,N_25396);
nor U25796 (N_25796,N_25349,N_25356);
xnor U25797 (N_25797,N_25435,N_25454);
and U25798 (N_25798,N_25253,N_25433);
or U25799 (N_25799,N_25202,N_25420);
nand U25800 (N_25800,N_25771,N_25774);
xor U25801 (N_25801,N_25672,N_25570);
or U25802 (N_25802,N_25562,N_25612);
and U25803 (N_25803,N_25662,N_25615);
and U25804 (N_25804,N_25682,N_25544);
xor U25805 (N_25805,N_25538,N_25709);
or U25806 (N_25806,N_25704,N_25553);
and U25807 (N_25807,N_25727,N_25623);
nand U25808 (N_25808,N_25724,N_25658);
or U25809 (N_25809,N_25655,N_25798);
nor U25810 (N_25810,N_25632,N_25780);
xor U25811 (N_25811,N_25740,N_25669);
nor U25812 (N_25812,N_25734,N_25700);
or U25813 (N_25813,N_25522,N_25576);
nor U25814 (N_25814,N_25664,N_25679);
nor U25815 (N_25815,N_25715,N_25573);
xor U25816 (N_25816,N_25775,N_25536);
or U25817 (N_25817,N_25566,N_25581);
xor U25818 (N_25818,N_25527,N_25747);
xnor U25819 (N_25819,N_25557,N_25512);
and U25820 (N_25820,N_25794,N_25607);
and U25821 (N_25821,N_25680,N_25735);
or U25822 (N_25822,N_25530,N_25706);
xor U25823 (N_25823,N_25641,N_25508);
or U25824 (N_25824,N_25653,N_25759);
nand U25825 (N_25825,N_25693,N_25502);
xnor U25826 (N_25826,N_25541,N_25587);
nand U25827 (N_25827,N_25618,N_25764);
xnor U25828 (N_25828,N_25796,N_25501);
nor U25829 (N_25829,N_25614,N_25517);
xnor U25830 (N_25830,N_25546,N_25762);
and U25831 (N_25831,N_25599,N_25580);
and U25832 (N_25832,N_25554,N_25627);
xnor U25833 (N_25833,N_25579,N_25716);
xor U25834 (N_25834,N_25500,N_25635);
xnor U25835 (N_25835,N_25751,N_25742);
or U25836 (N_25836,N_25708,N_25630);
or U25837 (N_25837,N_25650,N_25617);
nor U25838 (N_25838,N_25531,N_25763);
nand U25839 (N_25839,N_25535,N_25616);
or U25840 (N_25840,N_25745,N_25737);
xor U25841 (N_25841,N_25528,N_25703);
and U25842 (N_25842,N_25564,N_25783);
nor U25843 (N_25843,N_25729,N_25671);
or U25844 (N_25844,N_25768,N_25567);
and U25845 (N_25845,N_25743,N_25721);
nor U25846 (N_25846,N_25519,N_25640);
or U25847 (N_25847,N_25521,N_25651);
xor U25848 (N_25848,N_25789,N_25514);
nor U25849 (N_25849,N_25516,N_25643);
xor U25850 (N_25850,N_25565,N_25620);
or U25851 (N_25851,N_25539,N_25791);
nand U25852 (N_25852,N_25758,N_25639);
xnor U25853 (N_25853,N_25788,N_25532);
xor U25854 (N_25854,N_25606,N_25634);
or U25855 (N_25855,N_25660,N_25540);
or U25856 (N_25856,N_25642,N_25622);
xnor U25857 (N_25857,N_25547,N_25718);
nor U25858 (N_25858,N_25592,N_25585);
xor U25859 (N_25859,N_25707,N_25761);
or U25860 (N_25860,N_25503,N_25636);
xor U25861 (N_25861,N_25550,N_25736);
nor U25862 (N_25862,N_25694,N_25504);
nor U25863 (N_25863,N_25697,N_25558);
and U25864 (N_25864,N_25593,N_25604);
xnor U25865 (N_25865,N_25510,N_25511);
xnor U25866 (N_25866,N_25732,N_25770);
nor U25867 (N_25867,N_25760,N_25657);
and U25868 (N_25868,N_25730,N_25600);
and U25869 (N_25869,N_25792,N_25781);
or U25870 (N_25870,N_25691,N_25624);
nor U25871 (N_25871,N_25722,N_25506);
or U25872 (N_25872,N_25569,N_25690);
and U25873 (N_25873,N_25799,N_25583);
and U25874 (N_25874,N_25526,N_25685);
nor U25875 (N_25875,N_25534,N_25552);
nor U25876 (N_25876,N_25711,N_25753);
and U25877 (N_25877,N_25563,N_25505);
nor U25878 (N_25878,N_25601,N_25572);
xnor U25879 (N_25879,N_25668,N_25712);
or U25880 (N_25880,N_25665,N_25754);
xnor U25881 (N_25881,N_25752,N_25611);
xnor U25882 (N_25882,N_25595,N_25688);
and U25883 (N_25883,N_25725,N_25701);
xor U25884 (N_25884,N_25790,N_25686);
xnor U25885 (N_25885,N_25756,N_25598);
and U25886 (N_25886,N_25594,N_25631);
or U25887 (N_25887,N_25678,N_25705);
nor U25888 (N_25888,N_25741,N_25757);
xor U25889 (N_25889,N_25681,N_25551);
and U25890 (N_25890,N_25625,N_25591);
xor U25891 (N_25891,N_25596,N_25777);
nand U25892 (N_25892,N_25513,N_25561);
nand U25893 (N_25893,N_25590,N_25670);
nand U25894 (N_25894,N_25529,N_25609);
nand U25895 (N_25895,N_25648,N_25676);
nand U25896 (N_25896,N_25548,N_25793);
xnor U25897 (N_25897,N_25755,N_25786);
and U25898 (N_25898,N_25637,N_25647);
nor U25899 (N_25899,N_25602,N_25738);
nand U25900 (N_25900,N_25785,N_25698);
and U25901 (N_25901,N_25795,N_25537);
xor U25902 (N_25902,N_25677,N_25723);
xnor U25903 (N_25903,N_25719,N_25556);
and U25904 (N_25904,N_25767,N_25578);
and U25905 (N_25905,N_25577,N_25610);
and U25906 (N_25906,N_25520,N_25689);
and U25907 (N_25907,N_25597,N_25710);
nor U25908 (N_25908,N_25649,N_25518);
nor U25909 (N_25909,N_25714,N_25589);
nor U25910 (N_25910,N_25525,N_25524);
nand U25911 (N_25911,N_25568,N_25582);
nor U25912 (N_25912,N_25720,N_25750);
xor U25913 (N_25913,N_25687,N_25772);
xor U25914 (N_25914,N_25717,N_25666);
xor U25915 (N_25915,N_25702,N_25731);
xnor U25916 (N_25916,N_25739,N_25748);
and U25917 (N_25917,N_25695,N_25559);
nor U25918 (N_25918,N_25608,N_25773);
or U25919 (N_25919,N_25613,N_25683);
and U25920 (N_25920,N_25654,N_25543);
nand U25921 (N_25921,N_25776,N_25659);
nand U25922 (N_25922,N_25619,N_25769);
and U25923 (N_25923,N_25533,N_25628);
or U25924 (N_25924,N_25766,N_25603);
or U25925 (N_25925,N_25797,N_25684);
nor U25926 (N_25926,N_25699,N_25584);
or U25927 (N_25927,N_25646,N_25575);
or U25928 (N_25928,N_25778,N_25574);
or U25929 (N_25929,N_25746,N_25674);
and U25930 (N_25930,N_25515,N_25588);
or U25931 (N_25931,N_25549,N_25626);
nand U25932 (N_25932,N_25675,N_25629);
xnor U25933 (N_25933,N_25605,N_25726);
and U25934 (N_25934,N_25673,N_25586);
nor U25935 (N_25935,N_25509,N_25784);
nor U25936 (N_25936,N_25696,N_25555);
xnor U25937 (N_25937,N_25782,N_25560);
and U25938 (N_25938,N_25663,N_25667);
xnor U25939 (N_25939,N_25571,N_25507);
or U25940 (N_25940,N_25765,N_25645);
nand U25941 (N_25941,N_25542,N_25638);
or U25942 (N_25942,N_25656,N_25644);
xor U25943 (N_25943,N_25787,N_25621);
and U25944 (N_25944,N_25749,N_25661);
or U25945 (N_25945,N_25545,N_25692);
or U25946 (N_25946,N_25713,N_25523);
nand U25947 (N_25947,N_25733,N_25652);
and U25948 (N_25948,N_25779,N_25728);
nand U25949 (N_25949,N_25744,N_25633);
nand U25950 (N_25950,N_25510,N_25557);
nor U25951 (N_25951,N_25724,N_25561);
xnor U25952 (N_25952,N_25659,N_25525);
or U25953 (N_25953,N_25583,N_25767);
nand U25954 (N_25954,N_25651,N_25537);
nand U25955 (N_25955,N_25638,N_25764);
xor U25956 (N_25956,N_25522,N_25516);
nor U25957 (N_25957,N_25609,N_25578);
nand U25958 (N_25958,N_25703,N_25741);
nor U25959 (N_25959,N_25549,N_25636);
xor U25960 (N_25960,N_25569,N_25637);
nand U25961 (N_25961,N_25578,N_25565);
nand U25962 (N_25962,N_25645,N_25604);
or U25963 (N_25963,N_25619,N_25664);
xnor U25964 (N_25964,N_25651,N_25563);
or U25965 (N_25965,N_25501,N_25709);
xor U25966 (N_25966,N_25516,N_25675);
xnor U25967 (N_25967,N_25525,N_25786);
and U25968 (N_25968,N_25610,N_25686);
xnor U25969 (N_25969,N_25508,N_25794);
and U25970 (N_25970,N_25753,N_25560);
and U25971 (N_25971,N_25771,N_25676);
or U25972 (N_25972,N_25783,N_25769);
xnor U25973 (N_25973,N_25610,N_25612);
and U25974 (N_25974,N_25556,N_25775);
nor U25975 (N_25975,N_25703,N_25663);
and U25976 (N_25976,N_25578,N_25690);
or U25977 (N_25977,N_25550,N_25707);
nand U25978 (N_25978,N_25521,N_25680);
and U25979 (N_25979,N_25755,N_25706);
nand U25980 (N_25980,N_25573,N_25749);
nand U25981 (N_25981,N_25780,N_25764);
nor U25982 (N_25982,N_25546,N_25736);
or U25983 (N_25983,N_25609,N_25541);
nand U25984 (N_25984,N_25558,N_25699);
nor U25985 (N_25985,N_25792,N_25738);
or U25986 (N_25986,N_25721,N_25522);
nand U25987 (N_25987,N_25548,N_25612);
xnor U25988 (N_25988,N_25675,N_25607);
xnor U25989 (N_25989,N_25554,N_25691);
and U25990 (N_25990,N_25676,N_25779);
nand U25991 (N_25991,N_25782,N_25696);
or U25992 (N_25992,N_25700,N_25762);
nor U25993 (N_25993,N_25506,N_25638);
nand U25994 (N_25994,N_25744,N_25602);
xnor U25995 (N_25995,N_25569,N_25633);
and U25996 (N_25996,N_25691,N_25597);
nand U25997 (N_25997,N_25555,N_25602);
and U25998 (N_25998,N_25719,N_25578);
and U25999 (N_25999,N_25799,N_25662);
and U26000 (N_26000,N_25776,N_25582);
xor U26001 (N_26001,N_25783,N_25518);
and U26002 (N_26002,N_25623,N_25582);
nor U26003 (N_26003,N_25633,N_25593);
xor U26004 (N_26004,N_25656,N_25749);
or U26005 (N_26005,N_25737,N_25663);
or U26006 (N_26006,N_25595,N_25502);
nand U26007 (N_26007,N_25514,N_25595);
xor U26008 (N_26008,N_25656,N_25584);
and U26009 (N_26009,N_25546,N_25547);
nand U26010 (N_26010,N_25684,N_25591);
nor U26011 (N_26011,N_25542,N_25541);
xor U26012 (N_26012,N_25656,N_25652);
or U26013 (N_26013,N_25759,N_25567);
nand U26014 (N_26014,N_25502,N_25590);
xnor U26015 (N_26015,N_25698,N_25506);
xor U26016 (N_26016,N_25541,N_25598);
and U26017 (N_26017,N_25785,N_25576);
or U26018 (N_26018,N_25768,N_25520);
nor U26019 (N_26019,N_25744,N_25778);
or U26020 (N_26020,N_25549,N_25693);
or U26021 (N_26021,N_25777,N_25672);
nand U26022 (N_26022,N_25736,N_25609);
and U26023 (N_26023,N_25556,N_25783);
nand U26024 (N_26024,N_25728,N_25510);
nand U26025 (N_26025,N_25630,N_25744);
nand U26026 (N_26026,N_25551,N_25641);
nand U26027 (N_26027,N_25731,N_25798);
nand U26028 (N_26028,N_25723,N_25517);
and U26029 (N_26029,N_25613,N_25531);
nor U26030 (N_26030,N_25514,N_25569);
nor U26031 (N_26031,N_25707,N_25528);
or U26032 (N_26032,N_25532,N_25685);
and U26033 (N_26033,N_25602,N_25573);
or U26034 (N_26034,N_25778,N_25725);
or U26035 (N_26035,N_25567,N_25609);
or U26036 (N_26036,N_25777,N_25771);
and U26037 (N_26037,N_25649,N_25783);
xnor U26038 (N_26038,N_25577,N_25657);
or U26039 (N_26039,N_25540,N_25572);
and U26040 (N_26040,N_25684,N_25600);
nor U26041 (N_26041,N_25653,N_25604);
or U26042 (N_26042,N_25659,N_25599);
xor U26043 (N_26043,N_25548,N_25528);
nand U26044 (N_26044,N_25682,N_25627);
and U26045 (N_26045,N_25603,N_25782);
and U26046 (N_26046,N_25665,N_25711);
nand U26047 (N_26047,N_25540,N_25768);
xnor U26048 (N_26048,N_25683,N_25645);
and U26049 (N_26049,N_25749,N_25727);
and U26050 (N_26050,N_25505,N_25588);
and U26051 (N_26051,N_25606,N_25689);
nor U26052 (N_26052,N_25585,N_25535);
xor U26053 (N_26053,N_25712,N_25569);
and U26054 (N_26054,N_25541,N_25515);
or U26055 (N_26055,N_25524,N_25769);
xnor U26056 (N_26056,N_25557,N_25699);
nand U26057 (N_26057,N_25656,N_25545);
and U26058 (N_26058,N_25548,N_25594);
nor U26059 (N_26059,N_25664,N_25626);
nand U26060 (N_26060,N_25529,N_25766);
nor U26061 (N_26061,N_25622,N_25545);
or U26062 (N_26062,N_25797,N_25598);
nand U26063 (N_26063,N_25653,N_25557);
xor U26064 (N_26064,N_25511,N_25516);
xor U26065 (N_26065,N_25659,N_25581);
nor U26066 (N_26066,N_25511,N_25656);
and U26067 (N_26067,N_25598,N_25568);
xor U26068 (N_26068,N_25616,N_25682);
and U26069 (N_26069,N_25637,N_25604);
or U26070 (N_26070,N_25735,N_25764);
xor U26071 (N_26071,N_25570,N_25717);
or U26072 (N_26072,N_25749,N_25630);
and U26073 (N_26073,N_25757,N_25542);
nor U26074 (N_26074,N_25620,N_25630);
nor U26075 (N_26075,N_25558,N_25565);
nor U26076 (N_26076,N_25636,N_25770);
xnor U26077 (N_26077,N_25570,N_25750);
and U26078 (N_26078,N_25657,N_25536);
or U26079 (N_26079,N_25506,N_25584);
nand U26080 (N_26080,N_25548,N_25551);
nor U26081 (N_26081,N_25530,N_25621);
or U26082 (N_26082,N_25755,N_25788);
and U26083 (N_26083,N_25755,N_25543);
or U26084 (N_26084,N_25751,N_25537);
and U26085 (N_26085,N_25624,N_25548);
and U26086 (N_26086,N_25526,N_25562);
nor U26087 (N_26087,N_25583,N_25742);
nor U26088 (N_26088,N_25646,N_25764);
xor U26089 (N_26089,N_25603,N_25507);
and U26090 (N_26090,N_25529,N_25787);
or U26091 (N_26091,N_25602,N_25655);
nand U26092 (N_26092,N_25778,N_25676);
nor U26093 (N_26093,N_25512,N_25757);
and U26094 (N_26094,N_25579,N_25642);
xnor U26095 (N_26095,N_25574,N_25745);
or U26096 (N_26096,N_25784,N_25716);
xnor U26097 (N_26097,N_25720,N_25783);
nor U26098 (N_26098,N_25747,N_25629);
and U26099 (N_26099,N_25601,N_25741);
or U26100 (N_26100,N_25835,N_25815);
and U26101 (N_26101,N_25869,N_26008);
and U26102 (N_26102,N_25924,N_25840);
nand U26103 (N_26103,N_26012,N_25824);
nand U26104 (N_26104,N_26034,N_25827);
or U26105 (N_26105,N_25871,N_25851);
nor U26106 (N_26106,N_25881,N_25816);
xnor U26107 (N_26107,N_25966,N_26060);
xor U26108 (N_26108,N_25984,N_25848);
or U26109 (N_26109,N_25938,N_26098);
or U26110 (N_26110,N_25844,N_26004);
nand U26111 (N_26111,N_25847,N_25822);
nor U26112 (N_26112,N_25953,N_25829);
nor U26113 (N_26113,N_25809,N_25939);
and U26114 (N_26114,N_25807,N_25957);
nand U26115 (N_26115,N_25880,N_26038);
and U26116 (N_26116,N_26081,N_25862);
or U26117 (N_26117,N_25927,N_25887);
nand U26118 (N_26118,N_25944,N_26031);
nand U26119 (N_26119,N_26094,N_25911);
xor U26120 (N_26120,N_25898,N_26088);
or U26121 (N_26121,N_25930,N_25821);
xnor U26122 (N_26122,N_26040,N_26086);
or U26123 (N_26123,N_26052,N_26057);
nand U26124 (N_26124,N_25969,N_26002);
nand U26125 (N_26125,N_25876,N_25996);
nor U26126 (N_26126,N_26019,N_26048);
nor U26127 (N_26127,N_25842,N_25895);
or U26128 (N_26128,N_26033,N_26027);
xnor U26129 (N_26129,N_25900,N_25846);
nor U26130 (N_26130,N_25997,N_25933);
or U26131 (N_26131,N_25998,N_26064);
xor U26132 (N_26132,N_25982,N_26080);
and U26133 (N_26133,N_26077,N_25956);
or U26134 (N_26134,N_25987,N_25920);
nor U26135 (N_26135,N_26028,N_26076);
nor U26136 (N_26136,N_25905,N_25978);
nand U26137 (N_26137,N_25926,N_25834);
nand U26138 (N_26138,N_26083,N_26021);
xor U26139 (N_26139,N_25906,N_25903);
and U26140 (N_26140,N_25885,N_25909);
xnor U26141 (N_26141,N_25837,N_25979);
nor U26142 (N_26142,N_25802,N_25872);
or U26143 (N_26143,N_25845,N_25942);
or U26144 (N_26144,N_25878,N_25897);
and U26145 (N_26145,N_25819,N_25950);
nand U26146 (N_26146,N_25864,N_25908);
nor U26147 (N_26147,N_25931,N_26085);
or U26148 (N_26148,N_25891,N_26062);
nor U26149 (N_26149,N_25970,N_25983);
nor U26150 (N_26150,N_25877,N_25971);
nand U26151 (N_26151,N_26072,N_25910);
or U26152 (N_26152,N_26056,N_25855);
and U26153 (N_26153,N_25896,N_25940);
xor U26154 (N_26154,N_26001,N_26084);
nand U26155 (N_26155,N_26090,N_25951);
xnor U26156 (N_26156,N_26070,N_25865);
nor U26157 (N_26157,N_25935,N_26026);
and U26158 (N_26158,N_25858,N_26075);
or U26159 (N_26159,N_25919,N_25873);
nand U26160 (N_26160,N_25811,N_25921);
xnor U26161 (N_26161,N_25828,N_25886);
nand U26162 (N_26162,N_25976,N_25959);
or U26163 (N_26163,N_26013,N_25913);
xor U26164 (N_26164,N_25960,N_26032);
nand U26165 (N_26165,N_25985,N_26067);
and U26166 (N_26166,N_25946,N_25836);
and U26167 (N_26167,N_25831,N_25907);
and U26168 (N_26168,N_25949,N_25810);
and U26169 (N_26169,N_26010,N_25849);
or U26170 (N_26170,N_26018,N_26051);
xnor U26171 (N_26171,N_25964,N_26071);
nand U26172 (N_26172,N_25967,N_26069);
and U26173 (N_26173,N_25994,N_26082);
nor U26174 (N_26174,N_26055,N_26050);
or U26175 (N_26175,N_26065,N_26089);
and U26176 (N_26176,N_25936,N_25916);
nor U26177 (N_26177,N_26000,N_26005);
xor U26178 (N_26178,N_25820,N_25965);
and U26179 (N_26179,N_25805,N_25806);
nor U26180 (N_26180,N_26099,N_26023);
xnor U26181 (N_26181,N_25801,N_25986);
xor U26182 (N_26182,N_25952,N_26029);
xor U26183 (N_26183,N_26047,N_26046);
and U26184 (N_26184,N_25914,N_25902);
or U26185 (N_26185,N_25947,N_26003);
xor U26186 (N_26186,N_26014,N_25892);
or U26187 (N_26187,N_25859,N_25808);
or U26188 (N_26188,N_25812,N_26015);
nor U26189 (N_26189,N_26037,N_25974);
nand U26190 (N_26190,N_25863,N_25856);
nor U26191 (N_26191,N_26030,N_25826);
and U26192 (N_26192,N_26016,N_25899);
or U26193 (N_26193,N_26097,N_25825);
xnor U26194 (N_26194,N_25814,N_25961);
xor U26195 (N_26195,N_26078,N_25923);
and U26196 (N_26196,N_25830,N_26068);
nand U26197 (N_26197,N_25857,N_26039);
xnor U26198 (N_26198,N_25963,N_26035);
xnor U26199 (N_26199,N_25893,N_25925);
or U26200 (N_26200,N_26041,N_25884);
xnor U26201 (N_26201,N_25817,N_25813);
or U26202 (N_26202,N_25922,N_26009);
or U26203 (N_26203,N_25852,N_26092);
xnor U26204 (N_26204,N_25894,N_26073);
xnor U26205 (N_26205,N_25843,N_25975);
or U26206 (N_26206,N_25928,N_26061);
or U26207 (N_26207,N_26053,N_25932);
and U26208 (N_26208,N_25839,N_26045);
and U26209 (N_26209,N_26042,N_25883);
nor U26210 (N_26210,N_25934,N_25954);
and U26211 (N_26211,N_25992,N_25866);
and U26212 (N_26212,N_25838,N_25941);
xnor U26213 (N_26213,N_25929,N_25832);
nand U26214 (N_26214,N_25988,N_25853);
nor U26215 (N_26215,N_26058,N_25875);
xor U26216 (N_26216,N_25945,N_26066);
nor U26217 (N_26217,N_25868,N_26043);
xnor U26218 (N_26218,N_25990,N_26036);
nor U26219 (N_26219,N_26006,N_25993);
nand U26220 (N_26220,N_25989,N_25841);
nor U26221 (N_26221,N_26022,N_25948);
nand U26222 (N_26222,N_25850,N_26087);
nand U26223 (N_26223,N_25912,N_26024);
and U26224 (N_26224,N_26059,N_25882);
or U26225 (N_26225,N_26017,N_25980);
or U26226 (N_26226,N_26093,N_25823);
or U26227 (N_26227,N_25999,N_25870);
xnor U26228 (N_26228,N_26063,N_25800);
and U26229 (N_26229,N_26096,N_25943);
nand U26230 (N_26230,N_25888,N_25904);
nor U26231 (N_26231,N_25995,N_25901);
nand U26232 (N_26232,N_25972,N_25854);
xor U26233 (N_26233,N_26011,N_26049);
nor U26234 (N_26234,N_26020,N_25867);
nand U26235 (N_26235,N_26091,N_26095);
nor U26236 (N_26236,N_25861,N_25889);
nand U26237 (N_26237,N_25977,N_26007);
nand U26238 (N_26238,N_26044,N_25818);
nand U26239 (N_26239,N_25917,N_25937);
nand U26240 (N_26240,N_25958,N_25833);
and U26241 (N_26241,N_25879,N_25803);
nor U26242 (N_26242,N_26079,N_25981);
or U26243 (N_26243,N_25955,N_26025);
xnor U26244 (N_26244,N_26054,N_25874);
and U26245 (N_26245,N_25915,N_25962);
xor U26246 (N_26246,N_25860,N_25973);
nand U26247 (N_26247,N_25968,N_25918);
nor U26248 (N_26248,N_25991,N_25890);
nand U26249 (N_26249,N_25804,N_26074);
xor U26250 (N_26250,N_26004,N_25924);
and U26251 (N_26251,N_25886,N_25897);
nor U26252 (N_26252,N_26016,N_25999);
and U26253 (N_26253,N_25996,N_25973);
or U26254 (N_26254,N_26057,N_25864);
or U26255 (N_26255,N_26020,N_26040);
xnor U26256 (N_26256,N_25836,N_25933);
or U26257 (N_26257,N_25802,N_25815);
or U26258 (N_26258,N_26030,N_25809);
nand U26259 (N_26259,N_26029,N_25821);
xor U26260 (N_26260,N_25906,N_25982);
xnor U26261 (N_26261,N_25913,N_25959);
nor U26262 (N_26262,N_25844,N_25882);
nor U26263 (N_26263,N_25828,N_26076);
xor U26264 (N_26264,N_25806,N_25927);
nor U26265 (N_26265,N_25853,N_25836);
or U26266 (N_26266,N_25885,N_25841);
or U26267 (N_26267,N_26025,N_25877);
xor U26268 (N_26268,N_25883,N_26008);
or U26269 (N_26269,N_26058,N_25855);
xor U26270 (N_26270,N_25955,N_25997);
and U26271 (N_26271,N_25858,N_26071);
or U26272 (N_26272,N_25894,N_25980);
and U26273 (N_26273,N_26043,N_26076);
nor U26274 (N_26274,N_25948,N_26053);
nand U26275 (N_26275,N_26090,N_25918);
xnor U26276 (N_26276,N_25862,N_25811);
nor U26277 (N_26277,N_26049,N_25831);
xor U26278 (N_26278,N_26021,N_25836);
or U26279 (N_26279,N_25876,N_25844);
xnor U26280 (N_26280,N_26015,N_26030);
nand U26281 (N_26281,N_25905,N_26089);
nand U26282 (N_26282,N_26033,N_25939);
and U26283 (N_26283,N_25990,N_26058);
or U26284 (N_26284,N_26091,N_26022);
and U26285 (N_26285,N_26095,N_25897);
xor U26286 (N_26286,N_25908,N_26018);
or U26287 (N_26287,N_26039,N_26089);
xor U26288 (N_26288,N_25864,N_26075);
nor U26289 (N_26289,N_25808,N_25847);
and U26290 (N_26290,N_26082,N_26072);
nor U26291 (N_26291,N_25841,N_26076);
nor U26292 (N_26292,N_25869,N_25892);
xnor U26293 (N_26293,N_25889,N_26084);
or U26294 (N_26294,N_26036,N_25910);
nand U26295 (N_26295,N_25977,N_25947);
and U26296 (N_26296,N_26057,N_25841);
or U26297 (N_26297,N_25837,N_26042);
or U26298 (N_26298,N_26074,N_26097);
and U26299 (N_26299,N_25945,N_25918);
and U26300 (N_26300,N_25926,N_25912);
nand U26301 (N_26301,N_25887,N_26009);
xnor U26302 (N_26302,N_25963,N_25962);
nand U26303 (N_26303,N_25809,N_25937);
or U26304 (N_26304,N_25991,N_26074);
and U26305 (N_26305,N_25955,N_25941);
xor U26306 (N_26306,N_26080,N_25803);
xnor U26307 (N_26307,N_25989,N_26023);
and U26308 (N_26308,N_25930,N_26016);
xnor U26309 (N_26309,N_26042,N_26037);
nor U26310 (N_26310,N_25845,N_25972);
nor U26311 (N_26311,N_25963,N_26057);
xnor U26312 (N_26312,N_25806,N_25954);
nand U26313 (N_26313,N_25865,N_25972);
nor U26314 (N_26314,N_25835,N_26001);
nand U26315 (N_26315,N_25921,N_25801);
or U26316 (N_26316,N_25871,N_26011);
nand U26317 (N_26317,N_25896,N_25831);
nor U26318 (N_26318,N_25922,N_26029);
or U26319 (N_26319,N_25940,N_25948);
nand U26320 (N_26320,N_25938,N_26079);
and U26321 (N_26321,N_25863,N_25918);
and U26322 (N_26322,N_26057,N_25964);
or U26323 (N_26323,N_25857,N_25811);
nor U26324 (N_26324,N_26058,N_25835);
nand U26325 (N_26325,N_26011,N_25958);
nor U26326 (N_26326,N_25903,N_25949);
nand U26327 (N_26327,N_25871,N_25867);
nor U26328 (N_26328,N_26039,N_26052);
nand U26329 (N_26329,N_25916,N_26001);
nor U26330 (N_26330,N_25958,N_26089);
or U26331 (N_26331,N_25994,N_25884);
and U26332 (N_26332,N_25951,N_25958);
xnor U26333 (N_26333,N_25924,N_25841);
or U26334 (N_26334,N_25996,N_25851);
xor U26335 (N_26335,N_25905,N_25981);
or U26336 (N_26336,N_25831,N_25854);
nor U26337 (N_26337,N_25878,N_25886);
xnor U26338 (N_26338,N_26077,N_26021);
or U26339 (N_26339,N_26002,N_25817);
xnor U26340 (N_26340,N_26011,N_26025);
xnor U26341 (N_26341,N_25983,N_25960);
xor U26342 (N_26342,N_26009,N_25952);
and U26343 (N_26343,N_25947,N_25955);
or U26344 (N_26344,N_25824,N_26008);
nor U26345 (N_26345,N_25842,N_25906);
nor U26346 (N_26346,N_26093,N_25857);
or U26347 (N_26347,N_25825,N_25829);
xor U26348 (N_26348,N_25876,N_26016);
and U26349 (N_26349,N_25927,N_25989);
or U26350 (N_26350,N_25912,N_25996);
and U26351 (N_26351,N_25893,N_25834);
nand U26352 (N_26352,N_26085,N_25823);
and U26353 (N_26353,N_26040,N_25990);
nand U26354 (N_26354,N_25825,N_26026);
xor U26355 (N_26355,N_25929,N_25834);
nand U26356 (N_26356,N_26046,N_26023);
xnor U26357 (N_26357,N_26014,N_25876);
xnor U26358 (N_26358,N_26032,N_25894);
nor U26359 (N_26359,N_25992,N_25817);
and U26360 (N_26360,N_26046,N_26034);
nand U26361 (N_26361,N_25840,N_26021);
xnor U26362 (N_26362,N_26033,N_25908);
nand U26363 (N_26363,N_25960,N_25889);
and U26364 (N_26364,N_25887,N_25955);
or U26365 (N_26365,N_26059,N_25867);
nor U26366 (N_26366,N_25881,N_25867);
or U26367 (N_26367,N_25873,N_25938);
xor U26368 (N_26368,N_26070,N_25916);
nor U26369 (N_26369,N_25878,N_25972);
nor U26370 (N_26370,N_26049,N_26030);
xor U26371 (N_26371,N_26012,N_26085);
xnor U26372 (N_26372,N_26029,N_26027);
and U26373 (N_26373,N_25973,N_26076);
xor U26374 (N_26374,N_25857,N_26016);
nand U26375 (N_26375,N_26038,N_26077);
xnor U26376 (N_26376,N_25828,N_25933);
or U26377 (N_26377,N_25839,N_26067);
nand U26378 (N_26378,N_25847,N_25929);
nor U26379 (N_26379,N_25935,N_25922);
xor U26380 (N_26380,N_25925,N_25892);
nor U26381 (N_26381,N_25809,N_25955);
nor U26382 (N_26382,N_25872,N_26043);
or U26383 (N_26383,N_25833,N_25908);
nor U26384 (N_26384,N_26085,N_25937);
nand U26385 (N_26385,N_25875,N_26079);
and U26386 (N_26386,N_25925,N_25970);
xor U26387 (N_26387,N_26032,N_25904);
nor U26388 (N_26388,N_26026,N_25867);
nor U26389 (N_26389,N_25998,N_25904);
or U26390 (N_26390,N_25977,N_25934);
nand U26391 (N_26391,N_25960,N_25964);
and U26392 (N_26392,N_25878,N_26051);
or U26393 (N_26393,N_26016,N_25806);
and U26394 (N_26394,N_25928,N_25896);
nor U26395 (N_26395,N_26086,N_26002);
nand U26396 (N_26396,N_25851,N_25825);
nor U26397 (N_26397,N_26044,N_25999);
and U26398 (N_26398,N_25918,N_26003);
and U26399 (N_26399,N_25829,N_25970);
nand U26400 (N_26400,N_26126,N_26255);
nor U26401 (N_26401,N_26142,N_26278);
xor U26402 (N_26402,N_26220,N_26135);
nand U26403 (N_26403,N_26284,N_26140);
xnor U26404 (N_26404,N_26338,N_26151);
and U26405 (N_26405,N_26389,N_26305);
or U26406 (N_26406,N_26256,N_26211);
nand U26407 (N_26407,N_26311,N_26243);
nand U26408 (N_26408,N_26295,N_26346);
nor U26409 (N_26409,N_26349,N_26174);
and U26410 (N_26410,N_26313,N_26316);
or U26411 (N_26411,N_26351,N_26139);
nor U26412 (N_26412,N_26328,N_26108);
xnor U26413 (N_26413,N_26226,N_26297);
nor U26414 (N_26414,N_26285,N_26159);
or U26415 (N_26415,N_26114,N_26301);
xor U26416 (N_26416,N_26280,N_26384);
and U26417 (N_26417,N_26368,N_26250);
nand U26418 (N_26418,N_26204,N_26394);
and U26419 (N_26419,N_26375,N_26292);
and U26420 (N_26420,N_26132,N_26124);
nand U26421 (N_26421,N_26348,N_26342);
and U26422 (N_26422,N_26277,N_26373);
and U26423 (N_26423,N_26329,N_26109);
nand U26424 (N_26424,N_26196,N_26184);
or U26425 (N_26425,N_26296,N_26319);
and U26426 (N_26426,N_26261,N_26247);
or U26427 (N_26427,N_26272,N_26362);
nand U26428 (N_26428,N_26121,N_26339);
nand U26429 (N_26429,N_26103,N_26217);
nor U26430 (N_26430,N_26302,N_26252);
and U26431 (N_26431,N_26376,N_26123);
and U26432 (N_26432,N_26190,N_26183);
or U26433 (N_26433,N_26345,N_26265);
xor U26434 (N_26434,N_26393,N_26361);
xnor U26435 (N_26435,N_26344,N_26286);
and U26436 (N_26436,N_26372,N_26137);
or U26437 (N_26437,N_26143,N_26234);
nand U26438 (N_26438,N_26113,N_26175);
or U26439 (N_26439,N_26193,N_26206);
nor U26440 (N_26440,N_26288,N_26150);
nor U26441 (N_26441,N_26125,N_26299);
xor U26442 (N_26442,N_26101,N_26227);
nor U26443 (N_26443,N_26340,N_26127);
or U26444 (N_26444,N_26321,N_26100);
xor U26445 (N_26445,N_26177,N_26279);
or U26446 (N_26446,N_26399,N_26254);
xor U26447 (N_26447,N_26205,N_26326);
nand U26448 (N_26448,N_26336,N_26290);
nor U26449 (N_26449,N_26325,N_26385);
nand U26450 (N_26450,N_26129,N_26117);
nand U26451 (N_26451,N_26332,N_26187);
and U26452 (N_26452,N_26160,N_26240);
nor U26453 (N_26453,N_26315,N_26377);
or U26454 (N_26454,N_26179,N_26207);
and U26455 (N_26455,N_26337,N_26176);
nand U26456 (N_26456,N_26264,N_26270);
and U26457 (N_26457,N_26309,N_26102);
nor U26458 (N_26458,N_26221,N_26392);
or U26459 (N_26459,N_26259,N_26357);
nand U26460 (N_26460,N_26320,N_26324);
or U26461 (N_26461,N_26364,N_26171);
xnor U26462 (N_26462,N_26396,N_26258);
and U26463 (N_26463,N_26387,N_26267);
and U26464 (N_26464,N_26307,N_26369);
or U26465 (N_26465,N_26134,N_26147);
nand U26466 (N_26466,N_26225,N_26191);
nand U26467 (N_26467,N_26273,N_26363);
nand U26468 (N_26468,N_26120,N_26180);
and U26469 (N_26469,N_26386,N_26145);
xor U26470 (N_26470,N_26215,N_26287);
xnor U26471 (N_26471,N_26353,N_26249);
or U26472 (N_26472,N_26110,N_26367);
and U26473 (N_26473,N_26195,N_26189);
and U26474 (N_26474,N_26112,N_26341);
nor U26475 (N_26475,N_26209,N_26300);
nor U26476 (N_26476,N_26322,N_26167);
nand U26477 (N_26477,N_26383,N_26197);
and U26478 (N_26478,N_26260,N_26149);
and U26479 (N_26479,N_26323,N_26378);
nand U26480 (N_26480,N_26294,N_26172);
nand U26481 (N_26481,N_26158,N_26161);
nor U26482 (N_26482,N_26391,N_26350);
nor U26483 (N_26483,N_26192,N_26269);
or U26484 (N_26484,N_26238,N_26228);
xnor U26485 (N_26485,N_26388,N_26366);
and U26486 (N_26486,N_26154,N_26202);
nand U26487 (N_26487,N_26282,N_26356);
nand U26488 (N_26488,N_26198,N_26119);
or U26489 (N_26489,N_26186,N_26374);
and U26490 (N_26490,N_26116,N_26136);
or U26491 (N_26491,N_26153,N_26253);
and U26492 (N_26492,N_26141,N_26148);
nor U26493 (N_26493,N_26262,N_26105);
or U26494 (N_26494,N_26283,N_26230);
and U26495 (N_26495,N_26201,N_26168);
nor U26496 (N_26496,N_26232,N_26306);
or U26497 (N_26497,N_26334,N_26274);
xor U26498 (N_26498,N_26156,N_26185);
nand U26499 (N_26499,N_26303,N_26214);
nor U26500 (N_26500,N_26222,N_26398);
or U26501 (N_26501,N_26165,N_26241);
and U26502 (N_26502,N_26359,N_26251);
and U26503 (N_26503,N_26194,N_26268);
and U26504 (N_26504,N_26289,N_26219);
nor U26505 (N_26505,N_26163,N_26131);
or U26506 (N_26506,N_26347,N_26188);
nand U26507 (N_26507,N_26276,N_26263);
nand U26508 (N_26508,N_26178,N_26318);
and U26509 (N_26509,N_26275,N_26233);
nor U26510 (N_26510,N_26208,N_26162);
nor U26511 (N_26511,N_26212,N_26365);
xor U26512 (N_26512,N_26118,N_26371);
nor U26513 (N_26513,N_26293,N_26166);
or U26514 (N_26514,N_26379,N_26106);
nor U26515 (N_26515,N_26310,N_26128);
nor U26516 (N_26516,N_26257,N_26330);
xor U26517 (N_26517,N_26281,N_26200);
or U26518 (N_26518,N_26327,N_26354);
xnor U26519 (N_26519,N_26314,N_26170);
or U26520 (N_26520,N_26331,N_26104);
nand U26521 (N_26521,N_26130,N_26360);
nand U26522 (N_26522,N_26164,N_26111);
xnor U26523 (N_26523,N_26358,N_26155);
nor U26524 (N_26524,N_26199,N_26216);
nor U26525 (N_26525,N_26244,N_26245);
and U26526 (N_26526,N_26203,N_26237);
nor U26527 (N_26527,N_26146,N_26239);
xor U26528 (N_26528,N_26298,N_26304);
xor U26529 (N_26529,N_26213,N_26144);
xor U26530 (N_26530,N_26218,N_26169);
or U26531 (N_26531,N_26355,N_26246);
nor U26532 (N_26532,N_26390,N_26181);
nor U26533 (N_26533,N_26382,N_26395);
nand U26534 (N_26534,N_26173,N_26107);
nor U26535 (N_26535,N_26266,N_26224);
or U26536 (N_26536,N_26291,N_26122);
nor U26537 (N_26537,N_26271,N_26182);
and U26538 (N_26538,N_26223,N_26236);
nand U26539 (N_26539,N_26333,N_26157);
xor U26540 (N_26540,N_26308,N_26397);
nand U26541 (N_26541,N_26138,N_26115);
nor U26542 (N_26542,N_26317,N_26235);
and U26543 (N_26543,N_26312,N_26210);
or U26544 (N_26544,N_26229,N_26343);
nor U26545 (N_26545,N_26152,N_26370);
or U26546 (N_26546,N_26335,N_26381);
nand U26547 (N_26547,N_26248,N_26133);
nor U26548 (N_26548,N_26380,N_26231);
and U26549 (N_26549,N_26352,N_26242);
nor U26550 (N_26550,N_26286,N_26204);
or U26551 (N_26551,N_26167,N_26213);
nor U26552 (N_26552,N_26318,N_26260);
nand U26553 (N_26553,N_26186,N_26339);
nor U26554 (N_26554,N_26148,N_26323);
xnor U26555 (N_26555,N_26391,N_26318);
or U26556 (N_26556,N_26339,N_26345);
nand U26557 (N_26557,N_26236,N_26389);
nor U26558 (N_26558,N_26306,N_26271);
or U26559 (N_26559,N_26353,N_26190);
nand U26560 (N_26560,N_26354,N_26166);
nand U26561 (N_26561,N_26125,N_26126);
xnor U26562 (N_26562,N_26166,N_26382);
or U26563 (N_26563,N_26191,N_26359);
xnor U26564 (N_26564,N_26280,N_26293);
nand U26565 (N_26565,N_26287,N_26197);
or U26566 (N_26566,N_26269,N_26165);
or U26567 (N_26567,N_26102,N_26229);
or U26568 (N_26568,N_26208,N_26327);
and U26569 (N_26569,N_26365,N_26105);
nor U26570 (N_26570,N_26286,N_26358);
or U26571 (N_26571,N_26261,N_26103);
nor U26572 (N_26572,N_26320,N_26381);
or U26573 (N_26573,N_26140,N_26389);
or U26574 (N_26574,N_26300,N_26199);
nor U26575 (N_26575,N_26258,N_26357);
nand U26576 (N_26576,N_26359,N_26243);
xor U26577 (N_26577,N_26205,N_26266);
xnor U26578 (N_26578,N_26165,N_26385);
and U26579 (N_26579,N_26141,N_26305);
xnor U26580 (N_26580,N_26366,N_26111);
xnor U26581 (N_26581,N_26258,N_26288);
or U26582 (N_26582,N_26286,N_26289);
and U26583 (N_26583,N_26173,N_26135);
or U26584 (N_26584,N_26160,N_26354);
or U26585 (N_26585,N_26280,N_26271);
xor U26586 (N_26586,N_26197,N_26129);
nor U26587 (N_26587,N_26243,N_26127);
nand U26588 (N_26588,N_26233,N_26286);
nand U26589 (N_26589,N_26248,N_26356);
or U26590 (N_26590,N_26155,N_26236);
nand U26591 (N_26591,N_26206,N_26224);
xnor U26592 (N_26592,N_26342,N_26170);
nor U26593 (N_26593,N_26116,N_26110);
and U26594 (N_26594,N_26231,N_26370);
nand U26595 (N_26595,N_26395,N_26208);
nor U26596 (N_26596,N_26191,N_26246);
nand U26597 (N_26597,N_26234,N_26300);
or U26598 (N_26598,N_26181,N_26344);
and U26599 (N_26599,N_26137,N_26349);
nand U26600 (N_26600,N_26210,N_26354);
or U26601 (N_26601,N_26306,N_26377);
and U26602 (N_26602,N_26146,N_26268);
nand U26603 (N_26603,N_26304,N_26296);
xor U26604 (N_26604,N_26260,N_26388);
nor U26605 (N_26605,N_26329,N_26310);
and U26606 (N_26606,N_26277,N_26300);
nor U26607 (N_26607,N_26218,N_26323);
nor U26608 (N_26608,N_26192,N_26239);
xnor U26609 (N_26609,N_26190,N_26375);
xor U26610 (N_26610,N_26300,N_26136);
and U26611 (N_26611,N_26207,N_26320);
nor U26612 (N_26612,N_26140,N_26186);
nand U26613 (N_26613,N_26131,N_26176);
and U26614 (N_26614,N_26392,N_26182);
xor U26615 (N_26615,N_26144,N_26127);
and U26616 (N_26616,N_26306,N_26300);
nand U26617 (N_26617,N_26167,N_26366);
and U26618 (N_26618,N_26205,N_26251);
nor U26619 (N_26619,N_26257,N_26379);
xnor U26620 (N_26620,N_26162,N_26201);
and U26621 (N_26621,N_26281,N_26313);
and U26622 (N_26622,N_26130,N_26195);
or U26623 (N_26623,N_26362,N_26151);
nand U26624 (N_26624,N_26320,N_26238);
nand U26625 (N_26625,N_26216,N_26101);
nand U26626 (N_26626,N_26313,N_26166);
nor U26627 (N_26627,N_26250,N_26147);
nand U26628 (N_26628,N_26266,N_26238);
nand U26629 (N_26629,N_26304,N_26223);
nor U26630 (N_26630,N_26261,N_26381);
nor U26631 (N_26631,N_26204,N_26165);
nor U26632 (N_26632,N_26295,N_26259);
and U26633 (N_26633,N_26273,N_26251);
nand U26634 (N_26634,N_26255,N_26382);
and U26635 (N_26635,N_26212,N_26349);
and U26636 (N_26636,N_26314,N_26280);
nand U26637 (N_26637,N_26226,N_26113);
nand U26638 (N_26638,N_26142,N_26202);
xor U26639 (N_26639,N_26229,N_26275);
xnor U26640 (N_26640,N_26193,N_26299);
xor U26641 (N_26641,N_26132,N_26399);
and U26642 (N_26642,N_26276,N_26164);
or U26643 (N_26643,N_26212,N_26354);
and U26644 (N_26644,N_26246,N_26372);
or U26645 (N_26645,N_26382,N_26385);
nand U26646 (N_26646,N_26358,N_26378);
nand U26647 (N_26647,N_26251,N_26225);
nor U26648 (N_26648,N_26261,N_26289);
nand U26649 (N_26649,N_26167,N_26223);
xnor U26650 (N_26650,N_26328,N_26153);
nand U26651 (N_26651,N_26180,N_26302);
xor U26652 (N_26652,N_26140,N_26272);
xnor U26653 (N_26653,N_26327,N_26123);
nand U26654 (N_26654,N_26144,N_26108);
nand U26655 (N_26655,N_26356,N_26201);
nand U26656 (N_26656,N_26196,N_26360);
and U26657 (N_26657,N_26305,N_26107);
nand U26658 (N_26658,N_26131,N_26166);
nor U26659 (N_26659,N_26384,N_26117);
or U26660 (N_26660,N_26100,N_26177);
nor U26661 (N_26661,N_26281,N_26248);
nor U26662 (N_26662,N_26238,N_26237);
or U26663 (N_26663,N_26100,N_26199);
nand U26664 (N_26664,N_26154,N_26292);
xnor U26665 (N_26665,N_26320,N_26372);
xnor U26666 (N_26666,N_26387,N_26342);
xor U26667 (N_26667,N_26147,N_26229);
nand U26668 (N_26668,N_26226,N_26329);
or U26669 (N_26669,N_26347,N_26223);
nand U26670 (N_26670,N_26246,N_26361);
or U26671 (N_26671,N_26193,N_26103);
nand U26672 (N_26672,N_26329,N_26368);
xor U26673 (N_26673,N_26351,N_26338);
xnor U26674 (N_26674,N_26128,N_26175);
nand U26675 (N_26675,N_26286,N_26279);
nor U26676 (N_26676,N_26316,N_26153);
and U26677 (N_26677,N_26386,N_26304);
nor U26678 (N_26678,N_26345,N_26190);
or U26679 (N_26679,N_26287,N_26113);
nor U26680 (N_26680,N_26300,N_26180);
or U26681 (N_26681,N_26377,N_26121);
nor U26682 (N_26682,N_26113,N_26262);
or U26683 (N_26683,N_26258,N_26143);
xor U26684 (N_26684,N_26101,N_26394);
xnor U26685 (N_26685,N_26317,N_26370);
and U26686 (N_26686,N_26239,N_26150);
nand U26687 (N_26687,N_26246,N_26259);
and U26688 (N_26688,N_26146,N_26240);
xnor U26689 (N_26689,N_26247,N_26349);
nor U26690 (N_26690,N_26140,N_26168);
nand U26691 (N_26691,N_26131,N_26147);
nor U26692 (N_26692,N_26393,N_26125);
and U26693 (N_26693,N_26393,N_26246);
or U26694 (N_26694,N_26302,N_26381);
nor U26695 (N_26695,N_26175,N_26255);
nand U26696 (N_26696,N_26111,N_26119);
nand U26697 (N_26697,N_26348,N_26238);
nand U26698 (N_26698,N_26201,N_26335);
and U26699 (N_26699,N_26241,N_26354);
nand U26700 (N_26700,N_26532,N_26547);
or U26701 (N_26701,N_26697,N_26402);
xor U26702 (N_26702,N_26593,N_26699);
xor U26703 (N_26703,N_26613,N_26534);
xor U26704 (N_26704,N_26670,N_26644);
nand U26705 (N_26705,N_26612,N_26598);
xnor U26706 (N_26706,N_26431,N_26498);
or U26707 (N_26707,N_26489,N_26673);
and U26708 (N_26708,N_26496,N_26614);
nor U26709 (N_26709,N_26497,N_26453);
and U26710 (N_26710,N_26577,N_26422);
or U26711 (N_26711,N_26678,N_26521);
and U26712 (N_26712,N_26480,N_26597);
nor U26713 (N_26713,N_26579,N_26538);
and U26714 (N_26714,N_26416,N_26400);
nor U26715 (N_26715,N_26450,N_26500);
or U26716 (N_26716,N_26475,N_26466);
nor U26717 (N_26717,N_26444,N_26609);
or U26718 (N_26718,N_26533,N_26415);
nand U26719 (N_26719,N_26594,N_26565);
xor U26720 (N_26720,N_26640,N_26638);
or U26721 (N_26721,N_26601,N_26432);
and U26722 (N_26722,N_26523,N_26490);
nand U26723 (N_26723,N_26524,N_26441);
or U26724 (N_26724,N_26559,N_26504);
nor U26725 (N_26725,N_26560,N_26628);
and U26726 (N_26726,N_26464,N_26585);
nor U26727 (N_26727,N_26446,N_26478);
xnor U26728 (N_26728,N_26688,N_26588);
xor U26729 (N_26729,N_26417,N_26563);
xnor U26730 (N_26730,N_26470,N_26404);
and U26731 (N_26731,N_26541,N_26409);
and U26732 (N_26732,N_26539,N_26529);
or U26733 (N_26733,N_26526,N_26435);
and U26734 (N_26734,N_26590,N_26550);
xnor U26735 (N_26735,N_26557,N_26677);
and U26736 (N_26736,N_26462,N_26687);
nor U26737 (N_26737,N_26583,N_26679);
nor U26738 (N_26738,N_26611,N_26681);
and U26739 (N_26739,N_26499,N_26494);
nand U26740 (N_26740,N_26459,N_26599);
nor U26741 (N_26741,N_26692,N_26483);
xor U26742 (N_26742,N_26661,N_26669);
or U26743 (N_26743,N_26646,N_26648);
nor U26744 (N_26744,N_26554,N_26645);
or U26745 (N_26745,N_26680,N_26515);
nand U26746 (N_26746,N_26615,N_26649);
xnor U26747 (N_26747,N_26513,N_26682);
and U26748 (N_26748,N_26501,N_26636);
and U26749 (N_26749,N_26561,N_26549);
or U26750 (N_26750,N_26442,N_26476);
nor U26751 (N_26751,N_26572,N_26683);
xnor U26752 (N_26752,N_26684,N_26698);
xnor U26753 (N_26753,N_26627,N_26552);
nand U26754 (N_26754,N_26662,N_26642);
and U26755 (N_26755,N_26425,N_26472);
and U26756 (N_26756,N_26455,N_26535);
nand U26757 (N_26757,N_26405,N_26528);
and U26758 (N_26758,N_26508,N_26433);
or U26759 (N_26759,N_26482,N_26663);
nor U26760 (N_26760,N_26608,N_26568);
and U26761 (N_26761,N_26617,N_26545);
xor U26762 (N_26762,N_26510,N_26690);
or U26763 (N_26763,N_26492,N_26456);
or U26764 (N_26764,N_26556,N_26693);
nand U26765 (N_26765,N_26507,N_26695);
xor U26766 (N_26766,N_26516,N_26509);
nor U26767 (N_26767,N_26546,N_26481);
nor U26768 (N_26768,N_26460,N_26675);
or U26769 (N_26769,N_26449,N_26436);
or U26770 (N_26770,N_26471,N_26473);
and U26771 (N_26771,N_26465,N_26576);
and U26772 (N_26772,N_26625,N_26440);
nand U26773 (N_26773,N_26511,N_26424);
and U26774 (N_26774,N_26503,N_26639);
xor U26775 (N_26775,N_26401,N_26454);
or U26776 (N_26776,N_26600,N_26641);
nand U26777 (N_26777,N_26445,N_26610);
xor U26778 (N_26778,N_26578,N_26626);
nand U26779 (N_26779,N_26548,N_26637);
and U26780 (N_26780,N_26429,N_26451);
nor U26781 (N_26781,N_26696,N_26621);
nor U26782 (N_26782,N_26514,N_26660);
or U26783 (N_26783,N_26418,N_26652);
or U26784 (N_26784,N_26485,N_26408);
nor U26785 (N_26785,N_26537,N_26543);
and U26786 (N_26786,N_26536,N_26658);
nor U26787 (N_26787,N_26420,N_26562);
and U26788 (N_26788,N_26574,N_26634);
and U26789 (N_26789,N_26674,N_26421);
xor U26790 (N_26790,N_26635,N_26589);
and U26791 (N_26791,N_26691,N_26479);
nor U26792 (N_26792,N_26624,N_26604);
and U26793 (N_26793,N_26664,N_26522);
xor U26794 (N_26794,N_26527,N_26619);
nand U26795 (N_26795,N_26474,N_26505);
xor U26796 (N_26796,N_26566,N_26468);
and U26797 (N_26797,N_26668,N_26457);
or U26798 (N_26798,N_26428,N_26427);
nor U26799 (N_26799,N_26506,N_26406);
or U26800 (N_26800,N_26430,N_26676);
nand U26801 (N_26801,N_26419,N_26410);
xor U26802 (N_26802,N_26672,N_26407);
nor U26803 (N_26803,N_26423,N_26567);
or U26804 (N_26804,N_26651,N_26531);
or U26805 (N_26805,N_26493,N_26606);
and U26806 (N_26806,N_26438,N_26623);
nand U26807 (N_26807,N_26502,N_26631);
or U26808 (N_26808,N_26551,N_26656);
nand U26809 (N_26809,N_26517,N_26587);
and U26810 (N_26810,N_26582,N_26553);
nand U26811 (N_26811,N_26581,N_26512);
and U26812 (N_26812,N_26666,N_26484);
and U26813 (N_26813,N_26605,N_26592);
nand U26814 (N_26814,N_26458,N_26643);
nand U26815 (N_26815,N_26620,N_26414);
nand U26816 (N_26816,N_26654,N_26467);
or U26817 (N_26817,N_26530,N_26671);
and U26818 (N_26818,N_26540,N_26452);
or U26819 (N_26819,N_26632,N_26412);
nor U26820 (N_26820,N_26437,N_26443);
and U26821 (N_26821,N_26591,N_26448);
nand U26822 (N_26822,N_26580,N_26403);
or U26823 (N_26823,N_26665,N_26525);
or U26824 (N_26824,N_26469,N_26685);
nand U26825 (N_26825,N_26686,N_26463);
nor U26826 (N_26826,N_26573,N_26629);
and U26827 (N_26827,N_26518,N_26519);
nor U26828 (N_26828,N_26564,N_26477);
nor U26829 (N_26829,N_26439,N_26595);
or U26830 (N_26830,N_26495,N_26647);
nor U26831 (N_26831,N_26650,N_26630);
and U26832 (N_26832,N_26544,N_26426);
nor U26833 (N_26833,N_26689,N_26694);
nor U26834 (N_26834,N_26622,N_26602);
nand U26835 (N_26835,N_26520,N_26486);
nand U26836 (N_26836,N_26659,N_26570);
and U26837 (N_26837,N_26411,N_26571);
xnor U26838 (N_26838,N_26586,N_26667);
nand U26839 (N_26839,N_26555,N_26413);
xnor U26840 (N_26840,N_26653,N_26607);
nand U26841 (N_26841,N_26584,N_26542);
and U26842 (N_26842,N_26491,N_26603);
xnor U26843 (N_26843,N_26633,N_26434);
and U26844 (N_26844,N_26447,N_26487);
or U26845 (N_26845,N_26488,N_26616);
xor U26846 (N_26846,N_26596,N_26569);
or U26847 (N_26847,N_26657,N_26618);
and U26848 (N_26848,N_26558,N_26655);
nor U26849 (N_26849,N_26461,N_26575);
xor U26850 (N_26850,N_26688,N_26492);
xnor U26851 (N_26851,N_26627,N_26657);
nor U26852 (N_26852,N_26634,N_26540);
and U26853 (N_26853,N_26504,N_26627);
or U26854 (N_26854,N_26544,N_26599);
xnor U26855 (N_26855,N_26579,N_26420);
or U26856 (N_26856,N_26506,N_26453);
xnor U26857 (N_26857,N_26504,N_26448);
or U26858 (N_26858,N_26541,N_26486);
nand U26859 (N_26859,N_26618,N_26407);
nor U26860 (N_26860,N_26417,N_26490);
and U26861 (N_26861,N_26635,N_26578);
nor U26862 (N_26862,N_26412,N_26633);
xor U26863 (N_26863,N_26573,N_26649);
nand U26864 (N_26864,N_26651,N_26452);
or U26865 (N_26865,N_26479,N_26672);
nand U26866 (N_26866,N_26637,N_26635);
and U26867 (N_26867,N_26406,N_26593);
or U26868 (N_26868,N_26606,N_26596);
or U26869 (N_26869,N_26579,N_26481);
nor U26870 (N_26870,N_26611,N_26657);
xnor U26871 (N_26871,N_26629,N_26460);
or U26872 (N_26872,N_26453,N_26564);
or U26873 (N_26873,N_26499,N_26430);
nor U26874 (N_26874,N_26495,N_26636);
xor U26875 (N_26875,N_26447,N_26556);
nand U26876 (N_26876,N_26463,N_26507);
nor U26877 (N_26877,N_26616,N_26562);
and U26878 (N_26878,N_26604,N_26447);
or U26879 (N_26879,N_26596,N_26568);
or U26880 (N_26880,N_26695,N_26651);
nand U26881 (N_26881,N_26481,N_26695);
nand U26882 (N_26882,N_26678,N_26605);
nand U26883 (N_26883,N_26403,N_26696);
nand U26884 (N_26884,N_26401,N_26480);
nor U26885 (N_26885,N_26529,N_26442);
nor U26886 (N_26886,N_26407,N_26521);
and U26887 (N_26887,N_26610,N_26681);
or U26888 (N_26888,N_26461,N_26680);
xor U26889 (N_26889,N_26521,N_26657);
and U26890 (N_26890,N_26686,N_26516);
nand U26891 (N_26891,N_26498,N_26609);
nor U26892 (N_26892,N_26650,N_26452);
and U26893 (N_26893,N_26437,N_26536);
nor U26894 (N_26894,N_26542,N_26536);
and U26895 (N_26895,N_26542,N_26533);
and U26896 (N_26896,N_26694,N_26555);
xnor U26897 (N_26897,N_26530,N_26683);
nand U26898 (N_26898,N_26448,N_26618);
or U26899 (N_26899,N_26495,N_26442);
xor U26900 (N_26900,N_26411,N_26591);
nand U26901 (N_26901,N_26561,N_26525);
xor U26902 (N_26902,N_26633,N_26547);
nor U26903 (N_26903,N_26599,N_26421);
nor U26904 (N_26904,N_26417,N_26649);
nor U26905 (N_26905,N_26527,N_26636);
and U26906 (N_26906,N_26579,N_26468);
nand U26907 (N_26907,N_26579,N_26585);
xnor U26908 (N_26908,N_26572,N_26515);
or U26909 (N_26909,N_26450,N_26628);
or U26910 (N_26910,N_26493,N_26687);
nand U26911 (N_26911,N_26469,N_26425);
xor U26912 (N_26912,N_26610,N_26446);
nand U26913 (N_26913,N_26694,N_26514);
xnor U26914 (N_26914,N_26542,N_26435);
nand U26915 (N_26915,N_26563,N_26441);
nor U26916 (N_26916,N_26526,N_26410);
nand U26917 (N_26917,N_26560,N_26698);
nand U26918 (N_26918,N_26567,N_26534);
nand U26919 (N_26919,N_26410,N_26430);
xnor U26920 (N_26920,N_26537,N_26691);
or U26921 (N_26921,N_26607,N_26412);
and U26922 (N_26922,N_26546,N_26626);
or U26923 (N_26923,N_26653,N_26455);
or U26924 (N_26924,N_26617,N_26558);
nor U26925 (N_26925,N_26425,N_26426);
and U26926 (N_26926,N_26629,N_26451);
nor U26927 (N_26927,N_26618,N_26569);
nand U26928 (N_26928,N_26659,N_26483);
xor U26929 (N_26929,N_26659,N_26482);
xnor U26930 (N_26930,N_26408,N_26477);
nand U26931 (N_26931,N_26520,N_26415);
nor U26932 (N_26932,N_26490,N_26545);
xnor U26933 (N_26933,N_26492,N_26589);
nor U26934 (N_26934,N_26542,N_26530);
nand U26935 (N_26935,N_26585,N_26593);
or U26936 (N_26936,N_26666,N_26466);
xnor U26937 (N_26937,N_26628,N_26640);
xor U26938 (N_26938,N_26619,N_26523);
or U26939 (N_26939,N_26446,N_26667);
nand U26940 (N_26940,N_26603,N_26516);
nand U26941 (N_26941,N_26586,N_26576);
xnor U26942 (N_26942,N_26426,N_26442);
and U26943 (N_26943,N_26496,N_26445);
nand U26944 (N_26944,N_26482,N_26475);
nand U26945 (N_26945,N_26630,N_26616);
xor U26946 (N_26946,N_26447,N_26498);
or U26947 (N_26947,N_26489,N_26563);
nand U26948 (N_26948,N_26405,N_26494);
xnor U26949 (N_26949,N_26530,N_26537);
xnor U26950 (N_26950,N_26504,N_26694);
or U26951 (N_26951,N_26560,N_26490);
nand U26952 (N_26952,N_26690,N_26541);
nand U26953 (N_26953,N_26497,N_26403);
nor U26954 (N_26954,N_26671,N_26470);
nor U26955 (N_26955,N_26688,N_26490);
nand U26956 (N_26956,N_26607,N_26624);
xnor U26957 (N_26957,N_26479,N_26422);
xor U26958 (N_26958,N_26475,N_26556);
and U26959 (N_26959,N_26417,N_26529);
or U26960 (N_26960,N_26596,N_26501);
and U26961 (N_26961,N_26552,N_26599);
and U26962 (N_26962,N_26506,N_26584);
nor U26963 (N_26963,N_26636,N_26534);
nor U26964 (N_26964,N_26421,N_26571);
and U26965 (N_26965,N_26616,N_26486);
or U26966 (N_26966,N_26477,N_26461);
xor U26967 (N_26967,N_26539,N_26486);
xnor U26968 (N_26968,N_26562,N_26681);
xor U26969 (N_26969,N_26446,N_26659);
or U26970 (N_26970,N_26631,N_26580);
or U26971 (N_26971,N_26559,N_26508);
nand U26972 (N_26972,N_26411,N_26534);
and U26973 (N_26973,N_26681,N_26627);
nand U26974 (N_26974,N_26408,N_26657);
nor U26975 (N_26975,N_26565,N_26572);
nand U26976 (N_26976,N_26667,N_26550);
and U26977 (N_26977,N_26426,N_26637);
and U26978 (N_26978,N_26519,N_26543);
and U26979 (N_26979,N_26670,N_26590);
and U26980 (N_26980,N_26563,N_26535);
nand U26981 (N_26981,N_26571,N_26577);
and U26982 (N_26982,N_26658,N_26469);
nor U26983 (N_26983,N_26503,N_26466);
xnor U26984 (N_26984,N_26643,N_26487);
xor U26985 (N_26985,N_26524,N_26508);
or U26986 (N_26986,N_26522,N_26668);
nand U26987 (N_26987,N_26468,N_26439);
or U26988 (N_26988,N_26411,N_26440);
nor U26989 (N_26989,N_26587,N_26443);
nand U26990 (N_26990,N_26454,N_26416);
nand U26991 (N_26991,N_26685,N_26463);
xnor U26992 (N_26992,N_26407,N_26663);
nand U26993 (N_26993,N_26683,N_26632);
xnor U26994 (N_26994,N_26617,N_26556);
nor U26995 (N_26995,N_26503,N_26655);
or U26996 (N_26996,N_26421,N_26478);
or U26997 (N_26997,N_26656,N_26576);
or U26998 (N_26998,N_26410,N_26643);
xnor U26999 (N_26999,N_26429,N_26457);
nand U27000 (N_27000,N_26870,N_26966);
or U27001 (N_27001,N_26951,N_26715);
xor U27002 (N_27002,N_26842,N_26857);
nor U27003 (N_27003,N_26777,N_26821);
xnor U27004 (N_27004,N_26827,N_26930);
nor U27005 (N_27005,N_26820,N_26947);
and U27006 (N_27006,N_26853,N_26994);
or U27007 (N_27007,N_26750,N_26765);
or U27008 (N_27008,N_26868,N_26791);
nor U27009 (N_27009,N_26729,N_26969);
and U27010 (N_27010,N_26742,N_26976);
and U27011 (N_27011,N_26958,N_26898);
nor U27012 (N_27012,N_26788,N_26849);
xnor U27013 (N_27013,N_26984,N_26758);
nor U27014 (N_27014,N_26880,N_26978);
xnor U27015 (N_27015,N_26738,N_26812);
nor U27016 (N_27016,N_26957,N_26869);
nor U27017 (N_27017,N_26745,N_26997);
xor U27018 (N_27018,N_26771,N_26746);
xnor U27019 (N_27019,N_26814,N_26914);
or U27020 (N_27020,N_26961,N_26818);
xnor U27021 (N_27021,N_26916,N_26922);
or U27022 (N_27022,N_26942,N_26845);
or U27023 (N_27023,N_26907,N_26886);
nor U27024 (N_27024,N_26924,N_26761);
nand U27025 (N_27025,N_26800,N_26768);
nor U27026 (N_27026,N_26926,N_26720);
or U27027 (N_27027,N_26894,N_26811);
nor U27028 (N_27028,N_26776,N_26982);
nand U27029 (N_27029,N_26830,N_26872);
or U27030 (N_27030,N_26974,N_26784);
or U27031 (N_27031,N_26769,N_26836);
nand U27032 (N_27032,N_26902,N_26753);
nand U27033 (N_27033,N_26747,N_26712);
and U27034 (N_27034,N_26744,N_26834);
nand U27035 (N_27035,N_26877,N_26939);
nor U27036 (N_27036,N_26840,N_26838);
nand U27037 (N_27037,N_26839,N_26882);
or U27038 (N_27038,N_26911,N_26903);
and U27039 (N_27039,N_26835,N_26971);
or U27040 (N_27040,N_26987,N_26963);
xor U27041 (N_27041,N_26799,N_26796);
and U27042 (N_27042,N_26931,N_26708);
and U27043 (N_27043,N_26825,N_26783);
and U27044 (N_27044,N_26754,N_26908);
or U27045 (N_27045,N_26829,N_26970);
nand U27046 (N_27046,N_26779,N_26732);
and U27047 (N_27047,N_26837,N_26725);
nand U27048 (N_27048,N_26983,N_26988);
nor U27049 (N_27049,N_26833,N_26846);
nor U27050 (N_27050,N_26919,N_26756);
or U27051 (N_27051,N_26792,N_26852);
or U27052 (N_27052,N_26858,N_26824);
xnor U27053 (N_27053,N_26721,N_26941);
and U27054 (N_27054,N_26714,N_26813);
nand U27055 (N_27055,N_26881,N_26751);
xor U27056 (N_27056,N_26906,N_26933);
nand U27057 (N_27057,N_26900,N_26887);
xnor U27058 (N_27058,N_26936,N_26918);
and U27059 (N_27059,N_26782,N_26804);
and U27060 (N_27060,N_26706,N_26968);
nand U27061 (N_27061,N_26795,N_26920);
or U27062 (N_27062,N_26944,N_26895);
or U27063 (N_27063,N_26859,N_26901);
nand U27064 (N_27064,N_26705,N_26943);
nor U27065 (N_27065,N_26889,N_26938);
or U27066 (N_27066,N_26972,N_26703);
xor U27067 (N_27067,N_26711,N_26736);
or U27068 (N_27068,N_26992,N_26925);
or U27069 (N_27069,N_26945,N_26728);
nor U27070 (N_27070,N_26735,N_26989);
and U27071 (N_27071,N_26863,N_26798);
or U27072 (N_27072,N_26794,N_26921);
nor U27073 (N_27073,N_26910,N_26946);
and U27074 (N_27074,N_26831,N_26850);
xor U27075 (N_27075,N_26704,N_26733);
nor U27076 (N_27076,N_26977,N_26797);
or U27077 (N_27077,N_26937,N_26866);
and U27078 (N_27078,N_26897,N_26965);
and U27079 (N_27079,N_26803,N_26718);
nand U27080 (N_27080,N_26932,N_26973);
and U27081 (N_27081,N_26959,N_26826);
or U27082 (N_27082,N_26766,N_26995);
nor U27083 (N_27083,N_26905,N_26855);
or U27084 (N_27084,N_26752,N_26874);
nor U27085 (N_27085,N_26748,N_26785);
and U27086 (N_27086,N_26710,N_26847);
xnor U27087 (N_27087,N_26964,N_26888);
nand U27088 (N_27088,N_26891,N_26917);
or U27089 (N_27089,N_26913,N_26892);
and U27090 (N_27090,N_26861,N_26885);
and U27091 (N_27091,N_26760,N_26949);
nand U27092 (N_27092,N_26713,N_26884);
nor U27093 (N_27093,N_26876,N_26828);
nand U27094 (N_27094,N_26990,N_26979);
and U27095 (N_27095,N_26723,N_26808);
and U27096 (N_27096,N_26967,N_26865);
nand U27097 (N_27097,N_26896,N_26879);
xnor U27098 (N_27098,N_26817,N_26764);
or U27099 (N_27099,N_26991,N_26778);
or U27100 (N_27100,N_26755,N_26786);
nand U27101 (N_27101,N_26832,N_26940);
nor U27102 (N_27102,N_26890,N_26719);
xnor U27103 (N_27103,N_26962,N_26700);
and U27104 (N_27104,N_26860,N_26772);
or U27105 (N_27105,N_26999,N_26707);
xor U27106 (N_27106,N_26841,N_26993);
and U27107 (N_27107,N_26743,N_26802);
or U27108 (N_27108,N_26793,N_26727);
and U27109 (N_27109,N_26955,N_26734);
nand U27110 (N_27110,N_26717,N_26954);
nor U27111 (N_27111,N_26809,N_26960);
nor U27112 (N_27112,N_26883,N_26899);
or U27113 (N_27113,N_26815,N_26722);
xor U27114 (N_27114,N_26790,N_26843);
nand U27115 (N_27115,N_26774,N_26909);
nor U27116 (N_27116,N_26737,N_26929);
and U27117 (N_27117,N_26740,N_26948);
and U27118 (N_27118,N_26998,N_26819);
or U27119 (N_27119,N_26767,N_26867);
nor U27120 (N_27120,N_26851,N_26807);
nand U27121 (N_27121,N_26823,N_26844);
and U27122 (N_27122,N_26928,N_26981);
nand U27123 (N_27123,N_26780,N_26757);
nand U27124 (N_27124,N_26781,N_26856);
xor U27125 (N_27125,N_26953,N_26862);
and U27126 (N_27126,N_26775,N_26923);
and U27127 (N_27127,N_26854,N_26730);
nor U27128 (N_27128,N_26950,N_26875);
nand U27129 (N_27129,N_26816,N_26952);
nand U27130 (N_27130,N_26986,N_26935);
and U27131 (N_27131,N_26996,N_26805);
or U27132 (N_27132,N_26726,N_26980);
and U27133 (N_27133,N_26912,N_26975);
or U27134 (N_27134,N_26759,N_26770);
and U27135 (N_27135,N_26871,N_26864);
xor U27136 (N_27136,N_26701,N_26763);
xor U27137 (N_27137,N_26731,N_26724);
xor U27138 (N_27138,N_26773,N_26739);
nor U27139 (N_27139,N_26801,N_26985);
xnor U27140 (N_27140,N_26927,N_26787);
xnor U27141 (N_27141,N_26709,N_26822);
nor U27142 (N_27142,N_26702,N_26956);
xnor U27143 (N_27143,N_26915,N_26749);
or U27144 (N_27144,N_26810,N_26878);
and U27145 (N_27145,N_26716,N_26873);
xor U27146 (N_27146,N_26893,N_26741);
or U27147 (N_27147,N_26806,N_26789);
and U27148 (N_27148,N_26934,N_26762);
or U27149 (N_27149,N_26904,N_26848);
nor U27150 (N_27150,N_26763,N_26893);
nor U27151 (N_27151,N_26997,N_26880);
nand U27152 (N_27152,N_26954,N_26741);
xor U27153 (N_27153,N_26772,N_26839);
xnor U27154 (N_27154,N_26778,N_26951);
or U27155 (N_27155,N_26976,N_26963);
or U27156 (N_27156,N_26754,N_26964);
nand U27157 (N_27157,N_26853,N_26740);
xnor U27158 (N_27158,N_26889,N_26830);
nor U27159 (N_27159,N_26712,N_26714);
xnor U27160 (N_27160,N_26832,N_26992);
xnor U27161 (N_27161,N_26757,N_26739);
nor U27162 (N_27162,N_26771,N_26736);
or U27163 (N_27163,N_26750,N_26757);
nand U27164 (N_27164,N_26960,N_26885);
nor U27165 (N_27165,N_26938,N_26750);
and U27166 (N_27166,N_26848,N_26912);
or U27167 (N_27167,N_26991,N_26899);
or U27168 (N_27168,N_26807,N_26943);
nand U27169 (N_27169,N_26912,N_26718);
or U27170 (N_27170,N_26999,N_26717);
and U27171 (N_27171,N_26832,N_26994);
or U27172 (N_27172,N_26947,N_26831);
and U27173 (N_27173,N_26769,N_26731);
or U27174 (N_27174,N_26851,N_26981);
nor U27175 (N_27175,N_26715,N_26861);
or U27176 (N_27176,N_26728,N_26705);
nor U27177 (N_27177,N_26733,N_26868);
nand U27178 (N_27178,N_26850,N_26764);
xnor U27179 (N_27179,N_26898,N_26789);
xnor U27180 (N_27180,N_26706,N_26938);
and U27181 (N_27181,N_26943,N_26879);
or U27182 (N_27182,N_26809,N_26828);
nor U27183 (N_27183,N_26883,N_26927);
nand U27184 (N_27184,N_26728,N_26939);
nor U27185 (N_27185,N_26759,N_26900);
nand U27186 (N_27186,N_26912,N_26937);
or U27187 (N_27187,N_26980,N_26748);
and U27188 (N_27188,N_26952,N_26753);
xnor U27189 (N_27189,N_26889,N_26962);
or U27190 (N_27190,N_26712,N_26962);
nand U27191 (N_27191,N_26996,N_26764);
nor U27192 (N_27192,N_26988,N_26919);
nand U27193 (N_27193,N_26787,N_26929);
and U27194 (N_27194,N_26983,N_26852);
nor U27195 (N_27195,N_26856,N_26786);
or U27196 (N_27196,N_26846,N_26900);
or U27197 (N_27197,N_26963,N_26994);
nand U27198 (N_27198,N_26977,N_26724);
nor U27199 (N_27199,N_26855,N_26877);
nor U27200 (N_27200,N_26876,N_26989);
nand U27201 (N_27201,N_26755,N_26898);
or U27202 (N_27202,N_26850,N_26860);
and U27203 (N_27203,N_26991,N_26958);
nor U27204 (N_27204,N_26809,N_26791);
nand U27205 (N_27205,N_26728,N_26881);
or U27206 (N_27206,N_26865,N_26902);
xnor U27207 (N_27207,N_26885,N_26835);
and U27208 (N_27208,N_26991,N_26992);
nor U27209 (N_27209,N_26766,N_26789);
nand U27210 (N_27210,N_26823,N_26950);
and U27211 (N_27211,N_26830,N_26802);
and U27212 (N_27212,N_26817,N_26814);
nor U27213 (N_27213,N_26791,N_26843);
or U27214 (N_27214,N_26703,N_26899);
nor U27215 (N_27215,N_26799,N_26752);
nand U27216 (N_27216,N_26920,N_26759);
xor U27217 (N_27217,N_26896,N_26831);
xor U27218 (N_27218,N_26891,N_26960);
and U27219 (N_27219,N_26914,N_26996);
nand U27220 (N_27220,N_26992,N_26942);
and U27221 (N_27221,N_26799,N_26902);
and U27222 (N_27222,N_26956,N_26775);
or U27223 (N_27223,N_26750,N_26955);
or U27224 (N_27224,N_26981,N_26950);
xor U27225 (N_27225,N_26938,N_26856);
xor U27226 (N_27226,N_26842,N_26973);
or U27227 (N_27227,N_26774,N_26816);
nor U27228 (N_27228,N_26843,N_26769);
and U27229 (N_27229,N_26723,N_26977);
or U27230 (N_27230,N_26758,N_26924);
xnor U27231 (N_27231,N_26854,N_26856);
and U27232 (N_27232,N_26835,N_26832);
nand U27233 (N_27233,N_26806,N_26858);
nand U27234 (N_27234,N_26706,N_26704);
nand U27235 (N_27235,N_26827,N_26990);
and U27236 (N_27236,N_26753,N_26846);
nor U27237 (N_27237,N_26812,N_26802);
and U27238 (N_27238,N_26856,N_26971);
and U27239 (N_27239,N_26949,N_26771);
xnor U27240 (N_27240,N_26719,N_26782);
nor U27241 (N_27241,N_26769,N_26904);
nand U27242 (N_27242,N_26945,N_26865);
nand U27243 (N_27243,N_26941,N_26980);
or U27244 (N_27244,N_26975,N_26771);
nor U27245 (N_27245,N_26755,N_26970);
xor U27246 (N_27246,N_26990,N_26973);
or U27247 (N_27247,N_26864,N_26855);
xor U27248 (N_27248,N_26816,N_26715);
or U27249 (N_27249,N_26961,N_26856);
or U27250 (N_27250,N_26816,N_26724);
and U27251 (N_27251,N_26838,N_26766);
xnor U27252 (N_27252,N_26756,N_26835);
xnor U27253 (N_27253,N_26905,N_26717);
xnor U27254 (N_27254,N_26980,N_26786);
nor U27255 (N_27255,N_26743,N_26725);
or U27256 (N_27256,N_26964,N_26755);
and U27257 (N_27257,N_26756,N_26799);
or U27258 (N_27258,N_26950,N_26756);
nor U27259 (N_27259,N_26868,N_26871);
xor U27260 (N_27260,N_26846,N_26997);
xnor U27261 (N_27261,N_26943,N_26740);
xnor U27262 (N_27262,N_26788,N_26889);
nor U27263 (N_27263,N_26937,N_26828);
nor U27264 (N_27264,N_26810,N_26779);
nand U27265 (N_27265,N_26985,N_26879);
and U27266 (N_27266,N_26997,N_26986);
xor U27267 (N_27267,N_26823,N_26834);
and U27268 (N_27268,N_26912,N_26706);
nor U27269 (N_27269,N_26810,N_26807);
xor U27270 (N_27270,N_26837,N_26920);
nor U27271 (N_27271,N_26743,N_26998);
nor U27272 (N_27272,N_26744,N_26932);
xor U27273 (N_27273,N_26800,N_26989);
or U27274 (N_27274,N_26886,N_26959);
nor U27275 (N_27275,N_26860,N_26799);
nor U27276 (N_27276,N_26901,N_26898);
nand U27277 (N_27277,N_26897,N_26794);
and U27278 (N_27278,N_26880,N_26838);
nor U27279 (N_27279,N_26998,N_26737);
or U27280 (N_27280,N_26958,N_26899);
xor U27281 (N_27281,N_26717,N_26956);
or U27282 (N_27282,N_26804,N_26943);
or U27283 (N_27283,N_26775,N_26788);
and U27284 (N_27284,N_26876,N_26887);
nand U27285 (N_27285,N_26783,N_26743);
nand U27286 (N_27286,N_26929,N_26766);
xor U27287 (N_27287,N_26992,N_26952);
and U27288 (N_27288,N_26907,N_26813);
nor U27289 (N_27289,N_26888,N_26744);
and U27290 (N_27290,N_26909,N_26980);
xor U27291 (N_27291,N_26922,N_26731);
xor U27292 (N_27292,N_26889,N_26821);
and U27293 (N_27293,N_26938,N_26902);
and U27294 (N_27294,N_26731,N_26970);
xor U27295 (N_27295,N_26945,N_26887);
or U27296 (N_27296,N_26815,N_26971);
nor U27297 (N_27297,N_26911,N_26951);
nor U27298 (N_27298,N_26825,N_26980);
nand U27299 (N_27299,N_26794,N_26899);
xor U27300 (N_27300,N_27190,N_27281);
and U27301 (N_27301,N_27150,N_27160);
or U27302 (N_27302,N_27277,N_27103);
xor U27303 (N_27303,N_27020,N_27108);
and U27304 (N_27304,N_27253,N_27233);
nand U27305 (N_27305,N_27204,N_27180);
nor U27306 (N_27306,N_27000,N_27032);
and U27307 (N_27307,N_27275,N_27206);
nor U27308 (N_27308,N_27130,N_27066);
xnor U27309 (N_27309,N_27070,N_27057);
or U27310 (N_27310,N_27207,N_27231);
nand U27311 (N_27311,N_27126,N_27133);
nor U27312 (N_27312,N_27124,N_27143);
xor U27313 (N_27313,N_27257,N_27221);
nor U27314 (N_27314,N_27227,N_27240);
and U27315 (N_27315,N_27028,N_27251);
xnor U27316 (N_27316,N_27012,N_27282);
and U27317 (N_27317,N_27099,N_27080);
nor U27318 (N_27318,N_27236,N_27263);
nor U27319 (N_27319,N_27139,N_27129);
and U27320 (N_27320,N_27161,N_27094);
and U27321 (N_27321,N_27025,N_27211);
nand U27322 (N_27322,N_27093,N_27235);
xor U27323 (N_27323,N_27015,N_27260);
nand U27324 (N_27324,N_27258,N_27232);
and U27325 (N_27325,N_27069,N_27121);
nor U27326 (N_27326,N_27076,N_27247);
or U27327 (N_27327,N_27030,N_27174);
and U27328 (N_27328,N_27285,N_27119);
nand U27329 (N_27329,N_27220,N_27291);
and U27330 (N_27330,N_27064,N_27050);
nor U27331 (N_27331,N_27244,N_27265);
and U27332 (N_27332,N_27185,N_27138);
and U27333 (N_27333,N_27026,N_27092);
xor U27334 (N_27334,N_27001,N_27034);
nor U27335 (N_27335,N_27250,N_27131);
nor U27336 (N_27336,N_27033,N_27114);
or U27337 (N_27337,N_27072,N_27089);
xnor U27338 (N_27338,N_27088,N_27061);
xor U27339 (N_27339,N_27023,N_27037);
xnor U27340 (N_27340,N_27195,N_27154);
nor U27341 (N_27341,N_27128,N_27019);
and U27342 (N_27342,N_27002,N_27043);
xnor U27343 (N_27343,N_27065,N_27157);
nor U27344 (N_27344,N_27172,N_27073);
or U27345 (N_27345,N_27115,N_27009);
nand U27346 (N_27346,N_27175,N_27283);
xor U27347 (N_27347,N_27156,N_27010);
xnor U27348 (N_27348,N_27209,N_27219);
or U27349 (N_27349,N_27041,N_27212);
nand U27350 (N_27350,N_27270,N_27062);
nand U27351 (N_27351,N_27224,N_27152);
nand U27352 (N_27352,N_27040,N_27217);
xnor U27353 (N_27353,N_27113,N_27081);
and U27354 (N_27354,N_27038,N_27228);
nor U27355 (N_27355,N_27117,N_27239);
nand U27356 (N_27356,N_27045,N_27176);
nor U27357 (N_27357,N_27059,N_27036);
or U27358 (N_27358,N_27031,N_27159);
nand U27359 (N_27359,N_27162,N_27248);
nor U27360 (N_27360,N_27004,N_27086);
and U27361 (N_27361,N_27272,N_27183);
or U27362 (N_27362,N_27170,N_27268);
and U27363 (N_27363,N_27091,N_27196);
nor U27364 (N_27364,N_27218,N_27164);
and U27365 (N_27365,N_27027,N_27039);
nand U27366 (N_27366,N_27024,N_27169);
nand U27367 (N_27367,N_27163,N_27046);
and U27368 (N_27368,N_27137,N_27189);
and U27369 (N_27369,N_27238,N_27146);
nor U27370 (N_27370,N_27298,N_27029);
xnor U27371 (N_27371,N_27230,N_27111);
and U27372 (N_27372,N_27003,N_27063);
or U27373 (N_27373,N_27213,N_27256);
or U27374 (N_27374,N_27241,N_27179);
nand U27375 (N_27375,N_27123,N_27048);
nor U27376 (N_27376,N_27203,N_27118);
xor U27377 (N_27377,N_27278,N_27178);
nor U27378 (N_27378,N_27021,N_27249);
nand U27379 (N_27379,N_27171,N_27007);
nand U27380 (N_27380,N_27110,N_27293);
and U27381 (N_27381,N_27144,N_27142);
nand U27382 (N_27382,N_27223,N_27214);
and U27383 (N_27383,N_27229,N_27120);
nand U27384 (N_27384,N_27254,N_27056);
nor U27385 (N_27385,N_27096,N_27122);
xnor U27386 (N_27386,N_27284,N_27005);
xnor U27387 (N_27387,N_27077,N_27255);
nor U27388 (N_27388,N_27084,N_27177);
nand U27389 (N_27389,N_27273,N_27226);
nor U27390 (N_27390,N_27097,N_27058);
nor U27391 (N_27391,N_27068,N_27205);
and U27392 (N_27392,N_27181,N_27299);
xor U27393 (N_27393,N_27289,N_27071);
and U27394 (N_27394,N_27112,N_27262);
and U27395 (N_27395,N_27044,N_27132);
and U27396 (N_27396,N_27201,N_27271);
or U27397 (N_27397,N_27148,N_27053);
and U27398 (N_27398,N_27049,N_27018);
and U27399 (N_27399,N_27125,N_27098);
nand U27400 (N_27400,N_27100,N_27295);
xor U27401 (N_27401,N_27136,N_27075);
nor U27402 (N_27402,N_27290,N_27184);
or U27403 (N_27403,N_27165,N_27101);
nor U27404 (N_27404,N_27017,N_27167);
nor U27405 (N_27405,N_27149,N_27198);
nor U27406 (N_27406,N_27182,N_27286);
nand U27407 (N_27407,N_27067,N_27083);
xnor U27408 (N_27408,N_27274,N_27060);
xnor U27409 (N_27409,N_27259,N_27035);
nand U27410 (N_27410,N_27187,N_27013);
and U27411 (N_27411,N_27102,N_27085);
xor U27412 (N_27412,N_27192,N_27051);
nand U27413 (N_27413,N_27266,N_27145);
xnor U27414 (N_27414,N_27074,N_27042);
and U27415 (N_27415,N_27287,N_27104);
xor U27416 (N_27416,N_27246,N_27116);
and U27417 (N_27417,N_27261,N_27082);
or U27418 (N_27418,N_27155,N_27016);
nand U27419 (N_27419,N_27078,N_27158);
nand U27420 (N_27420,N_27216,N_27210);
xor U27421 (N_27421,N_27140,N_27193);
or U27422 (N_27422,N_27200,N_27276);
nor U27423 (N_27423,N_27197,N_27186);
nand U27424 (N_27424,N_27269,N_27279);
or U27425 (N_27425,N_27014,N_27141);
and U27426 (N_27426,N_27134,N_27052);
or U27427 (N_27427,N_27264,N_27234);
nor U27428 (N_27428,N_27127,N_27090);
xnor U27429 (N_27429,N_27106,N_27225);
nand U27430 (N_27430,N_27055,N_27054);
nand U27431 (N_27431,N_27222,N_27199);
nand U27432 (N_27432,N_27296,N_27087);
and U27433 (N_27433,N_27135,N_27011);
or U27434 (N_27434,N_27188,N_27107);
nor U27435 (N_27435,N_27022,N_27297);
nor U27436 (N_27436,N_27292,N_27153);
nor U27437 (N_27437,N_27243,N_27006);
and U27438 (N_27438,N_27105,N_27267);
or U27439 (N_27439,N_27215,N_27242);
or U27440 (N_27440,N_27151,N_27095);
xor U27441 (N_27441,N_27245,N_27194);
xor U27442 (N_27442,N_27237,N_27047);
xor U27443 (N_27443,N_27008,N_27294);
or U27444 (N_27444,N_27166,N_27147);
xnor U27445 (N_27445,N_27168,N_27202);
nand U27446 (N_27446,N_27191,N_27208);
nor U27447 (N_27447,N_27173,N_27280);
or U27448 (N_27448,N_27288,N_27252);
and U27449 (N_27449,N_27079,N_27109);
or U27450 (N_27450,N_27082,N_27198);
xnor U27451 (N_27451,N_27076,N_27221);
nor U27452 (N_27452,N_27121,N_27043);
nor U27453 (N_27453,N_27252,N_27193);
nor U27454 (N_27454,N_27179,N_27146);
nand U27455 (N_27455,N_27159,N_27086);
or U27456 (N_27456,N_27108,N_27032);
nor U27457 (N_27457,N_27035,N_27014);
nand U27458 (N_27458,N_27124,N_27169);
nor U27459 (N_27459,N_27207,N_27298);
nor U27460 (N_27460,N_27281,N_27139);
or U27461 (N_27461,N_27002,N_27293);
nand U27462 (N_27462,N_27087,N_27098);
nor U27463 (N_27463,N_27066,N_27154);
nand U27464 (N_27464,N_27195,N_27185);
xor U27465 (N_27465,N_27224,N_27290);
nor U27466 (N_27466,N_27070,N_27142);
or U27467 (N_27467,N_27116,N_27064);
nor U27468 (N_27468,N_27108,N_27298);
xnor U27469 (N_27469,N_27143,N_27114);
or U27470 (N_27470,N_27143,N_27253);
nor U27471 (N_27471,N_27094,N_27056);
or U27472 (N_27472,N_27260,N_27212);
nor U27473 (N_27473,N_27051,N_27012);
nor U27474 (N_27474,N_27179,N_27240);
or U27475 (N_27475,N_27278,N_27125);
xor U27476 (N_27476,N_27169,N_27242);
nand U27477 (N_27477,N_27233,N_27076);
nand U27478 (N_27478,N_27049,N_27256);
nor U27479 (N_27479,N_27167,N_27243);
nor U27480 (N_27480,N_27127,N_27164);
and U27481 (N_27481,N_27197,N_27036);
nand U27482 (N_27482,N_27273,N_27126);
nor U27483 (N_27483,N_27266,N_27101);
or U27484 (N_27484,N_27148,N_27107);
nor U27485 (N_27485,N_27159,N_27089);
or U27486 (N_27486,N_27245,N_27230);
nor U27487 (N_27487,N_27021,N_27158);
and U27488 (N_27488,N_27197,N_27002);
and U27489 (N_27489,N_27230,N_27244);
and U27490 (N_27490,N_27097,N_27155);
xnor U27491 (N_27491,N_27282,N_27043);
nand U27492 (N_27492,N_27036,N_27035);
nand U27493 (N_27493,N_27284,N_27175);
and U27494 (N_27494,N_27058,N_27059);
and U27495 (N_27495,N_27044,N_27040);
or U27496 (N_27496,N_27034,N_27234);
nor U27497 (N_27497,N_27134,N_27189);
nand U27498 (N_27498,N_27162,N_27028);
xor U27499 (N_27499,N_27029,N_27212);
nand U27500 (N_27500,N_27047,N_27126);
or U27501 (N_27501,N_27233,N_27200);
nor U27502 (N_27502,N_27216,N_27173);
xnor U27503 (N_27503,N_27262,N_27216);
or U27504 (N_27504,N_27109,N_27074);
and U27505 (N_27505,N_27100,N_27141);
xnor U27506 (N_27506,N_27099,N_27151);
nand U27507 (N_27507,N_27040,N_27097);
nor U27508 (N_27508,N_27185,N_27220);
xnor U27509 (N_27509,N_27141,N_27200);
and U27510 (N_27510,N_27208,N_27033);
nand U27511 (N_27511,N_27273,N_27014);
nand U27512 (N_27512,N_27095,N_27154);
nor U27513 (N_27513,N_27236,N_27035);
nand U27514 (N_27514,N_27194,N_27216);
nor U27515 (N_27515,N_27166,N_27038);
and U27516 (N_27516,N_27127,N_27054);
xor U27517 (N_27517,N_27125,N_27095);
xor U27518 (N_27518,N_27220,N_27150);
nand U27519 (N_27519,N_27112,N_27292);
or U27520 (N_27520,N_27122,N_27105);
nor U27521 (N_27521,N_27227,N_27140);
xor U27522 (N_27522,N_27207,N_27156);
nor U27523 (N_27523,N_27147,N_27177);
nor U27524 (N_27524,N_27237,N_27094);
or U27525 (N_27525,N_27229,N_27137);
nand U27526 (N_27526,N_27154,N_27013);
nand U27527 (N_27527,N_27059,N_27248);
or U27528 (N_27528,N_27063,N_27120);
xor U27529 (N_27529,N_27052,N_27241);
and U27530 (N_27530,N_27109,N_27296);
nor U27531 (N_27531,N_27219,N_27295);
nand U27532 (N_27532,N_27184,N_27130);
nand U27533 (N_27533,N_27112,N_27046);
or U27534 (N_27534,N_27153,N_27023);
and U27535 (N_27535,N_27044,N_27240);
or U27536 (N_27536,N_27210,N_27184);
and U27537 (N_27537,N_27168,N_27286);
xor U27538 (N_27538,N_27243,N_27146);
and U27539 (N_27539,N_27226,N_27167);
or U27540 (N_27540,N_27263,N_27205);
nor U27541 (N_27541,N_27058,N_27089);
nand U27542 (N_27542,N_27088,N_27277);
or U27543 (N_27543,N_27208,N_27254);
and U27544 (N_27544,N_27210,N_27061);
and U27545 (N_27545,N_27115,N_27291);
nand U27546 (N_27546,N_27298,N_27132);
or U27547 (N_27547,N_27053,N_27161);
xor U27548 (N_27548,N_27124,N_27234);
xor U27549 (N_27549,N_27073,N_27050);
nand U27550 (N_27550,N_27244,N_27063);
nand U27551 (N_27551,N_27159,N_27098);
xor U27552 (N_27552,N_27194,N_27284);
xor U27553 (N_27553,N_27158,N_27201);
nand U27554 (N_27554,N_27034,N_27173);
xor U27555 (N_27555,N_27122,N_27042);
xor U27556 (N_27556,N_27120,N_27075);
nor U27557 (N_27557,N_27299,N_27138);
nor U27558 (N_27558,N_27072,N_27183);
or U27559 (N_27559,N_27227,N_27111);
or U27560 (N_27560,N_27224,N_27173);
nor U27561 (N_27561,N_27070,N_27263);
and U27562 (N_27562,N_27038,N_27199);
or U27563 (N_27563,N_27219,N_27200);
and U27564 (N_27564,N_27258,N_27011);
nor U27565 (N_27565,N_27161,N_27275);
or U27566 (N_27566,N_27086,N_27239);
nand U27567 (N_27567,N_27153,N_27035);
xor U27568 (N_27568,N_27159,N_27264);
xnor U27569 (N_27569,N_27100,N_27142);
nor U27570 (N_27570,N_27030,N_27130);
nor U27571 (N_27571,N_27151,N_27152);
and U27572 (N_27572,N_27151,N_27145);
nor U27573 (N_27573,N_27224,N_27104);
xor U27574 (N_27574,N_27111,N_27279);
and U27575 (N_27575,N_27097,N_27026);
nor U27576 (N_27576,N_27080,N_27180);
and U27577 (N_27577,N_27039,N_27238);
nor U27578 (N_27578,N_27053,N_27020);
xor U27579 (N_27579,N_27134,N_27008);
nor U27580 (N_27580,N_27139,N_27188);
or U27581 (N_27581,N_27258,N_27085);
xor U27582 (N_27582,N_27276,N_27092);
nand U27583 (N_27583,N_27196,N_27224);
and U27584 (N_27584,N_27124,N_27179);
and U27585 (N_27585,N_27006,N_27110);
nand U27586 (N_27586,N_27001,N_27270);
nand U27587 (N_27587,N_27159,N_27039);
and U27588 (N_27588,N_27045,N_27061);
nor U27589 (N_27589,N_27254,N_27083);
nor U27590 (N_27590,N_27270,N_27294);
nor U27591 (N_27591,N_27138,N_27036);
nor U27592 (N_27592,N_27220,N_27009);
or U27593 (N_27593,N_27087,N_27115);
nor U27594 (N_27594,N_27214,N_27100);
xnor U27595 (N_27595,N_27288,N_27025);
or U27596 (N_27596,N_27268,N_27088);
or U27597 (N_27597,N_27181,N_27290);
nor U27598 (N_27598,N_27199,N_27057);
nand U27599 (N_27599,N_27295,N_27128);
nor U27600 (N_27600,N_27350,N_27375);
nand U27601 (N_27601,N_27589,N_27318);
and U27602 (N_27602,N_27416,N_27396);
nor U27603 (N_27603,N_27307,N_27436);
nand U27604 (N_27604,N_27370,N_27344);
xnor U27605 (N_27605,N_27486,N_27468);
or U27606 (N_27606,N_27551,N_27517);
and U27607 (N_27607,N_27553,N_27478);
and U27608 (N_27608,N_27431,N_27395);
nor U27609 (N_27609,N_27561,N_27479);
xnor U27610 (N_27610,N_27536,N_27335);
and U27611 (N_27611,N_27562,N_27348);
or U27612 (N_27612,N_27456,N_27437);
xnor U27613 (N_27613,N_27461,N_27360);
nand U27614 (N_27614,N_27550,N_27484);
nor U27615 (N_27615,N_27342,N_27546);
and U27616 (N_27616,N_27330,N_27398);
and U27617 (N_27617,N_27412,N_27469);
or U27618 (N_27618,N_27378,N_27414);
nand U27619 (N_27619,N_27343,N_27497);
nand U27620 (N_27620,N_27397,N_27331);
nor U27621 (N_27621,N_27582,N_27539);
nand U27622 (N_27622,N_27579,N_27376);
nand U27623 (N_27623,N_27495,N_27522);
or U27624 (N_27624,N_27424,N_27560);
or U27625 (N_27625,N_27555,N_27568);
nand U27626 (N_27626,N_27598,N_27512);
or U27627 (N_27627,N_27308,N_27459);
xnor U27628 (N_27628,N_27453,N_27518);
nor U27629 (N_27629,N_27314,N_27520);
xor U27630 (N_27630,N_27305,N_27439);
xor U27631 (N_27631,N_27340,N_27463);
or U27632 (N_27632,N_27316,N_27445);
or U27633 (N_27633,N_27557,N_27429);
nand U27634 (N_27634,N_27441,N_27574);
xor U27635 (N_27635,N_27361,N_27403);
xor U27636 (N_27636,N_27473,N_27324);
and U27637 (N_27637,N_27580,N_27417);
or U27638 (N_27638,N_27339,N_27571);
nand U27639 (N_27639,N_27465,N_27491);
nor U27640 (N_27640,N_27500,N_27438);
nor U27641 (N_27641,N_27559,N_27482);
or U27642 (N_27642,N_27504,N_27362);
or U27643 (N_27643,N_27509,N_27508);
or U27644 (N_27644,N_27368,N_27547);
or U27645 (N_27645,N_27379,N_27367);
and U27646 (N_27646,N_27531,N_27443);
xor U27647 (N_27647,N_27496,N_27347);
or U27648 (N_27648,N_27444,N_27467);
and U27649 (N_27649,N_27385,N_27351);
nor U27650 (N_27650,N_27426,N_27599);
and U27651 (N_27651,N_27353,N_27399);
and U27652 (N_27652,N_27538,N_27516);
nand U27653 (N_27653,N_27534,N_27489);
and U27654 (N_27654,N_27358,N_27471);
or U27655 (N_27655,N_27355,N_27503);
or U27656 (N_27656,N_27329,N_27383);
nor U27657 (N_27657,N_27597,N_27460);
and U27658 (N_27658,N_27388,N_27513);
nand U27659 (N_27659,N_27446,N_27333);
and U27660 (N_27660,N_27573,N_27594);
nand U27661 (N_27661,N_27498,N_27413);
and U27662 (N_27662,N_27541,N_27457);
or U27663 (N_27663,N_27514,N_27476);
xnor U27664 (N_27664,N_27591,N_27549);
xnor U27665 (N_27665,N_27556,N_27451);
and U27666 (N_27666,N_27359,N_27499);
and U27667 (N_27667,N_27535,N_27302);
and U27668 (N_27668,N_27410,N_27366);
nand U27669 (N_27669,N_27328,N_27435);
and U27670 (N_27670,N_27406,N_27381);
and U27671 (N_27671,N_27474,N_27587);
nand U27672 (N_27672,N_27391,N_27552);
xor U27673 (N_27673,N_27427,N_27583);
and U27674 (N_27674,N_27332,N_27543);
or U27675 (N_27675,N_27554,N_27458);
xnor U27676 (N_27676,N_27593,N_27525);
nor U27677 (N_27677,N_27405,N_27304);
and U27678 (N_27678,N_27402,N_27558);
nor U27679 (N_27679,N_27390,N_27354);
nand U27680 (N_27680,N_27317,N_27450);
or U27681 (N_27681,N_27528,N_27430);
and U27682 (N_27682,N_27336,N_27372);
and U27683 (N_27683,N_27510,N_27448);
nor U27684 (N_27684,N_27357,N_27346);
or U27685 (N_27685,N_27581,N_27481);
and U27686 (N_27686,N_27565,N_27519);
nand U27687 (N_27687,N_27363,N_27407);
nor U27688 (N_27688,N_27452,N_27483);
xor U27689 (N_27689,N_27488,N_27349);
nor U27690 (N_27690,N_27433,N_27400);
and U27691 (N_27691,N_27327,N_27529);
xor U27692 (N_27692,N_27309,N_27596);
xnor U27693 (N_27693,N_27530,N_27592);
or U27694 (N_27694,N_27373,N_27411);
xor U27695 (N_27695,N_27315,N_27454);
nor U27696 (N_27696,N_27423,N_27544);
xor U27697 (N_27697,N_27477,N_27590);
and U27698 (N_27698,N_27401,N_27566);
nor U27699 (N_27699,N_27532,N_27303);
and U27700 (N_27700,N_27409,N_27321);
or U27701 (N_27701,N_27382,N_27404);
or U27702 (N_27702,N_27466,N_27319);
nand U27703 (N_27703,N_27511,N_27480);
xnor U27704 (N_27704,N_27575,N_27523);
or U27705 (N_27705,N_27386,N_27310);
and U27706 (N_27706,N_27485,N_27365);
or U27707 (N_27707,N_27364,N_27595);
nand U27708 (N_27708,N_27420,N_27493);
or U27709 (N_27709,N_27501,N_27537);
and U27710 (N_27710,N_27415,N_27301);
nand U27711 (N_27711,N_27462,N_27564);
nor U27712 (N_27712,N_27392,N_27322);
xnor U27713 (N_27713,N_27313,N_27325);
nor U27714 (N_27714,N_27380,N_27506);
nor U27715 (N_27715,N_27369,N_27428);
nand U27716 (N_27716,N_27408,N_27578);
or U27717 (N_27717,N_27584,N_27371);
nor U27718 (N_27718,N_27312,N_27341);
and U27719 (N_27719,N_27545,N_27533);
nor U27720 (N_27720,N_27492,N_27338);
and U27721 (N_27721,N_27393,N_27425);
xor U27722 (N_27722,N_27548,N_27394);
nand U27723 (N_27723,N_27337,N_27323);
xor U27724 (N_27724,N_27515,N_27389);
or U27725 (N_27725,N_27387,N_27311);
nor U27726 (N_27726,N_27526,N_27563);
and U27727 (N_27727,N_27569,N_27356);
and U27728 (N_27728,N_27334,N_27524);
or U27729 (N_27729,N_27490,N_27494);
or U27730 (N_27730,N_27505,N_27374);
nand U27731 (N_27731,N_27464,N_27326);
nor U27732 (N_27732,N_27572,N_27577);
nand U27733 (N_27733,N_27527,N_27487);
and U27734 (N_27734,N_27567,N_27475);
or U27735 (N_27735,N_27418,N_27449);
nand U27736 (N_27736,N_27434,N_27576);
xnor U27737 (N_27737,N_27419,N_27300);
and U27738 (N_27738,N_27306,N_27345);
nand U27739 (N_27739,N_27442,N_27542);
and U27740 (N_27740,N_27455,N_27440);
nor U27741 (N_27741,N_27320,N_27352);
nand U27742 (N_27742,N_27585,N_27432);
nand U27743 (N_27743,N_27507,N_27570);
or U27744 (N_27744,N_27421,N_27377);
and U27745 (N_27745,N_27470,N_27540);
nor U27746 (N_27746,N_27586,N_27502);
nor U27747 (N_27747,N_27521,N_27588);
nand U27748 (N_27748,N_27447,N_27472);
nor U27749 (N_27749,N_27384,N_27422);
nor U27750 (N_27750,N_27385,N_27556);
and U27751 (N_27751,N_27552,N_27383);
xnor U27752 (N_27752,N_27413,N_27400);
nor U27753 (N_27753,N_27403,N_27383);
xor U27754 (N_27754,N_27375,N_27447);
nand U27755 (N_27755,N_27403,N_27534);
or U27756 (N_27756,N_27367,N_27443);
and U27757 (N_27757,N_27316,N_27463);
or U27758 (N_27758,N_27567,N_27324);
nand U27759 (N_27759,N_27355,N_27582);
or U27760 (N_27760,N_27474,N_27487);
nor U27761 (N_27761,N_27497,N_27394);
xor U27762 (N_27762,N_27477,N_27496);
and U27763 (N_27763,N_27370,N_27358);
xor U27764 (N_27764,N_27595,N_27462);
xnor U27765 (N_27765,N_27458,N_27586);
xnor U27766 (N_27766,N_27412,N_27428);
and U27767 (N_27767,N_27534,N_27487);
xnor U27768 (N_27768,N_27367,N_27534);
nand U27769 (N_27769,N_27505,N_27395);
nand U27770 (N_27770,N_27521,N_27327);
xnor U27771 (N_27771,N_27500,N_27421);
nand U27772 (N_27772,N_27435,N_27552);
and U27773 (N_27773,N_27599,N_27557);
or U27774 (N_27774,N_27405,N_27520);
nand U27775 (N_27775,N_27530,N_27421);
xnor U27776 (N_27776,N_27561,N_27566);
xor U27777 (N_27777,N_27566,N_27390);
or U27778 (N_27778,N_27470,N_27554);
or U27779 (N_27779,N_27516,N_27337);
and U27780 (N_27780,N_27523,N_27579);
xor U27781 (N_27781,N_27389,N_27560);
nand U27782 (N_27782,N_27429,N_27384);
xnor U27783 (N_27783,N_27487,N_27513);
nand U27784 (N_27784,N_27369,N_27303);
xnor U27785 (N_27785,N_27582,N_27388);
nor U27786 (N_27786,N_27339,N_27508);
and U27787 (N_27787,N_27530,N_27476);
nand U27788 (N_27788,N_27567,N_27513);
and U27789 (N_27789,N_27328,N_27572);
xor U27790 (N_27790,N_27347,N_27580);
nand U27791 (N_27791,N_27478,N_27393);
or U27792 (N_27792,N_27487,N_27574);
or U27793 (N_27793,N_27552,N_27397);
nand U27794 (N_27794,N_27465,N_27574);
or U27795 (N_27795,N_27396,N_27459);
and U27796 (N_27796,N_27312,N_27585);
nor U27797 (N_27797,N_27533,N_27404);
and U27798 (N_27798,N_27592,N_27439);
nor U27799 (N_27799,N_27530,N_27383);
nand U27800 (N_27800,N_27514,N_27322);
and U27801 (N_27801,N_27328,N_27590);
xor U27802 (N_27802,N_27431,N_27422);
nor U27803 (N_27803,N_27390,N_27527);
nand U27804 (N_27804,N_27448,N_27541);
or U27805 (N_27805,N_27522,N_27316);
nor U27806 (N_27806,N_27387,N_27526);
nor U27807 (N_27807,N_27331,N_27407);
or U27808 (N_27808,N_27496,N_27388);
or U27809 (N_27809,N_27432,N_27530);
nand U27810 (N_27810,N_27598,N_27439);
nor U27811 (N_27811,N_27461,N_27401);
nor U27812 (N_27812,N_27364,N_27381);
and U27813 (N_27813,N_27553,N_27317);
nor U27814 (N_27814,N_27411,N_27353);
nand U27815 (N_27815,N_27415,N_27426);
nand U27816 (N_27816,N_27316,N_27430);
or U27817 (N_27817,N_27567,N_27314);
xor U27818 (N_27818,N_27379,N_27358);
and U27819 (N_27819,N_27476,N_27523);
xor U27820 (N_27820,N_27419,N_27577);
nand U27821 (N_27821,N_27553,N_27565);
and U27822 (N_27822,N_27432,N_27570);
and U27823 (N_27823,N_27507,N_27558);
nand U27824 (N_27824,N_27419,N_27552);
or U27825 (N_27825,N_27567,N_27345);
or U27826 (N_27826,N_27320,N_27588);
nand U27827 (N_27827,N_27593,N_27339);
or U27828 (N_27828,N_27355,N_27440);
or U27829 (N_27829,N_27324,N_27393);
nor U27830 (N_27830,N_27428,N_27333);
and U27831 (N_27831,N_27548,N_27318);
or U27832 (N_27832,N_27594,N_27360);
or U27833 (N_27833,N_27557,N_27519);
or U27834 (N_27834,N_27580,N_27534);
xor U27835 (N_27835,N_27405,N_27556);
and U27836 (N_27836,N_27305,N_27594);
nor U27837 (N_27837,N_27429,N_27376);
or U27838 (N_27838,N_27459,N_27397);
and U27839 (N_27839,N_27432,N_27430);
xor U27840 (N_27840,N_27390,N_27305);
or U27841 (N_27841,N_27378,N_27471);
nor U27842 (N_27842,N_27592,N_27341);
or U27843 (N_27843,N_27518,N_27370);
and U27844 (N_27844,N_27408,N_27548);
nor U27845 (N_27845,N_27598,N_27551);
nand U27846 (N_27846,N_27501,N_27394);
xor U27847 (N_27847,N_27471,N_27496);
nor U27848 (N_27848,N_27408,N_27308);
nor U27849 (N_27849,N_27386,N_27462);
nand U27850 (N_27850,N_27469,N_27339);
and U27851 (N_27851,N_27387,N_27584);
nand U27852 (N_27852,N_27420,N_27406);
and U27853 (N_27853,N_27325,N_27508);
xor U27854 (N_27854,N_27447,N_27539);
nor U27855 (N_27855,N_27442,N_27351);
nor U27856 (N_27856,N_27484,N_27347);
xnor U27857 (N_27857,N_27531,N_27487);
nor U27858 (N_27858,N_27492,N_27429);
nor U27859 (N_27859,N_27508,N_27531);
nand U27860 (N_27860,N_27388,N_27446);
or U27861 (N_27861,N_27423,N_27394);
or U27862 (N_27862,N_27411,N_27365);
xnor U27863 (N_27863,N_27459,N_27475);
or U27864 (N_27864,N_27533,N_27408);
nand U27865 (N_27865,N_27532,N_27393);
xnor U27866 (N_27866,N_27473,N_27500);
and U27867 (N_27867,N_27302,N_27439);
and U27868 (N_27868,N_27343,N_27336);
and U27869 (N_27869,N_27589,N_27314);
and U27870 (N_27870,N_27321,N_27566);
xnor U27871 (N_27871,N_27336,N_27447);
nor U27872 (N_27872,N_27338,N_27543);
or U27873 (N_27873,N_27326,N_27420);
and U27874 (N_27874,N_27495,N_27357);
nor U27875 (N_27875,N_27449,N_27520);
xor U27876 (N_27876,N_27413,N_27556);
xnor U27877 (N_27877,N_27551,N_27323);
nand U27878 (N_27878,N_27337,N_27317);
xnor U27879 (N_27879,N_27576,N_27410);
and U27880 (N_27880,N_27428,N_27306);
or U27881 (N_27881,N_27564,N_27446);
or U27882 (N_27882,N_27495,N_27523);
xor U27883 (N_27883,N_27408,N_27575);
or U27884 (N_27884,N_27594,N_27434);
nor U27885 (N_27885,N_27487,N_27500);
or U27886 (N_27886,N_27385,N_27329);
xnor U27887 (N_27887,N_27535,N_27594);
and U27888 (N_27888,N_27391,N_27591);
nand U27889 (N_27889,N_27574,N_27568);
or U27890 (N_27890,N_27303,N_27365);
and U27891 (N_27891,N_27384,N_27446);
nand U27892 (N_27892,N_27485,N_27304);
and U27893 (N_27893,N_27501,N_27448);
and U27894 (N_27894,N_27306,N_27500);
nor U27895 (N_27895,N_27351,N_27492);
nor U27896 (N_27896,N_27342,N_27307);
nand U27897 (N_27897,N_27370,N_27504);
and U27898 (N_27898,N_27412,N_27414);
or U27899 (N_27899,N_27334,N_27536);
or U27900 (N_27900,N_27689,N_27722);
and U27901 (N_27901,N_27863,N_27801);
and U27902 (N_27902,N_27843,N_27797);
or U27903 (N_27903,N_27852,N_27693);
xor U27904 (N_27904,N_27826,N_27653);
or U27905 (N_27905,N_27765,N_27790);
nor U27906 (N_27906,N_27870,N_27887);
xnor U27907 (N_27907,N_27636,N_27720);
or U27908 (N_27908,N_27794,N_27782);
nand U27909 (N_27909,N_27638,N_27710);
or U27910 (N_27910,N_27777,N_27877);
xnor U27911 (N_27911,N_27847,N_27833);
nor U27912 (N_27912,N_27651,N_27813);
or U27913 (N_27913,N_27775,N_27652);
and U27914 (N_27914,N_27807,N_27809);
nor U27915 (N_27915,N_27889,N_27711);
and U27916 (N_27916,N_27642,N_27654);
nor U27917 (N_27917,N_27845,N_27754);
and U27918 (N_27918,N_27612,N_27672);
nand U27919 (N_27919,N_27763,N_27753);
nor U27920 (N_27920,N_27671,N_27627);
nor U27921 (N_27921,N_27674,N_27610);
nor U27922 (N_27922,N_27882,N_27861);
xor U27923 (N_27923,N_27675,N_27886);
nand U27924 (N_27924,N_27781,N_27773);
or U27925 (N_27925,N_27669,N_27729);
xor U27926 (N_27926,N_27602,N_27623);
or U27927 (N_27927,N_27832,N_27684);
nor U27928 (N_27928,N_27855,N_27740);
xnor U27929 (N_27929,N_27876,N_27734);
and U27930 (N_27930,N_27766,N_27819);
nand U27931 (N_27931,N_27772,N_27691);
and U27932 (N_27932,N_27696,N_27851);
and U27933 (N_27933,N_27685,N_27834);
or U27934 (N_27934,N_27897,N_27838);
nor U27935 (N_27935,N_27830,N_27702);
nand U27936 (N_27936,N_27787,N_27725);
and U27937 (N_27937,N_27622,N_27835);
nor U27938 (N_27938,N_27893,N_27601);
xnor U27939 (N_27939,N_27774,N_27755);
or U27940 (N_27940,N_27697,N_27871);
nor U27941 (N_27941,N_27665,N_27785);
and U27942 (N_27942,N_27824,N_27837);
nand U27943 (N_27943,N_27733,N_27600);
xor U27944 (N_27944,N_27780,N_27706);
or U27945 (N_27945,N_27692,N_27761);
or U27946 (N_27946,N_27898,N_27786);
and U27947 (N_27947,N_27816,N_27853);
nand U27948 (N_27948,N_27791,N_27655);
nor U27949 (N_27949,N_27858,N_27730);
nand U27950 (N_27950,N_27822,N_27737);
xnor U27951 (N_27951,N_27707,N_27621);
or U27952 (N_27952,N_27817,N_27603);
nand U27953 (N_27953,N_27727,N_27724);
or U27954 (N_27954,N_27634,N_27798);
nand U27955 (N_27955,N_27803,N_27842);
xnor U27956 (N_27956,N_27840,N_27821);
or U27957 (N_27957,N_27703,N_27649);
and U27958 (N_27958,N_27614,N_27644);
xnor U27959 (N_27959,N_27872,N_27629);
nor U27960 (N_27960,N_27645,N_27613);
xor U27961 (N_27961,N_27860,N_27681);
or U27962 (N_27962,N_27701,N_27869);
nor U27963 (N_27963,N_27704,N_27719);
and U27964 (N_27964,N_27770,N_27618);
nand U27965 (N_27965,N_27750,N_27836);
nor U27966 (N_27966,N_27687,N_27815);
nand U27967 (N_27967,N_27769,N_27757);
nand U27968 (N_27968,N_27828,N_27866);
or U27969 (N_27969,N_27633,N_27616);
nor U27970 (N_27970,N_27605,N_27732);
or U27971 (N_27971,N_27611,N_27690);
or U27972 (N_27972,N_27742,N_27749);
nor U27973 (N_27973,N_27714,N_27812);
and U27974 (N_27974,N_27746,N_27660);
xor U27975 (N_27975,N_27667,N_27678);
and U27976 (N_27976,N_27796,N_27670);
xor U27977 (N_27977,N_27844,N_27609);
or U27978 (N_27978,N_27850,N_27745);
nand U27979 (N_27979,N_27762,N_27771);
nand U27980 (N_27980,N_27888,N_27625);
nand U27981 (N_27981,N_27626,N_27677);
and U27982 (N_27982,N_27839,N_27736);
or U27983 (N_27983,N_27874,N_27890);
nor U27984 (N_27984,N_27825,N_27668);
or U27985 (N_27985,N_27641,N_27880);
nand U27986 (N_27986,N_27718,N_27873);
or U27987 (N_27987,N_27778,N_27799);
nand U27988 (N_27988,N_27841,N_27747);
or U27989 (N_27989,N_27628,N_27883);
and U27990 (N_27990,N_27806,N_27680);
nand U27991 (N_27991,N_27862,N_27639);
nand U27992 (N_27992,N_27808,N_27864);
nand U27993 (N_27993,N_27606,N_27624);
xnor U27994 (N_27994,N_27751,N_27615);
nor U27995 (N_27995,N_27617,N_27741);
and U27996 (N_27996,N_27676,N_27712);
or U27997 (N_27997,N_27632,N_27752);
nand U27998 (N_27998,N_27739,N_27859);
nor U27999 (N_27999,N_27744,N_27683);
nor U28000 (N_28000,N_27865,N_27695);
nor U28001 (N_28001,N_27640,N_27726);
and U28002 (N_28002,N_27648,N_27848);
nand U28003 (N_28003,N_27708,N_27656);
or U28004 (N_28004,N_27875,N_27878);
or U28005 (N_28005,N_27607,N_27810);
nor U28006 (N_28006,N_27802,N_27779);
and U28007 (N_28007,N_27795,N_27716);
and U28008 (N_28008,N_27658,N_27688);
nand U28009 (N_28009,N_27659,N_27760);
nor U28010 (N_28010,N_27879,N_27679);
nand U28011 (N_28011,N_27756,N_27831);
or U28012 (N_28012,N_27792,N_27804);
xor U28013 (N_28013,N_27788,N_27743);
nor U28014 (N_28014,N_27620,N_27846);
nand U28015 (N_28015,N_27764,N_27814);
nor U28016 (N_28016,N_27604,N_27827);
or U28017 (N_28017,N_27818,N_27715);
nand U28018 (N_28018,N_27784,N_27661);
or U28019 (N_28019,N_27666,N_27698);
nor U28020 (N_28020,N_27643,N_27705);
and U28021 (N_28021,N_27635,N_27776);
nand U28022 (N_28022,N_27728,N_27896);
nor U28023 (N_28023,N_27738,N_27686);
xor U28024 (N_28024,N_27823,N_27673);
nor U28025 (N_28025,N_27857,N_27713);
and U28026 (N_28026,N_27881,N_27721);
xor U28027 (N_28027,N_27892,N_27789);
xnor U28028 (N_28028,N_27868,N_27650);
and U28029 (N_28029,N_27664,N_27699);
and U28030 (N_28030,N_27891,N_27748);
nor U28031 (N_28031,N_27856,N_27805);
xor U28032 (N_28032,N_27717,N_27630);
and U28033 (N_28033,N_27884,N_27608);
or U28034 (N_28034,N_27854,N_27662);
and U28035 (N_28035,N_27829,N_27758);
and U28036 (N_28036,N_27631,N_27849);
nor U28037 (N_28037,N_27767,N_27894);
xnor U28038 (N_28038,N_27709,N_27647);
and U28039 (N_28039,N_27682,N_27731);
nand U28040 (N_28040,N_27723,N_27811);
nor U28041 (N_28041,N_27820,N_27619);
nor U28042 (N_28042,N_27759,N_27700);
xnor U28043 (N_28043,N_27735,N_27783);
and U28044 (N_28044,N_27663,N_27899);
and U28045 (N_28045,N_27867,N_27768);
or U28046 (N_28046,N_27657,N_27885);
nand U28047 (N_28047,N_27646,N_27895);
xnor U28048 (N_28048,N_27793,N_27637);
or U28049 (N_28049,N_27800,N_27694);
xnor U28050 (N_28050,N_27845,N_27745);
nand U28051 (N_28051,N_27754,N_27810);
or U28052 (N_28052,N_27604,N_27668);
or U28053 (N_28053,N_27816,N_27767);
nor U28054 (N_28054,N_27858,N_27617);
xnor U28055 (N_28055,N_27804,N_27605);
and U28056 (N_28056,N_27885,N_27621);
xor U28057 (N_28057,N_27770,N_27765);
or U28058 (N_28058,N_27664,N_27607);
nand U28059 (N_28059,N_27898,N_27865);
nor U28060 (N_28060,N_27705,N_27792);
xor U28061 (N_28061,N_27744,N_27834);
xor U28062 (N_28062,N_27655,N_27649);
or U28063 (N_28063,N_27754,N_27777);
or U28064 (N_28064,N_27715,N_27887);
and U28065 (N_28065,N_27798,N_27698);
nor U28066 (N_28066,N_27896,N_27788);
xnor U28067 (N_28067,N_27763,N_27871);
nand U28068 (N_28068,N_27798,N_27789);
and U28069 (N_28069,N_27622,N_27645);
nand U28070 (N_28070,N_27892,N_27841);
xnor U28071 (N_28071,N_27812,N_27600);
and U28072 (N_28072,N_27870,N_27698);
and U28073 (N_28073,N_27705,N_27811);
nor U28074 (N_28074,N_27808,N_27788);
and U28075 (N_28075,N_27816,N_27794);
xnor U28076 (N_28076,N_27793,N_27780);
nand U28077 (N_28077,N_27817,N_27706);
and U28078 (N_28078,N_27808,N_27895);
nor U28079 (N_28079,N_27700,N_27866);
and U28080 (N_28080,N_27745,N_27832);
and U28081 (N_28081,N_27779,N_27791);
nand U28082 (N_28082,N_27866,N_27725);
nor U28083 (N_28083,N_27632,N_27747);
xnor U28084 (N_28084,N_27876,N_27765);
xnor U28085 (N_28085,N_27613,N_27825);
and U28086 (N_28086,N_27859,N_27752);
and U28087 (N_28087,N_27735,N_27674);
nor U28088 (N_28088,N_27827,N_27655);
or U28089 (N_28089,N_27700,N_27704);
or U28090 (N_28090,N_27682,N_27816);
nand U28091 (N_28091,N_27803,N_27835);
nor U28092 (N_28092,N_27719,N_27690);
nor U28093 (N_28093,N_27829,N_27713);
nand U28094 (N_28094,N_27641,N_27683);
xnor U28095 (N_28095,N_27660,N_27896);
and U28096 (N_28096,N_27720,N_27806);
nor U28097 (N_28097,N_27655,N_27724);
or U28098 (N_28098,N_27651,N_27750);
and U28099 (N_28099,N_27611,N_27671);
nand U28100 (N_28100,N_27692,N_27807);
and U28101 (N_28101,N_27778,N_27749);
nor U28102 (N_28102,N_27786,N_27677);
nand U28103 (N_28103,N_27755,N_27635);
nor U28104 (N_28104,N_27816,N_27663);
xnor U28105 (N_28105,N_27631,N_27852);
or U28106 (N_28106,N_27731,N_27888);
and U28107 (N_28107,N_27888,N_27898);
nor U28108 (N_28108,N_27891,N_27602);
and U28109 (N_28109,N_27776,N_27664);
or U28110 (N_28110,N_27607,N_27651);
xnor U28111 (N_28111,N_27632,N_27634);
and U28112 (N_28112,N_27852,N_27735);
and U28113 (N_28113,N_27713,N_27680);
xnor U28114 (N_28114,N_27838,N_27784);
nand U28115 (N_28115,N_27658,N_27824);
xor U28116 (N_28116,N_27844,N_27855);
nor U28117 (N_28117,N_27795,N_27656);
or U28118 (N_28118,N_27819,N_27873);
nand U28119 (N_28119,N_27615,N_27771);
and U28120 (N_28120,N_27866,N_27616);
or U28121 (N_28121,N_27838,N_27608);
and U28122 (N_28122,N_27643,N_27660);
nand U28123 (N_28123,N_27864,N_27730);
nand U28124 (N_28124,N_27771,N_27801);
and U28125 (N_28125,N_27747,N_27759);
xor U28126 (N_28126,N_27694,N_27652);
and U28127 (N_28127,N_27890,N_27803);
xor U28128 (N_28128,N_27821,N_27849);
xor U28129 (N_28129,N_27602,N_27862);
nand U28130 (N_28130,N_27779,N_27638);
and U28131 (N_28131,N_27744,N_27718);
xnor U28132 (N_28132,N_27688,N_27836);
xor U28133 (N_28133,N_27773,N_27635);
xnor U28134 (N_28134,N_27695,N_27751);
xor U28135 (N_28135,N_27871,N_27709);
xnor U28136 (N_28136,N_27737,N_27628);
or U28137 (N_28137,N_27638,N_27648);
nor U28138 (N_28138,N_27823,N_27701);
and U28139 (N_28139,N_27615,N_27823);
xor U28140 (N_28140,N_27666,N_27609);
or U28141 (N_28141,N_27788,N_27895);
nor U28142 (N_28142,N_27792,N_27832);
nand U28143 (N_28143,N_27812,N_27803);
nand U28144 (N_28144,N_27806,N_27725);
nor U28145 (N_28145,N_27860,N_27803);
nor U28146 (N_28146,N_27792,N_27819);
xnor U28147 (N_28147,N_27713,N_27693);
or U28148 (N_28148,N_27703,N_27674);
nor U28149 (N_28149,N_27872,N_27709);
or U28150 (N_28150,N_27684,N_27839);
nand U28151 (N_28151,N_27842,N_27677);
and U28152 (N_28152,N_27884,N_27870);
xor U28153 (N_28153,N_27876,N_27610);
nor U28154 (N_28154,N_27888,N_27876);
nand U28155 (N_28155,N_27779,N_27660);
xor U28156 (N_28156,N_27713,N_27716);
and U28157 (N_28157,N_27646,N_27850);
nor U28158 (N_28158,N_27853,N_27689);
nor U28159 (N_28159,N_27803,N_27686);
xor U28160 (N_28160,N_27637,N_27895);
nand U28161 (N_28161,N_27667,N_27688);
nor U28162 (N_28162,N_27702,N_27648);
nor U28163 (N_28163,N_27702,N_27672);
and U28164 (N_28164,N_27644,N_27824);
and U28165 (N_28165,N_27852,N_27879);
xor U28166 (N_28166,N_27834,N_27835);
nand U28167 (N_28167,N_27890,N_27617);
xor U28168 (N_28168,N_27692,N_27659);
and U28169 (N_28169,N_27859,N_27620);
or U28170 (N_28170,N_27708,N_27621);
xor U28171 (N_28171,N_27855,N_27794);
xnor U28172 (N_28172,N_27787,N_27806);
xnor U28173 (N_28173,N_27658,N_27614);
or U28174 (N_28174,N_27753,N_27616);
xor U28175 (N_28175,N_27684,N_27817);
xor U28176 (N_28176,N_27790,N_27633);
nor U28177 (N_28177,N_27617,N_27691);
nor U28178 (N_28178,N_27862,N_27863);
and U28179 (N_28179,N_27739,N_27762);
xor U28180 (N_28180,N_27889,N_27701);
xor U28181 (N_28181,N_27714,N_27793);
nand U28182 (N_28182,N_27691,N_27644);
and U28183 (N_28183,N_27802,N_27754);
nor U28184 (N_28184,N_27678,N_27637);
nand U28185 (N_28185,N_27705,N_27703);
or U28186 (N_28186,N_27634,N_27739);
and U28187 (N_28187,N_27739,N_27832);
or U28188 (N_28188,N_27723,N_27808);
and U28189 (N_28189,N_27641,N_27703);
or U28190 (N_28190,N_27883,N_27640);
and U28191 (N_28191,N_27761,N_27858);
or U28192 (N_28192,N_27600,N_27866);
nand U28193 (N_28193,N_27648,N_27815);
nand U28194 (N_28194,N_27739,N_27870);
nor U28195 (N_28195,N_27726,N_27627);
nand U28196 (N_28196,N_27845,N_27610);
or U28197 (N_28197,N_27725,N_27731);
nand U28198 (N_28198,N_27728,N_27888);
nand U28199 (N_28199,N_27708,N_27814);
xnor U28200 (N_28200,N_28190,N_28065);
nor U28201 (N_28201,N_27937,N_28150);
nor U28202 (N_28202,N_28127,N_28154);
nand U28203 (N_28203,N_28097,N_28178);
and U28204 (N_28204,N_27916,N_28111);
or U28205 (N_28205,N_27917,N_27901);
nor U28206 (N_28206,N_28013,N_28096);
nor U28207 (N_28207,N_28188,N_28018);
nand U28208 (N_28208,N_28109,N_28005);
nor U28209 (N_28209,N_27921,N_28051);
or U28210 (N_28210,N_28172,N_27957);
nand U28211 (N_28211,N_28141,N_28099);
nand U28212 (N_28212,N_28068,N_28126);
and U28213 (N_28213,N_28050,N_28125);
and U28214 (N_28214,N_27965,N_28027);
nand U28215 (N_28215,N_28161,N_28158);
nor U28216 (N_28216,N_28081,N_28070);
nand U28217 (N_28217,N_28010,N_27982);
nand U28218 (N_28218,N_28114,N_28199);
or U28219 (N_28219,N_28057,N_28086);
xor U28220 (N_28220,N_28159,N_28198);
xnor U28221 (N_28221,N_27929,N_28019);
xnor U28222 (N_28222,N_27961,N_27902);
nor U28223 (N_28223,N_27946,N_28148);
nor U28224 (N_28224,N_28045,N_27908);
nor U28225 (N_28225,N_28184,N_28100);
and U28226 (N_28226,N_28082,N_27983);
xor U28227 (N_28227,N_27962,N_28156);
nand U28228 (N_28228,N_28192,N_28144);
nor U28229 (N_28229,N_28007,N_27928);
or U28230 (N_28230,N_28102,N_27927);
and U28231 (N_28231,N_27906,N_28104);
nand U28232 (N_28232,N_28160,N_28056);
and U28233 (N_28233,N_28153,N_28142);
nand U28234 (N_28234,N_27963,N_28146);
and U28235 (N_28235,N_28121,N_28166);
or U28236 (N_28236,N_28077,N_28181);
xor U28237 (N_28237,N_27924,N_28123);
or U28238 (N_28238,N_28042,N_27934);
and U28239 (N_28239,N_27956,N_28066);
and U28240 (N_28240,N_28014,N_28021);
and U28241 (N_28241,N_28179,N_28191);
xnor U28242 (N_28242,N_28006,N_28015);
nor U28243 (N_28243,N_28037,N_27973);
and U28244 (N_28244,N_28175,N_28060);
or U28245 (N_28245,N_28108,N_28106);
nor U28246 (N_28246,N_28038,N_27948);
nand U28247 (N_28247,N_28061,N_28138);
or U28248 (N_28248,N_27967,N_28053);
nand U28249 (N_28249,N_28083,N_27975);
nand U28250 (N_28250,N_27931,N_27964);
nand U28251 (N_28251,N_28117,N_28035);
or U28252 (N_28252,N_27925,N_28147);
and U28253 (N_28253,N_27991,N_28069);
nor U28254 (N_28254,N_27919,N_28196);
nor U28255 (N_28255,N_27920,N_28119);
nand U28256 (N_28256,N_28167,N_28047);
xnor U28257 (N_28257,N_27992,N_27979);
or U28258 (N_28258,N_28101,N_28112);
or U28259 (N_28259,N_28093,N_27996);
nor U28260 (N_28260,N_28054,N_27945);
nor U28261 (N_28261,N_28110,N_28132);
nand U28262 (N_28262,N_28180,N_28091);
xnor U28263 (N_28263,N_28030,N_28094);
nand U28264 (N_28264,N_28124,N_27999);
and U28265 (N_28265,N_27977,N_28187);
nor U28266 (N_28266,N_27985,N_28011);
xor U28267 (N_28267,N_27930,N_27905);
xor U28268 (N_28268,N_28194,N_27938);
xnor U28269 (N_28269,N_27976,N_28195);
or U28270 (N_28270,N_28089,N_28048);
xnor U28271 (N_28271,N_27986,N_27959);
xnor U28272 (N_28272,N_27910,N_27997);
nand U28273 (N_28273,N_28064,N_28088);
xor U28274 (N_28274,N_28028,N_28185);
and U28275 (N_28275,N_27984,N_28118);
xor U28276 (N_28276,N_28165,N_28087);
or U28277 (N_28277,N_28071,N_28197);
nand U28278 (N_28278,N_28063,N_27940);
nor U28279 (N_28279,N_28031,N_28116);
and U28280 (N_28280,N_28043,N_28008);
xnor U28281 (N_28281,N_27918,N_28041);
nor U28282 (N_28282,N_28078,N_28079);
xnor U28283 (N_28283,N_28120,N_27935);
nand U28284 (N_28284,N_27942,N_28134);
and U28285 (N_28285,N_27974,N_27969);
and U28286 (N_28286,N_28036,N_27971);
nand U28287 (N_28287,N_27926,N_27955);
nor U28288 (N_28288,N_28128,N_28052);
nor U28289 (N_28289,N_28107,N_28095);
or U28290 (N_28290,N_27941,N_28177);
xor U28291 (N_28291,N_28169,N_28164);
or U28292 (N_28292,N_28044,N_28189);
or U28293 (N_28293,N_27911,N_28067);
xor U28294 (N_28294,N_28152,N_28136);
nor U28295 (N_28295,N_28129,N_27912);
nor U28296 (N_28296,N_28140,N_28076);
and U28297 (N_28297,N_28105,N_27966);
xnor U28298 (N_28298,N_27990,N_27989);
nand U28299 (N_28299,N_28135,N_28098);
or U28300 (N_28300,N_28039,N_27943);
and U28301 (N_28301,N_28025,N_27904);
nor U28302 (N_28302,N_28168,N_28029);
and U28303 (N_28303,N_28145,N_28151);
xor U28304 (N_28304,N_27987,N_27968);
nand U28305 (N_28305,N_27903,N_28046);
or U28306 (N_28306,N_28170,N_28130);
xor U28307 (N_28307,N_28012,N_28032);
nand U28308 (N_28308,N_28062,N_28020);
nand U28309 (N_28309,N_28004,N_27960);
or U28310 (N_28310,N_28131,N_28072);
nor U28311 (N_28311,N_27932,N_27915);
or U28312 (N_28312,N_27947,N_28193);
nor U28313 (N_28313,N_28000,N_28002);
nand U28314 (N_28314,N_28186,N_28174);
and U28315 (N_28315,N_28090,N_27922);
xor U28316 (N_28316,N_27951,N_27914);
or U28317 (N_28317,N_27953,N_28113);
nor U28318 (N_28318,N_28074,N_28171);
or U28319 (N_28319,N_27936,N_27923);
and U28320 (N_28320,N_28157,N_28162);
or U28321 (N_28321,N_28122,N_28022);
nor U28322 (N_28322,N_27913,N_28023);
nand U28323 (N_28323,N_27950,N_27993);
or U28324 (N_28324,N_27939,N_28173);
nand U28325 (N_28325,N_27981,N_27958);
and U28326 (N_28326,N_27933,N_28080);
xnor U28327 (N_28327,N_28085,N_28026);
or U28328 (N_28328,N_28034,N_27970);
and U28329 (N_28329,N_27907,N_28092);
xor U28330 (N_28330,N_28115,N_27978);
and U28331 (N_28331,N_28059,N_28163);
or U28332 (N_28332,N_28001,N_28182);
nor U28333 (N_28333,N_28017,N_28055);
and U28334 (N_28334,N_28075,N_28049);
xor U28335 (N_28335,N_27944,N_27900);
or U28336 (N_28336,N_28024,N_28103);
nor U28337 (N_28337,N_28133,N_27909);
or U28338 (N_28338,N_28176,N_28016);
nor U28339 (N_28339,N_27954,N_28040);
xor U28340 (N_28340,N_28084,N_28009);
xnor U28341 (N_28341,N_27949,N_28137);
xnor U28342 (N_28342,N_28073,N_27972);
and U28343 (N_28343,N_27995,N_28033);
and U28344 (N_28344,N_27952,N_27980);
xnor U28345 (N_28345,N_27998,N_27988);
xnor U28346 (N_28346,N_28155,N_28003);
nand U28347 (N_28347,N_28058,N_28143);
and U28348 (N_28348,N_28183,N_28149);
or U28349 (N_28349,N_28139,N_27994);
nand U28350 (N_28350,N_28045,N_28125);
or U28351 (N_28351,N_28024,N_28149);
and U28352 (N_28352,N_28113,N_27917);
xnor U28353 (N_28353,N_28139,N_27984);
or U28354 (N_28354,N_28157,N_27978);
or U28355 (N_28355,N_28167,N_28098);
and U28356 (N_28356,N_27938,N_27946);
xor U28357 (N_28357,N_28073,N_28132);
and U28358 (N_28358,N_28024,N_28127);
nand U28359 (N_28359,N_27978,N_27909);
and U28360 (N_28360,N_27995,N_27984);
nor U28361 (N_28361,N_28035,N_28172);
nand U28362 (N_28362,N_28123,N_27979);
nor U28363 (N_28363,N_27916,N_27942);
nand U28364 (N_28364,N_28131,N_28025);
or U28365 (N_28365,N_27981,N_27985);
and U28366 (N_28366,N_28158,N_28057);
nand U28367 (N_28367,N_27951,N_27930);
nor U28368 (N_28368,N_28171,N_28187);
or U28369 (N_28369,N_28180,N_28078);
and U28370 (N_28370,N_28049,N_28106);
nand U28371 (N_28371,N_28071,N_27916);
xor U28372 (N_28372,N_27911,N_27925);
and U28373 (N_28373,N_27989,N_28175);
or U28374 (N_28374,N_28094,N_28117);
nand U28375 (N_28375,N_27919,N_27980);
or U28376 (N_28376,N_27998,N_28085);
nor U28377 (N_28377,N_28036,N_28003);
and U28378 (N_28378,N_28113,N_27926);
nor U28379 (N_28379,N_27947,N_28022);
xnor U28380 (N_28380,N_27946,N_28128);
and U28381 (N_28381,N_28198,N_28055);
xnor U28382 (N_28382,N_28052,N_28106);
nand U28383 (N_28383,N_28102,N_27962);
or U28384 (N_28384,N_28038,N_27933);
or U28385 (N_28385,N_27905,N_28151);
nor U28386 (N_28386,N_28042,N_27903);
nand U28387 (N_28387,N_28031,N_27941);
and U28388 (N_28388,N_28129,N_28115);
or U28389 (N_28389,N_28185,N_27966);
or U28390 (N_28390,N_28127,N_28023);
nand U28391 (N_28391,N_27964,N_28170);
and U28392 (N_28392,N_27993,N_28013);
and U28393 (N_28393,N_28006,N_28165);
and U28394 (N_28394,N_28173,N_28049);
and U28395 (N_28395,N_28172,N_27986);
nand U28396 (N_28396,N_28077,N_28080);
nor U28397 (N_28397,N_27993,N_28136);
xor U28398 (N_28398,N_28127,N_28116);
and U28399 (N_28399,N_28126,N_28098);
and U28400 (N_28400,N_28164,N_28160);
nor U28401 (N_28401,N_28198,N_27986);
nand U28402 (N_28402,N_27995,N_28089);
xor U28403 (N_28403,N_28080,N_28097);
nor U28404 (N_28404,N_28017,N_28076);
xnor U28405 (N_28405,N_27921,N_28053);
xnor U28406 (N_28406,N_28034,N_28058);
nor U28407 (N_28407,N_28102,N_28158);
or U28408 (N_28408,N_28032,N_27957);
and U28409 (N_28409,N_28085,N_27931);
nand U28410 (N_28410,N_28099,N_27925);
nor U28411 (N_28411,N_28043,N_28196);
nand U28412 (N_28412,N_28080,N_28009);
and U28413 (N_28413,N_28139,N_27966);
nor U28414 (N_28414,N_27908,N_28095);
nand U28415 (N_28415,N_28173,N_28006);
nor U28416 (N_28416,N_28084,N_28158);
nand U28417 (N_28417,N_28109,N_27915);
nor U28418 (N_28418,N_28094,N_28037);
and U28419 (N_28419,N_27927,N_28198);
nand U28420 (N_28420,N_28121,N_28102);
or U28421 (N_28421,N_27982,N_28002);
and U28422 (N_28422,N_27987,N_28127);
xnor U28423 (N_28423,N_28108,N_27997);
nand U28424 (N_28424,N_27949,N_27919);
nand U28425 (N_28425,N_28114,N_28189);
nor U28426 (N_28426,N_28043,N_27994);
or U28427 (N_28427,N_28066,N_28057);
or U28428 (N_28428,N_28165,N_28182);
nor U28429 (N_28429,N_28009,N_28136);
nand U28430 (N_28430,N_27932,N_28060);
xnor U28431 (N_28431,N_28073,N_27933);
or U28432 (N_28432,N_28007,N_28184);
or U28433 (N_28433,N_28058,N_28153);
or U28434 (N_28434,N_27973,N_27906);
and U28435 (N_28435,N_28048,N_28172);
xnor U28436 (N_28436,N_27995,N_28035);
xor U28437 (N_28437,N_28112,N_28012);
or U28438 (N_28438,N_28055,N_28093);
and U28439 (N_28439,N_28070,N_28068);
xor U28440 (N_28440,N_27989,N_27941);
nand U28441 (N_28441,N_27922,N_27984);
xnor U28442 (N_28442,N_27982,N_28129);
nand U28443 (N_28443,N_27901,N_28126);
and U28444 (N_28444,N_27932,N_28075);
nor U28445 (N_28445,N_28152,N_28138);
and U28446 (N_28446,N_28082,N_28091);
xnor U28447 (N_28447,N_28161,N_28076);
xnor U28448 (N_28448,N_28098,N_27911);
nand U28449 (N_28449,N_28084,N_27924);
nor U28450 (N_28450,N_28039,N_28163);
nand U28451 (N_28451,N_27976,N_28026);
and U28452 (N_28452,N_27931,N_28141);
or U28453 (N_28453,N_28110,N_28141);
nor U28454 (N_28454,N_28174,N_28120);
nor U28455 (N_28455,N_28033,N_28081);
xnor U28456 (N_28456,N_27973,N_28059);
or U28457 (N_28457,N_27981,N_27943);
or U28458 (N_28458,N_28028,N_28052);
or U28459 (N_28459,N_28176,N_27990);
nand U28460 (N_28460,N_28123,N_28162);
and U28461 (N_28461,N_27948,N_28015);
and U28462 (N_28462,N_27942,N_28117);
xor U28463 (N_28463,N_28081,N_27915);
or U28464 (N_28464,N_28048,N_27966);
and U28465 (N_28465,N_28020,N_28025);
nand U28466 (N_28466,N_28051,N_27967);
or U28467 (N_28467,N_28158,N_28182);
and U28468 (N_28468,N_28007,N_28114);
xor U28469 (N_28469,N_27930,N_28071);
or U28470 (N_28470,N_27952,N_28192);
nand U28471 (N_28471,N_27921,N_28001);
nor U28472 (N_28472,N_28090,N_28116);
nor U28473 (N_28473,N_27960,N_28141);
nand U28474 (N_28474,N_28139,N_28145);
and U28475 (N_28475,N_28087,N_28123);
nor U28476 (N_28476,N_28094,N_28124);
and U28477 (N_28477,N_27929,N_28018);
xnor U28478 (N_28478,N_28087,N_28003);
xnor U28479 (N_28479,N_28065,N_27933);
nor U28480 (N_28480,N_28079,N_28151);
and U28481 (N_28481,N_28037,N_28177);
nor U28482 (N_28482,N_28156,N_28060);
nor U28483 (N_28483,N_27997,N_28055);
nor U28484 (N_28484,N_28173,N_28167);
xor U28485 (N_28485,N_27962,N_27934);
nand U28486 (N_28486,N_28065,N_27922);
nor U28487 (N_28487,N_27992,N_28153);
and U28488 (N_28488,N_28113,N_28018);
xor U28489 (N_28489,N_28171,N_28085);
nor U28490 (N_28490,N_27980,N_27960);
nor U28491 (N_28491,N_28117,N_27916);
nor U28492 (N_28492,N_27933,N_28128);
xnor U28493 (N_28493,N_27917,N_28021);
nor U28494 (N_28494,N_27916,N_28062);
xor U28495 (N_28495,N_28094,N_28161);
or U28496 (N_28496,N_28031,N_28115);
or U28497 (N_28497,N_28084,N_27955);
xnor U28498 (N_28498,N_28134,N_28154);
xor U28499 (N_28499,N_27924,N_27939);
nor U28500 (N_28500,N_28466,N_28426);
and U28501 (N_28501,N_28315,N_28327);
and U28502 (N_28502,N_28260,N_28477);
xnor U28503 (N_28503,N_28333,N_28335);
xnor U28504 (N_28504,N_28236,N_28310);
nor U28505 (N_28505,N_28432,N_28252);
nand U28506 (N_28506,N_28206,N_28225);
nor U28507 (N_28507,N_28301,N_28235);
nand U28508 (N_28508,N_28233,N_28283);
and U28509 (N_28509,N_28438,N_28314);
or U28510 (N_28510,N_28340,N_28448);
nand U28511 (N_28511,N_28378,N_28353);
nand U28512 (N_28512,N_28482,N_28462);
and U28513 (N_28513,N_28433,N_28223);
or U28514 (N_28514,N_28326,N_28384);
nand U28515 (N_28515,N_28291,N_28268);
nor U28516 (N_28516,N_28275,N_28460);
nor U28517 (N_28517,N_28309,N_28272);
nand U28518 (N_28518,N_28342,N_28253);
nor U28519 (N_28519,N_28211,N_28496);
nand U28520 (N_28520,N_28422,N_28456);
and U28521 (N_28521,N_28352,N_28481);
xor U28522 (N_28522,N_28437,N_28490);
and U28523 (N_28523,N_28232,N_28436);
nor U28524 (N_28524,N_28341,N_28351);
or U28525 (N_28525,N_28423,N_28312);
nand U28526 (N_28526,N_28300,N_28402);
xor U28527 (N_28527,N_28304,N_28418);
nor U28528 (N_28528,N_28397,N_28488);
xnor U28529 (N_28529,N_28344,N_28396);
xor U28530 (N_28530,N_28284,N_28205);
nand U28531 (N_28531,N_28201,N_28263);
or U28532 (N_28532,N_28428,N_28487);
nor U28533 (N_28533,N_28354,N_28350);
nor U28534 (N_28534,N_28246,N_28322);
nor U28535 (N_28535,N_28209,N_28323);
or U28536 (N_28536,N_28416,N_28439);
nand U28537 (N_28537,N_28240,N_28227);
nand U28538 (N_28538,N_28474,N_28492);
xnor U28539 (N_28539,N_28243,N_28425);
nand U28540 (N_28540,N_28364,N_28299);
nor U28541 (N_28541,N_28334,N_28228);
xnor U28542 (N_28542,N_28365,N_28415);
nor U28543 (N_28543,N_28319,N_28339);
nand U28544 (N_28544,N_28497,N_28398);
and U28545 (N_28545,N_28403,N_28271);
nand U28546 (N_28546,N_28208,N_28214);
nand U28547 (N_28547,N_28347,N_28287);
and U28548 (N_28548,N_28368,N_28348);
xor U28549 (N_28549,N_28220,N_28358);
xnor U28550 (N_28550,N_28336,N_28254);
nor U28551 (N_28551,N_28213,N_28495);
xnor U28552 (N_28552,N_28306,N_28251);
xnor U28553 (N_28553,N_28421,N_28371);
and U28554 (N_28554,N_28385,N_28391);
nand U28555 (N_28555,N_28210,N_28412);
and U28556 (N_28556,N_28294,N_28404);
or U28557 (N_28557,N_28229,N_28349);
nor U28558 (N_28558,N_28429,N_28467);
nor U28559 (N_28559,N_28461,N_28362);
nand U28560 (N_28560,N_28269,N_28231);
nor U28561 (N_28561,N_28443,N_28386);
xor U28562 (N_28562,N_28454,N_28457);
xor U28563 (N_28563,N_28279,N_28498);
or U28564 (N_28564,N_28472,N_28313);
or U28565 (N_28565,N_28376,N_28224);
xnor U28566 (N_28566,N_28255,N_28302);
nand U28567 (N_28567,N_28463,N_28483);
and U28568 (N_28568,N_28381,N_28395);
and U28569 (N_28569,N_28289,N_28222);
xnor U28570 (N_28570,N_28346,N_28247);
nand U28571 (N_28571,N_28435,N_28297);
nand U28572 (N_28572,N_28379,N_28394);
nor U28573 (N_28573,N_28264,N_28370);
nand U28574 (N_28574,N_28484,N_28331);
and U28575 (N_28575,N_28296,N_28245);
and U28576 (N_28576,N_28455,N_28382);
and U28577 (N_28577,N_28337,N_28430);
nor U28578 (N_28578,N_28413,N_28444);
xnor U28579 (N_28579,N_28308,N_28285);
or U28580 (N_28580,N_28345,N_28311);
nor U28581 (N_28581,N_28372,N_28321);
nor U28582 (N_28582,N_28401,N_28499);
or U28583 (N_28583,N_28475,N_28389);
nand U28584 (N_28584,N_28355,N_28257);
nand U28585 (N_28585,N_28249,N_28357);
and U28586 (N_28586,N_28274,N_28410);
and U28587 (N_28587,N_28479,N_28238);
nand U28588 (N_28588,N_28375,N_28441);
xor U28589 (N_28589,N_28219,N_28281);
nor U28590 (N_28590,N_28261,N_28226);
or U28591 (N_28591,N_28452,N_28248);
and U28592 (N_28592,N_28307,N_28414);
and U28593 (N_28593,N_28465,N_28303);
or U28594 (N_28594,N_28325,N_28278);
and U28595 (N_28595,N_28380,N_28359);
xnor U28596 (N_28596,N_28200,N_28361);
nor U28597 (N_28597,N_28332,N_28434);
xnor U28598 (N_28598,N_28305,N_28320);
nand U28599 (N_28599,N_28318,N_28242);
and U28600 (N_28600,N_28230,N_28393);
nand U28601 (N_28601,N_28471,N_28377);
nor U28602 (N_28602,N_28446,N_28366);
or U28603 (N_28603,N_28316,N_28400);
xor U28604 (N_28604,N_28241,N_28215);
nand U28605 (N_28605,N_28470,N_28343);
and U28606 (N_28606,N_28330,N_28324);
and U28607 (N_28607,N_28203,N_28478);
xnor U28608 (N_28608,N_28445,N_28480);
and U28609 (N_28609,N_28221,N_28383);
nand U28610 (N_28610,N_28292,N_28207);
or U28611 (N_28611,N_28374,N_28329);
and U28612 (N_28612,N_28202,N_28392);
nor U28613 (N_28613,N_28237,N_28280);
nor U28614 (N_28614,N_28388,N_28411);
nand U28615 (N_28615,N_28258,N_28420);
nand U28616 (N_28616,N_28464,N_28390);
nand U28617 (N_28617,N_28204,N_28486);
nand U28618 (N_28618,N_28266,N_28458);
or U28619 (N_28619,N_28494,N_28459);
or U28620 (N_28620,N_28276,N_28367);
nor U28621 (N_28621,N_28338,N_28363);
or U28622 (N_28622,N_28239,N_28409);
xnor U28623 (N_28623,N_28405,N_28369);
and U28624 (N_28624,N_28449,N_28493);
xnor U28625 (N_28625,N_28267,N_28262);
xnor U28626 (N_28626,N_28298,N_28408);
xnor U28627 (N_28627,N_28451,N_28427);
nand U28628 (N_28628,N_28256,N_28442);
xnor U28629 (N_28629,N_28212,N_28476);
nand U28630 (N_28630,N_28440,N_28360);
and U28631 (N_28631,N_28469,N_28216);
nor U28632 (N_28632,N_28419,N_28295);
or U28633 (N_28633,N_28288,N_28282);
or U28634 (N_28634,N_28234,N_28489);
or U28635 (N_28635,N_28265,N_28290);
xnor U28636 (N_28636,N_28485,N_28406);
xor U28637 (N_28637,N_28431,N_28447);
nor U28638 (N_28638,N_28356,N_28317);
and U28639 (N_28639,N_28468,N_28277);
nor U28640 (N_28640,N_28399,N_28259);
nor U28641 (N_28641,N_28491,N_28250);
nand U28642 (N_28642,N_28387,N_28270);
or U28643 (N_28643,N_28373,N_28407);
nor U28644 (N_28644,N_28273,N_28293);
nor U28645 (N_28645,N_28244,N_28424);
nand U28646 (N_28646,N_28286,N_28450);
and U28647 (N_28647,N_28453,N_28217);
or U28648 (N_28648,N_28328,N_28473);
or U28649 (N_28649,N_28218,N_28417);
and U28650 (N_28650,N_28283,N_28296);
or U28651 (N_28651,N_28259,N_28354);
or U28652 (N_28652,N_28307,N_28421);
nand U28653 (N_28653,N_28474,N_28359);
nand U28654 (N_28654,N_28352,N_28489);
nand U28655 (N_28655,N_28222,N_28260);
and U28656 (N_28656,N_28231,N_28347);
xnor U28657 (N_28657,N_28423,N_28341);
and U28658 (N_28658,N_28459,N_28292);
or U28659 (N_28659,N_28270,N_28295);
and U28660 (N_28660,N_28447,N_28485);
and U28661 (N_28661,N_28450,N_28477);
nor U28662 (N_28662,N_28276,N_28451);
or U28663 (N_28663,N_28466,N_28423);
nand U28664 (N_28664,N_28465,N_28373);
xnor U28665 (N_28665,N_28333,N_28247);
xor U28666 (N_28666,N_28266,N_28219);
nor U28667 (N_28667,N_28238,N_28385);
and U28668 (N_28668,N_28371,N_28229);
and U28669 (N_28669,N_28251,N_28350);
nand U28670 (N_28670,N_28231,N_28391);
and U28671 (N_28671,N_28472,N_28438);
or U28672 (N_28672,N_28234,N_28276);
nand U28673 (N_28673,N_28421,N_28381);
nand U28674 (N_28674,N_28349,N_28468);
nor U28675 (N_28675,N_28259,N_28429);
and U28676 (N_28676,N_28210,N_28431);
nand U28677 (N_28677,N_28246,N_28357);
xnor U28678 (N_28678,N_28352,N_28201);
xnor U28679 (N_28679,N_28464,N_28415);
xnor U28680 (N_28680,N_28395,N_28207);
xor U28681 (N_28681,N_28372,N_28475);
nand U28682 (N_28682,N_28303,N_28263);
or U28683 (N_28683,N_28369,N_28201);
nand U28684 (N_28684,N_28345,N_28278);
or U28685 (N_28685,N_28338,N_28256);
nor U28686 (N_28686,N_28352,N_28454);
nor U28687 (N_28687,N_28461,N_28206);
and U28688 (N_28688,N_28410,N_28235);
nor U28689 (N_28689,N_28254,N_28342);
or U28690 (N_28690,N_28207,N_28490);
xor U28691 (N_28691,N_28303,N_28299);
and U28692 (N_28692,N_28289,N_28447);
nand U28693 (N_28693,N_28430,N_28448);
nand U28694 (N_28694,N_28299,N_28411);
xnor U28695 (N_28695,N_28293,N_28356);
or U28696 (N_28696,N_28473,N_28438);
nand U28697 (N_28697,N_28276,N_28294);
or U28698 (N_28698,N_28480,N_28336);
and U28699 (N_28699,N_28432,N_28462);
nor U28700 (N_28700,N_28212,N_28370);
and U28701 (N_28701,N_28453,N_28406);
nand U28702 (N_28702,N_28461,N_28279);
nor U28703 (N_28703,N_28348,N_28319);
nor U28704 (N_28704,N_28415,N_28498);
nand U28705 (N_28705,N_28434,N_28264);
nand U28706 (N_28706,N_28326,N_28471);
nor U28707 (N_28707,N_28278,N_28330);
nand U28708 (N_28708,N_28496,N_28284);
nor U28709 (N_28709,N_28474,N_28230);
and U28710 (N_28710,N_28300,N_28384);
nor U28711 (N_28711,N_28422,N_28386);
xor U28712 (N_28712,N_28470,N_28204);
xor U28713 (N_28713,N_28331,N_28434);
and U28714 (N_28714,N_28212,N_28407);
nand U28715 (N_28715,N_28446,N_28483);
xor U28716 (N_28716,N_28260,N_28241);
nand U28717 (N_28717,N_28224,N_28317);
nand U28718 (N_28718,N_28205,N_28351);
or U28719 (N_28719,N_28349,N_28447);
xnor U28720 (N_28720,N_28253,N_28415);
nor U28721 (N_28721,N_28224,N_28307);
xnor U28722 (N_28722,N_28340,N_28400);
xor U28723 (N_28723,N_28327,N_28434);
nand U28724 (N_28724,N_28200,N_28490);
and U28725 (N_28725,N_28312,N_28402);
xor U28726 (N_28726,N_28434,N_28413);
nand U28727 (N_28727,N_28326,N_28306);
or U28728 (N_28728,N_28441,N_28207);
or U28729 (N_28729,N_28330,N_28251);
and U28730 (N_28730,N_28300,N_28455);
or U28731 (N_28731,N_28271,N_28362);
and U28732 (N_28732,N_28315,N_28407);
nor U28733 (N_28733,N_28385,N_28227);
or U28734 (N_28734,N_28207,N_28332);
or U28735 (N_28735,N_28350,N_28311);
xnor U28736 (N_28736,N_28206,N_28349);
and U28737 (N_28737,N_28355,N_28350);
and U28738 (N_28738,N_28308,N_28250);
xnor U28739 (N_28739,N_28343,N_28440);
and U28740 (N_28740,N_28232,N_28300);
and U28741 (N_28741,N_28293,N_28452);
or U28742 (N_28742,N_28470,N_28451);
or U28743 (N_28743,N_28442,N_28254);
nand U28744 (N_28744,N_28494,N_28241);
or U28745 (N_28745,N_28447,N_28293);
or U28746 (N_28746,N_28298,N_28271);
xor U28747 (N_28747,N_28234,N_28222);
and U28748 (N_28748,N_28279,N_28360);
nor U28749 (N_28749,N_28390,N_28470);
or U28750 (N_28750,N_28328,N_28275);
and U28751 (N_28751,N_28419,N_28336);
nor U28752 (N_28752,N_28249,N_28356);
and U28753 (N_28753,N_28392,N_28276);
nor U28754 (N_28754,N_28315,N_28458);
nand U28755 (N_28755,N_28447,N_28328);
nand U28756 (N_28756,N_28212,N_28293);
xnor U28757 (N_28757,N_28457,N_28467);
and U28758 (N_28758,N_28486,N_28303);
or U28759 (N_28759,N_28405,N_28370);
or U28760 (N_28760,N_28470,N_28278);
nand U28761 (N_28761,N_28410,N_28446);
and U28762 (N_28762,N_28434,N_28382);
and U28763 (N_28763,N_28481,N_28322);
or U28764 (N_28764,N_28447,N_28207);
or U28765 (N_28765,N_28434,N_28401);
nor U28766 (N_28766,N_28481,N_28488);
nand U28767 (N_28767,N_28387,N_28414);
nand U28768 (N_28768,N_28225,N_28330);
xor U28769 (N_28769,N_28383,N_28358);
nor U28770 (N_28770,N_28255,N_28409);
xor U28771 (N_28771,N_28385,N_28321);
or U28772 (N_28772,N_28419,N_28434);
or U28773 (N_28773,N_28210,N_28421);
xor U28774 (N_28774,N_28320,N_28333);
xor U28775 (N_28775,N_28261,N_28472);
nand U28776 (N_28776,N_28212,N_28259);
xor U28777 (N_28777,N_28436,N_28308);
nor U28778 (N_28778,N_28295,N_28237);
xor U28779 (N_28779,N_28361,N_28496);
xnor U28780 (N_28780,N_28460,N_28348);
nor U28781 (N_28781,N_28216,N_28259);
and U28782 (N_28782,N_28495,N_28405);
nor U28783 (N_28783,N_28400,N_28289);
nand U28784 (N_28784,N_28351,N_28406);
or U28785 (N_28785,N_28268,N_28279);
nand U28786 (N_28786,N_28414,N_28489);
and U28787 (N_28787,N_28325,N_28202);
or U28788 (N_28788,N_28228,N_28274);
nand U28789 (N_28789,N_28253,N_28354);
or U28790 (N_28790,N_28303,N_28396);
and U28791 (N_28791,N_28358,N_28282);
nor U28792 (N_28792,N_28297,N_28267);
nor U28793 (N_28793,N_28392,N_28324);
nor U28794 (N_28794,N_28347,N_28324);
and U28795 (N_28795,N_28499,N_28399);
and U28796 (N_28796,N_28365,N_28283);
xnor U28797 (N_28797,N_28273,N_28254);
xor U28798 (N_28798,N_28495,N_28481);
nor U28799 (N_28799,N_28404,N_28280);
nand U28800 (N_28800,N_28556,N_28626);
nor U28801 (N_28801,N_28663,N_28680);
xnor U28802 (N_28802,N_28686,N_28796);
nor U28803 (N_28803,N_28532,N_28718);
xnor U28804 (N_28804,N_28531,N_28620);
nor U28805 (N_28805,N_28522,N_28535);
nand U28806 (N_28806,N_28662,N_28669);
nand U28807 (N_28807,N_28752,N_28761);
nand U28808 (N_28808,N_28629,N_28731);
nand U28809 (N_28809,N_28638,N_28739);
and U28810 (N_28810,N_28505,N_28746);
nand U28811 (N_28811,N_28719,N_28735);
or U28812 (N_28812,N_28644,N_28655);
xnor U28813 (N_28813,N_28722,N_28727);
xnor U28814 (N_28814,N_28592,N_28706);
or U28815 (N_28815,N_28519,N_28747);
xor U28816 (N_28816,N_28695,N_28616);
nor U28817 (N_28817,N_28676,N_28681);
nand U28818 (N_28818,N_28593,N_28760);
and U28819 (N_28819,N_28691,N_28788);
nand U28820 (N_28820,N_28774,N_28643);
nor U28821 (N_28821,N_28512,N_28555);
and U28822 (N_28822,N_28503,N_28653);
and U28823 (N_28823,N_28603,N_28530);
nor U28824 (N_28824,N_28633,N_28732);
nor U28825 (N_28825,N_28553,N_28594);
nor U28826 (N_28826,N_28674,N_28725);
and U28827 (N_28827,N_28795,N_28610);
nand U28828 (N_28828,N_28640,N_28697);
and U28829 (N_28829,N_28611,N_28584);
xnor U28830 (N_28830,N_28587,N_28736);
and U28831 (N_28831,N_28692,N_28576);
or U28832 (N_28832,N_28600,N_28518);
nand U28833 (N_28833,N_28789,N_28609);
and U28834 (N_28834,N_28661,N_28766);
nor U28835 (N_28835,N_28758,N_28744);
and U28836 (N_28836,N_28711,N_28548);
xor U28837 (N_28837,N_28776,N_28597);
nand U28838 (N_28838,N_28544,N_28536);
xor U28839 (N_28839,N_28724,N_28621);
and U28840 (N_28840,N_28690,N_28707);
xor U28841 (N_28841,N_28688,N_28702);
or U28842 (N_28842,N_28666,N_28667);
nor U28843 (N_28843,N_28525,N_28660);
xor U28844 (N_28844,N_28684,N_28772);
and U28845 (N_28845,N_28743,N_28648);
and U28846 (N_28846,N_28786,N_28582);
or U28847 (N_28847,N_28765,N_28751);
xnor U28848 (N_28848,N_28793,N_28524);
or U28849 (N_28849,N_28658,N_28750);
xnor U28850 (N_28850,N_28665,N_28779);
nor U28851 (N_28851,N_28654,N_28650);
nor U28852 (N_28852,N_28710,N_28708);
nor U28853 (N_28853,N_28717,N_28683);
nor U28854 (N_28854,N_28664,N_28798);
or U28855 (N_28855,N_28539,N_28685);
xnor U28856 (N_28856,N_28678,N_28615);
nand U28857 (N_28857,N_28714,N_28755);
or U28858 (N_28858,N_28728,N_28769);
nor U28859 (N_28859,N_28740,N_28699);
xor U28860 (N_28860,N_28618,N_28780);
nor U28861 (N_28861,N_28602,N_28627);
and U28862 (N_28862,N_28726,N_28687);
xnor U28863 (N_28863,N_28575,N_28723);
xor U28864 (N_28864,N_28785,N_28570);
or U28865 (N_28865,N_28645,N_28546);
and U28866 (N_28866,N_28799,N_28513);
nor U28867 (N_28867,N_28639,N_28588);
nand U28868 (N_28868,N_28730,N_28696);
and U28869 (N_28869,N_28567,N_28698);
or U28870 (N_28870,N_28533,N_28565);
nand U28871 (N_28871,N_28578,N_28738);
nor U28872 (N_28872,N_28500,N_28560);
xor U28873 (N_28873,N_28734,N_28541);
or U28874 (N_28874,N_28506,N_28689);
or U28875 (N_28875,N_28651,N_28540);
nor U28876 (N_28876,N_28713,N_28599);
xor U28877 (N_28877,N_28613,N_28514);
and U28878 (N_28878,N_28516,N_28771);
nand U28879 (N_28879,N_28564,N_28538);
nor U28880 (N_28880,N_28794,N_28583);
or U28881 (N_28881,N_28557,N_28569);
or U28882 (N_28882,N_28781,N_28608);
or U28883 (N_28883,N_28579,N_28580);
xor U28884 (N_28884,N_28716,N_28501);
nor U28885 (N_28885,N_28652,N_28762);
xnor U28886 (N_28886,N_28756,N_28659);
nor U28887 (N_28887,N_28612,N_28574);
or U28888 (N_28888,N_28768,N_28549);
xnor U28889 (N_28889,N_28764,N_28721);
xor U28890 (N_28890,N_28649,N_28502);
xnor U28891 (N_28891,N_28797,N_28631);
and U28892 (N_28892,N_28509,N_28563);
and U28893 (N_28893,N_28550,N_28586);
nor U28894 (N_28894,N_28517,N_28700);
nand U28895 (N_28895,N_28508,N_28606);
nor U28896 (N_28896,N_28623,N_28720);
nor U28897 (N_28897,N_28705,N_28537);
nor U28898 (N_28898,N_28520,N_28529);
and U28899 (N_28899,N_28635,N_28694);
and U28900 (N_28900,N_28775,N_28715);
nand U28901 (N_28901,N_28693,N_28634);
or U28902 (N_28902,N_28784,N_28677);
and U28903 (N_28903,N_28742,N_28757);
xor U28904 (N_28904,N_28543,N_28767);
nand U28905 (N_28905,N_28754,N_28581);
xnor U28906 (N_28906,N_28624,N_28590);
nand U28907 (N_28907,N_28679,N_28577);
nor U28908 (N_28908,N_28542,N_28632);
and U28909 (N_28909,N_28783,N_28507);
nor U28910 (N_28910,N_28657,N_28559);
and U28911 (N_28911,N_28607,N_28511);
and U28912 (N_28912,N_28791,N_28673);
and U28913 (N_28913,N_28668,N_28670);
and U28914 (N_28914,N_28605,N_28562);
xnor U28915 (N_28915,N_28656,N_28534);
nand U28916 (N_28916,N_28753,N_28545);
or U28917 (N_28917,N_28598,N_28561);
nor U28918 (N_28918,N_28790,N_28571);
and U28919 (N_28919,N_28749,N_28778);
nand U28920 (N_28920,N_28617,N_28777);
nand U28921 (N_28921,N_28646,N_28625);
and U28922 (N_28922,N_28733,N_28591);
nor U28923 (N_28923,N_28709,N_28782);
and U28924 (N_28924,N_28601,N_28787);
xor U28925 (N_28925,N_28675,N_28748);
nor U28926 (N_28926,N_28745,N_28573);
nand U28927 (N_28927,N_28630,N_28712);
nor U28928 (N_28928,N_28595,N_28528);
or U28929 (N_28929,N_28510,N_28763);
and U28930 (N_28930,N_28547,N_28642);
or U28931 (N_28931,N_28554,N_28589);
and U28932 (N_28932,N_28729,N_28704);
nand U28933 (N_28933,N_28770,N_28641);
nand U28934 (N_28934,N_28604,N_28527);
nand U28935 (N_28935,N_28566,N_28622);
nand U28936 (N_28936,N_28628,N_28682);
or U28937 (N_28937,N_28596,N_28572);
xor U28938 (N_28938,N_28647,N_28741);
or U28939 (N_28939,N_28552,N_28585);
nor U28940 (N_28940,N_28672,N_28636);
and U28941 (N_28941,N_28737,N_28701);
and U28942 (N_28942,N_28792,N_28504);
nand U28943 (N_28943,N_28521,N_28515);
xnor U28944 (N_28944,N_28568,N_28558);
nor U28945 (N_28945,N_28614,N_28703);
nand U28946 (N_28946,N_28551,N_28526);
and U28947 (N_28947,N_28759,N_28619);
nand U28948 (N_28948,N_28773,N_28637);
or U28949 (N_28949,N_28523,N_28671);
xor U28950 (N_28950,N_28574,N_28731);
nand U28951 (N_28951,N_28770,N_28534);
nor U28952 (N_28952,N_28712,N_28695);
nand U28953 (N_28953,N_28641,N_28562);
or U28954 (N_28954,N_28519,N_28772);
and U28955 (N_28955,N_28652,N_28615);
and U28956 (N_28956,N_28577,N_28511);
nand U28957 (N_28957,N_28739,N_28650);
xor U28958 (N_28958,N_28762,N_28595);
nand U28959 (N_28959,N_28745,N_28542);
nand U28960 (N_28960,N_28769,N_28612);
nand U28961 (N_28961,N_28559,N_28537);
and U28962 (N_28962,N_28652,N_28609);
nand U28963 (N_28963,N_28527,N_28759);
and U28964 (N_28964,N_28774,N_28740);
nor U28965 (N_28965,N_28697,N_28574);
or U28966 (N_28966,N_28721,N_28625);
or U28967 (N_28967,N_28681,N_28758);
nand U28968 (N_28968,N_28687,N_28698);
nand U28969 (N_28969,N_28731,N_28730);
or U28970 (N_28970,N_28623,N_28552);
or U28971 (N_28971,N_28616,N_28539);
nand U28972 (N_28972,N_28722,N_28723);
nand U28973 (N_28973,N_28574,N_28666);
xnor U28974 (N_28974,N_28721,N_28716);
and U28975 (N_28975,N_28752,N_28555);
or U28976 (N_28976,N_28572,N_28789);
xor U28977 (N_28977,N_28775,N_28777);
nand U28978 (N_28978,N_28572,N_28546);
xor U28979 (N_28979,N_28700,N_28759);
or U28980 (N_28980,N_28660,N_28553);
xnor U28981 (N_28981,N_28524,N_28530);
and U28982 (N_28982,N_28663,N_28736);
nand U28983 (N_28983,N_28713,N_28743);
nor U28984 (N_28984,N_28778,N_28651);
nand U28985 (N_28985,N_28732,N_28651);
and U28986 (N_28986,N_28676,N_28501);
nor U28987 (N_28987,N_28753,N_28593);
nand U28988 (N_28988,N_28662,N_28646);
or U28989 (N_28989,N_28765,N_28643);
xnor U28990 (N_28990,N_28524,N_28659);
nor U28991 (N_28991,N_28788,N_28714);
and U28992 (N_28992,N_28705,N_28781);
or U28993 (N_28993,N_28516,N_28562);
or U28994 (N_28994,N_28638,N_28756);
nor U28995 (N_28995,N_28616,N_28697);
and U28996 (N_28996,N_28766,N_28550);
nor U28997 (N_28997,N_28697,N_28683);
nor U28998 (N_28998,N_28717,N_28703);
nand U28999 (N_28999,N_28782,N_28547);
xnor U29000 (N_29000,N_28699,N_28791);
or U29001 (N_29001,N_28504,N_28588);
and U29002 (N_29002,N_28736,N_28784);
nand U29003 (N_29003,N_28563,N_28624);
or U29004 (N_29004,N_28634,N_28616);
nand U29005 (N_29005,N_28601,N_28501);
and U29006 (N_29006,N_28722,N_28744);
nand U29007 (N_29007,N_28650,N_28543);
xor U29008 (N_29008,N_28676,N_28554);
xor U29009 (N_29009,N_28513,N_28510);
xor U29010 (N_29010,N_28645,N_28658);
xnor U29011 (N_29011,N_28684,N_28606);
and U29012 (N_29012,N_28763,N_28545);
xnor U29013 (N_29013,N_28750,N_28771);
and U29014 (N_29014,N_28579,N_28510);
or U29015 (N_29015,N_28591,N_28667);
xor U29016 (N_29016,N_28657,N_28525);
xnor U29017 (N_29017,N_28609,N_28558);
nand U29018 (N_29018,N_28539,N_28569);
xnor U29019 (N_29019,N_28768,N_28789);
nor U29020 (N_29020,N_28702,N_28526);
and U29021 (N_29021,N_28667,N_28548);
and U29022 (N_29022,N_28784,N_28778);
nor U29023 (N_29023,N_28655,N_28791);
or U29024 (N_29024,N_28537,N_28601);
nand U29025 (N_29025,N_28752,N_28523);
xor U29026 (N_29026,N_28721,N_28572);
nor U29027 (N_29027,N_28656,N_28681);
nor U29028 (N_29028,N_28548,N_28590);
nand U29029 (N_29029,N_28598,N_28514);
xor U29030 (N_29030,N_28594,N_28781);
and U29031 (N_29031,N_28647,N_28679);
or U29032 (N_29032,N_28740,N_28688);
nand U29033 (N_29033,N_28507,N_28598);
xor U29034 (N_29034,N_28503,N_28589);
nor U29035 (N_29035,N_28738,N_28575);
nor U29036 (N_29036,N_28799,N_28732);
xnor U29037 (N_29037,N_28518,N_28690);
xor U29038 (N_29038,N_28577,N_28509);
nor U29039 (N_29039,N_28529,N_28516);
nor U29040 (N_29040,N_28600,N_28589);
or U29041 (N_29041,N_28757,N_28513);
nand U29042 (N_29042,N_28775,N_28792);
nand U29043 (N_29043,N_28592,N_28757);
and U29044 (N_29044,N_28537,N_28598);
or U29045 (N_29045,N_28779,N_28721);
xor U29046 (N_29046,N_28739,N_28675);
or U29047 (N_29047,N_28519,N_28724);
or U29048 (N_29048,N_28648,N_28557);
or U29049 (N_29049,N_28604,N_28665);
nand U29050 (N_29050,N_28587,N_28744);
or U29051 (N_29051,N_28655,N_28720);
nand U29052 (N_29052,N_28737,N_28775);
nand U29053 (N_29053,N_28740,N_28516);
and U29054 (N_29054,N_28617,N_28512);
or U29055 (N_29055,N_28786,N_28665);
nand U29056 (N_29056,N_28608,N_28631);
nor U29057 (N_29057,N_28646,N_28740);
xor U29058 (N_29058,N_28778,N_28742);
or U29059 (N_29059,N_28602,N_28547);
xnor U29060 (N_29060,N_28678,N_28744);
nor U29061 (N_29061,N_28600,N_28712);
and U29062 (N_29062,N_28639,N_28567);
xor U29063 (N_29063,N_28542,N_28618);
or U29064 (N_29064,N_28713,N_28546);
nand U29065 (N_29065,N_28693,N_28506);
or U29066 (N_29066,N_28773,N_28743);
nand U29067 (N_29067,N_28636,N_28688);
and U29068 (N_29068,N_28669,N_28541);
or U29069 (N_29069,N_28736,N_28578);
and U29070 (N_29070,N_28760,N_28704);
and U29071 (N_29071,N_28710,N_28692);
and U29072 (N_29072,N_28568,N_28680);
and U29073 (N_29073,N_28653,N_28536);
nor U29074 (N_29074,N_28629,N_28557);
nor U29075 (N_29075,N_28688,N_28551);
nand U29076 (N_29076,N_28790,N_28618);
xor U29077 (N_29077,N_28681,N_28555);
nand U29078 (N_29078,N_28694,N_28753);
or U29079 (N_29079,N_28595,N_28679);
or U29080 (N_29080,N_28686,N_28565);
nand U29081 (N_29081,N_28702,N_28661);
xor U29082 (N_29082,N_28735,N_28617);
and U29083 (N_29083,N_28680,N_28616);
nor U29084 (N_29084,N_28749,N_28605);
or U29085 (N_29085,N_28754,N_28543);
or U29086 (N_29086,N_28773,N_28509);
nor U29087 (N_29087,N_28782,N_28741);
xnor U29088 (N_29088,N_28666,N_28604);
xnor U29089 (N_29089,N_28648,N_28585);
nand U29090 (N_29090,N_28586,N_28574);
and U29091 (N_29091,N_28704,N_28685);
nand U29092 (N_29092,N_28628,N_28674);
or U29093 (N_29093,N_28751,N_28692);
and U29094 (N_29094,N_28681,N_28662);
and U29095 (N_29095,N_28738,N_28632);
xnor U29096 (N_29096,N_28523,N_28783);
and U29097 (N_29097,N_28525,N_28769);
nor U29098 (N_29098,N_28577,N_28740);
nand U29099 (N_29099,N_28782,N_28723);
and U29100 (N_29100,N_29018,N_28996);
nor U29101 (N_29101,N_29041,N_29000);
nand U29102 (N_29102,N_28958,N_28927);
or U29103 (N_29103,N_29017,N_28872);
nand U29104 (N_29104,N_28881,N_29039);
nand U29105 (N_29105,N_28863,N_28959);
and U29106 (N_29106,N_28875,N_29050);
nor U29107 (N_29107,N_29015,N_28809);
nor U29108 (N_29108,N_28906,N_29055);
xor U29109 (N_29109,N_29023,N_28861);
nand U29110 (N_29110,N_29026,N_28912);
xor U29111 (N_29111,N_29074,N_29020);
and U29112 (N_29112,N_28911,N_28807);
xnor U29113 (N_29113,N_29064,N_29006);
nor U29114 (N_29114,N_28888,N_28883);
or U29115 (N_29115,N_28843,N_29066);
or U29116 (N_29116,N_28823,N_28926);
or U29117 (N_29117,N_28878,N_29051);
nor U29118 (N_29118,N_28924,N_28934);
or U29119 (N_29119,N_29057,N_29071);
and U29120 (N_29120,N_29032,N_28837);
nor U29121 (N_29121,N_28916,N_29084);
nand U29122 (N_29122,N_29007,N_29036);
and U29123 (N_29123,N_28860,N_28938);
nor U29124 (N_29124,N_29009,N_28824);
or U29125 (N_29125,N_28955,N_28902);
and U29126 (N_29126,N_28848,N_28873);
or U29127 (N_29127,N_29087,N_28856);
and U29128 (N_29128,N_28967,N_29003);
xnor U29129 (N_29129,N_28846,N_28830);
nor U29130 (N_29130,N_29070,N_28877);
or U29131 (N_29131,N_29053,N_28909);
xnor U29132 (N_29132,N_29092,N_28854);
or U29133 (N_29133,N_28914,N_28960);
nand U29134 (N_29134,N_29011,N_28948);
xnor U29135 (N_29135,N_28835,N_28812);
and U29136 (N_29136,N_29061,N_29079);
xor U29137 (N_29137,N_28841,N_28983);
xor U29138 (N_29138,N_28920,N_28966);
or U29139 (N_29139,N_28870,N_29088);
xnor U29140 (N_29140,N_28853,N_29042);
and U29141 (N_29141,N_28820,N_29052);
and U29142 (N_29142,N_28842,N_29027);
or U29143 (N_29143,N_28831,N_29096);
xnor U29144 (N_29144,N_28851,N_28867);
nor U29145 (N_29145,N_28918,N_28845);
and U29146 (N_29146,N_28847,N_29002);
and U29147 (N_29147,N_29033,N_28836);
nand U29148 (N_29148,N_28986,N_29037);
nand U29149 (N_29149,N_29025,N_29090);
and U29150 (N_29150,N_28972,N_29086);
and U29151 (N_29151,N_29010,N_28969);
nor U29152 (N_29152,N_28975,N_28995);
or U29153 (N_29153,N_28976,N_28989);
nor U29154 (N_29154,N_29004,N_28892);
nor U29155 (N_29155,N_29067,N_28801);
or U29156 (N_29156,N_28947,N_28868);
or U29157 (N_29157,N_28990,N_29091);
and U29158 (N_29158,N_28803,N_28827);
xor U29159 (N_29159,N_29034,N_29062);
xor U29160 (N_29160,N_29093,N_28855);
or U29161 (N_29161,N_28805,N_28915);
xor U29162 (N_29162,N_28961,N_28997);
and U29163 (N_29163,N_28862,N_29013);
nor U29164 (N_29164,N_29058,N_29063);
xor U29165 (N_29165,N_28815,N_28840);
or U29166 (N_29166,N_28818,N_28814);
nand U29167 (N_29167,N_28932,N_28882);
xor U29168 (N_29168,N_29045,N_28890);
or U29169 (N_29169,N_28925,N_28931);
nor U29170 (N_29170,N_28802,N_28844);
or U29171 (N_29171,N_28944,N_28866);
nor U29172 (N_29172,N_29097,N_29035);
nand U29173 (N_29173,N_28808,N_29077);
or U29174 (N_29174,N_28923,N_28834);
nand U29175 (N_29175,N_28813,N_29095);
or U29176 (N_29176,N_28833,N_28933);
nor U29177 (N_29177,N_28919,N_29082);
nor U29178 (N_29178,N_28858,N_28945);
or U29179 (N_29179,N_28968,N_28810);
or U29180 (N_29180,N_29016,N_28826);
and U29181 (N_29181,N_28994,N_29073);
nand U29182 (N_29182,N_28998,N_28921);
nor U29183 (N_29183,N_28825,N_28942);
xnor U29184 (N_29184,N_28937,N_29075);
xnor U29185 (N_29185,N_29040,N_28965);
nand U29186 (N_29186,N_28889,N_29048);
or U29187 (N_29187,N_29081,N_28832);
and U29188 (N_29188,N_29046,N_28839);
nor U29189 (N_29189,N_29054,N_28884);
and U29190 (N_29190,N_29043,N_28903);
or U29191 (N_29191,N_29012,N_28964);
nand U29192 (N_29192,N_28829,N_28979);
nor U29193 (N_29193,N_28849,N_28816);
nor U29194 (N_29194,N_29069,N_28900);
or U29195 (N_29195,N_28895,N_28864);
nor U29196 (N_29196,N_28984,N_29028);
nand U29197 (N_29197,N_28800,N_28822);
nor U29198 (N_29198,N_29014,N_29021);
xnor U29199 (N_29199,N_28904,N_28897);
and U29200 (N_29200,N_29068,N_29065);
nor U29201 (N_29201,N_28974,N_28930);
nor U29202 (N_29202,N_28894,N_29029);
xor U29203 (N_29203,N_28950,N_28946);
and U29204 (N_29204,N_28896,N_28988);
or U29205 (N_29205,N_28804,N_28879);
nand U29206 (N_29206,N_29019,N_28908);
and U29207 (N_29207,N_28939,N_29022);
nor U29208 (N_29208,N_28876,N_28865);
xnor U29209 (N_29209,N_29005,N_28999);
nand U29210 (N_29210,N_28907,N_28817);
xor U29211 (N_29211,N_28949,N_28905);
nand U29212 (N_29212,N_28913,N_28940);
nand U29213 (N_29213,N_28898,N_28891);
and U29214 (N_29214,N_29024,N_29056);
xnor U29215 (N_29215,N_29001,N_28970);
or U29216 (N_29216,N_28985,N_28929);
nand U29217 (N_29217,N_28982,N_28887);
nand U29218 (N_29218,N_29030,N_28901);
or U29219 (N_29219,N_29049,N_28941);
nor U29220 (N_29220,N_28981,N_28917);
or U29221 (N_29221,N_28819,N_28859);
nand U29222 (N_29222,N_28936,N_28828);
xor U29223 (N_29223,N_28992,N_28971);
and U29224 (N_29224,N_28957,N_28821);
xnor U29225 (N_29225,N_28977,N_28811);
nand U29226 (N_29226,N_28993,N_28953);
and U29227 (N_29227,N_28899,N_28838);
xnor U29228 (N_29228,N_28922,N_29047);
nand U29229 (N_29229,N_28951,N_28869);
and U29230 (N_29230,N_28991,N_29098);
nor U29231 (N_29231,N_28963,N_28850);
or U29232 (N_29232,N_29072,N_29038);
nand U29233 (N_29233,N_28852,N_29099);
or U29234 (N_29234,N_29059,N_28956);
nand U29235 (N_29235,N_29078,N_29008);
xnor U29236 (N_29236,N_28857,N_28987);
xor U29237 (N_29237,N_29060,N_28910);
or U29238 (N_29238,N_29089,N_28886);
xor U29239 (N_29239,N_29094,N_29083);
and U29240 (N_29240,N_28978,N_28806);
and U29241 (N_29241,N_28943,N_28928);
nand U29242 (N_29242,N_28973,N_28935);
and U29243 (N_29243,N_29080,N_28880);
and U29244 (N_29244,N_29076,N_29031);
and U29245 (N_29245,N_28952,N_28871);
nor U29246 (N_29246,N_28980,N_28962);
nand U29247 (N_29247,N_28885,N_29044);
xor U29248 (N_29248,N_28954,N_28874);
xnor U29249 (N_29249,N_29085,N_28893);
xor U29250 (N_29250,N_28843,N_29000);
xor U29251 (N_29251,N_28972,N_28834);
nand U29252 (N_29252,N_28816,N_28986);
or U29253 (N_29253,N_28906,N_28883);
nor U29254 (N_29254,N_28832,N_28844);
and U29255 (N_29255,N_29042,N_29041);
xor U29256 (N_29256,N_28987,N_28971);
nand U29257 (N_29257,N_28844,N_28927);
nor U29258 (N_29258,N_28866,N_29035);
nand U29259 (N_29259,N_29096,N_28945);
or U29260 (N_29260,N_29070,N_28840);
xor U29261 (N_29261,N_28854,N_28978);
nor U29262 (N_29262,N_28869,N_29054);
xor U29263 (N_29263,N_29002,N_28965);
and U29264 (N_29264,N_28946,N_29068);
and U29265 (N_29265,N_28868,N_28873);
nor U29266 (N_29266,N_29038,N_28847);
or U29267 (N_29267,N_28848,N_28923);
xor U29268 (N_29268,N_28927,N_29095);
xnor U29269 (N_29269,N_28895,N_28973);
or U29270 (N_29270,N_28859,N_29073);
and U29271 (N_29271,N_28982,N_29099);
nor U29272 (N_29272,N_28934,N_28855);
or U29273 (N_29273,N_28898,N_29071);
nand U29274 (N_29274,N_28908,N_29013);
and U29275 (N_29275,N_28856,N_28804);
or U29276 (N_29276,N_28951,N_29065);
or U29277 (N_29277,N_29098,N_29074);
nor U29278 (N_29278,N_29025,N_28991);
or U29279 (N_29279,N_29037,N_28947);
nand U29280 (N_29280,N_28961,N_28844);
or U29281 (N_29281,N_28900,N_29098);
or U29282 (N_29282,N_29083,N_28974);
nand U29283 (N_29283,N_28984,N_28833);
nor U29284 (N_29284,N_28950,N_29003);
nor U29285 (N_29285,N_28876,N_28980);
nand U29286 (N_29286,N_28820,N_29099);
or U29287 (N_29287,N_28954,N_29037);
xnor U29288 (N_29288,N_28876,N_29077);
nand U29289 (N_29289,N_28951,N_28847);
xnor U29290 (N_29290,N_29013,N_28830);
xor U29291 (N_29291,N_29065,N_29097);
xor U29292 (N_29292,N_29077,N_28891);
nor U29293 (N_29293,N_28837,N_28817);
and U29294 (N_29294,N_28987,N_29054);
and U29295 (N_29295,N_28866,N_28978);
xor U29296 (N_29296,N_28906,N_28951);
nor U29297 (N_29297,N_28893,N_29089);
xnor U29298 (N_29298,N_29018,N_28993);
or U29299 (N_29299,N_28806,N_29019);
nand U29300 (N_29300,N_29025,N_28908);
xnor U29301 (N_29301,N_28864,N_28885);
xnor U29302 (N_29302,N_28820,N_29054);
xnor U29303 (N_29303,N_28919,N_28857);
nand U29304 (N_29304,N_28917,N_29027);
and U29305 (N_29305,N_28965,N_29015);
or U29306 (N_29306,N_29028,N_28822);
xnor U29307 (N_29307,N_29010,N_28894);
or U29308 (N_29308,N_28929,N_28890);
xor U29309 (N_29309,N_28891,N_28841);
or U29310 (N_29310,N_28801,N_28876);
and U29311 (N_29311,N_28884,N_28864);
xnor U29312 (N_29312,N_29013,N_28982);
or U29313 (N_29313,N_29069,N_29077);
and U29314 (N_29314,N_28860,N_28927);
xor U29315 (N_29315,N_28897,N_29021);
nor U29316 (N_29316,N_29086,N_28893);
nor U29317 (N_29317,N_28938,N_29007);
or U29318 (N_29318,N_28984,N_29019);
nand U29319 (N_29319,N_29010,N_28887);
nand U29320 (N_29320,N_28888,N_29083);
and U29321 (N_29321,N_29084,N_29033);
nor U29322 (N_29322,N_28988,N_28848);
or U29323 (N_29323,N_28918,N_28971);
nor U29324 (N_29324,N_28963,N_28905);
nand U29325 (N_29325,N_29069,N_28988);
xnor U29326 (N_29326,N_29088,N_29032);
nor U29327 (N_29327,N_28963,N_28852);
and U29328 (N_29328,N_28893,N_29062);
or U29329 (N_29329,N_28873,N_28887);
or U29330 (N_29330,N_28833,N_29000);
nor U29331 (N_29331,N_28950,N_29084);
and U29332 (N_29332,N_28858,N_28859);
or U29333 (N_29333,N_29068,N_28966);
nor U29334 (N_29334,N_28877,N_29005);
nor U29335 (N_29335,N_29076,N_29061);
nand U29336 (N_29336,N_28996,N_29059);
nor U29337 (N_29337,N_28806,N_28994);
and U29338 (N_29338,N_28898,N_29070);
nor U29339 (N_29339,N_29016,N_29075);
nor U29340 (N_29340,N_29062,N_28810);
xor U29341 (N_29341,N_28953,N_28801);
nand U29342 (N_29342,N_28855,N_29034);
xor U29343 (N_29343,N_29058,N_28960);
xnor U29344 (N_29344,N_28883,N_29095);
nor U29345 (N_29345,N_28871,N_29077);
or U29346 (N_29346,N_29073,N_29028);
and U29347 (N_29347,N_28999,N_28972);
or U29348 (N_29348,N_28943,N_28978);
and U29349 (N_29349,N_28803,N_28991);
nand U29350 (N_29350,N_29073,N_28970);
or U29351 (N_29351,N_28890,N_28969);
nand U29352 (N_29352,N_29088,N_28868);
and U29353 (N_29353,N_29025,N_29027);
or U29354 (N_29354,N_28832,N_28886);
or U29355 (N_29355,N_28815,N_29088);
and U29356 (N_29356,N_28815,N_28943);
nand U29357 (N_29357,N_28902,N_29026);
xor U29358 (N_29358,N_28834,N_28976);
or U29359 (N_29359,N_28957,N_28942);
xnor U29360 (N_29360,N_28825,N_29072);
nand U29361 (N_29361,N_28998,N_28839);
xnor U29362 (N_29362,N_28862,N_28967);
xor U29363 (N_29363,N_28935,N_29001);
nor U29364 (N_29364,N_29058,N_28973);
nor U29365 (N_29365,N_28840,N_28877);
xnor U29366 (N_29366,N_28861,N_29026);
xor U29367 (N_29367,N_29017,N_28822);
or U29368 (N_29368,N_28948,N_28868);
xnor U29369 (N_29369,N_28940,N_29056);
xnor U29370 (N_29370,N_28956,N_28947);
xnor U29371 (N_29371,N_28984,N_29092);
nor U29372 (N_29372,N_28878,N_28829);
and U29373 (N_29373,N_29011,N_29006);
and U29374 (N_29374,N_28809,N_28878);
xnor U29375 (N_29375,N_28987,N_29066);
and U29376 (N_29376,N_29062,N_28960);
or U29377 (N_29377,N_28810,N_28856);
nor U29378 (N_29378,N_29059,N_28966);
nor U29379 (N_29379,N_28970,N_28826);
nor U29380 (N_29380,N_29012,N_29018);
nor U29381 (N_29381,N_29080,N_28985);
or U29382 (N_29382,N_28941,N_28976);
or U29383 (N_29383,N_28969,N_28898);
nor U29384 (N_29384,N_28936,N_29072);
and U29385 (N_29385,N_28995,N_29008);
and U29386 (N_29386,N_29011,N_29055);
nor U29387 (N_29387,N_29013,N_29015);
nand U29388 (N_29388,N_28825,N_29005);
xnor U29389 (N_29389,N_28886,N_28804);
nand U29390 (N_29390,N_28969,N_28887);
or U29391 (N_29391,N_28904,N_28900);
xor U29392 (N_29392,N_28831,N_29031);
xor U29393 (N_29393,N_29053,N_28867);
nor U29394 (N_29394,N_28851,N_29098);
nand U29395 (N_29395,N_29085,N_29010);
or U29396 (N_29396,N_29035,N_28867);
or U29397 (N_29397,N_29007,N_29008);
nand U29398 (N_29398,N_28871,N_28880);
and U29399 (N_29399,N_29058,N_28956);
and U29400 (N_29400,N_29267,N_29231);
xnor U29401 (N_29401,N_29192,N_29165);
or U29402 (N_29402,N_29246,N_29304);
xor U29403 (N_29403,N_29268,N_29162);
nand U29404 (N_29404,N_29291,N_29187);
xnor U29405 (N_29405,N_29326,N_29128);
or U29406 (N_29406,N_29196,N_29110);
nand U29407 (N_29407,N_29101,N_29182);
nand U29408 (N_29408,N_29360,N_29365);
and U29409 (N_29409,N_29315,N_29371);
nor U29410 (N_29410,N_29299,N_29166);
xnor U29411 (N_29411,N_29153,N_29222);
nand U29412 (N_29412,N_29236,N_29136);
xor U29413 (N_29413,N_29366,N_29282);
and U29414 (N_29414,N_29381,N_29240);
xor U29415 (N_29415,N_29188,N_29105);
and U29416 (N_29416,N_29145,N_29120);
xnor U29417 (N_29417,N_29241,N_29249);
xor U29418 (N_29418,N_29102,N_29167);
or U29419 (N_29419,N_29151,N_29221);
or U29420 (N_29420,N_29296,N_29184);
or U29421 (N_29421,N_29270,N_29186);
or U29422 (N_29422,N_29312,N_29100);
nor U29423 (N_29423,N_29223,N_29287);
nand U29424 (N_29424,N_29321,N_29212);
and U29425 (N_29425,N_29252,N_29313);
and U29426 (N_29426,N_29301,N_29297);
or U29427 (N_29427,N_29202,N_29256);
and U29428 (N_29428,N_29342,N_29379);
nor U29429 (N_29429,N_29131,N_29298);
nor U29430 (N_29430,N_29335,N_29199);
or U29431 (N_29431,N_29115,N_29230);
and U29432 (N_29432,N_29229,N_29107);
nand U29433 (N_29433,N_29354,N_29149);
or U29434 (N_29434,N_29311,N_29349);
or U29435 (N_29435,N_29373,N_29344);
nor U29436 (N_29436,N_29109,N_29302);
xor U29437 (N_29437,N_29370,N_29262);
or U29438 (N_29438,N_29164,N_29198);
or U29439 (N_29439,N_29314,N_29347);
xor U29440 (N_29440,N_29398,N_29260);
nand U29441 (N_29441,N_29111,N_29168);
and U29442 (N_29442,N_29396,N_29190);
nor U29443 (N_29443,N_29332,N_29169);
or U29444 (N_29444,N_29320,N_29272);
nand U29445 (N_29445,N_29113,N_29132);
or U29446 (N_29446,N_29234,N_29263);
nor U29447 (N_29447,N_29306,N_29337);
nand U29448 (N_29448,N_29159,N_29123);
nor U29449 (N_29449,N_29243,N_29285);
nor U29450 (N_29450,N_29181,N_29305);
nand U29451 (N_29451,N_29141,N_29194);
and U29452 (N_29452,N_29170,N_29351);
nor U29453 (N_29453,N_29137,N_29280);
nor U29454 (N_29454,N_29108,N_29389);
nand U29455 (N_29455,N_29255,N_29248);
nand U29456 (N_29456,N_29395,N_29226);
or U29457 (N_29457,N_29308,N_29251);
nor U29458 (N_29458,N_29247,N_29121);
nand U29459 (N_29459,N_29380,N_29334);
nand U29460 (N_29460,N_29237,N_29368);
or U29461 (N_29461,N_29144,N_29265);
nand U29462 (N_29462,N_29340,N_29235);
nand U29463 (N_29463,N_29300,N_29205);
nand U29464 (N_29464,N_29195,N_29264);
nand U29465 (N_29465,N_29173,N_29273);
xor U29466 (N_29466,N_29220,N_29177);
nor U29467 (N_29467,N_29322,N_29390);
nor U29468 (N_29468,N_29375,N_29204);
and U29469 (N_29469,N_29271,N_29218);
nand U29470 (N_29470,N_29376,N_29250);
xor U29471 (N_29471,N_29112,N_29135);
and U29472 (N_29472,N_29118,N_29388);
xor U29473 (N_29473,N_29327,N_29382);
and U29474 (N_29474,N_29261,N_29139);
xor U29475 (N_29475,N_29233,N_29348);
or U29476 (N_29476,N_29127,N_29309);
nor U29477 (N_29477,N_29362,N_29152);
nor U29478 (N_29478,N_29384,N_29274);
and U29479 (N_29479,N_29155,N_29179);
nand U29480 (N_29480,N_29180,N_29171);
nand U29481 (N_29481,N_29355,N_29392);
nand U29482 (N_29482,N_29232,N_29129);
nand U29483 (N_29483,N_29269,N_29385);
or U29484 (N_29484,N_29160,N_29161);
and U29485 (N_29485,N_29259,N_29275);
nor U29486 (N_29486,N_29193,N_29213);
nor U29487 (N_29487,N_29116,N_29174);
nor U29488 (N_29488,N_29185,N_29266);
xnor U29489 (N_29489,N_29352,N_29393);
and U29490 (N_29490,N_29253,N_29245);
nand U29491 (N_29491,N_29117,N_29227);
and U29492 (N_29492,N_29286,N_29143);
xnor U29493 (N_29493,N_29377,N_29200);
nand U29494 (N_29494,N_29276,N_29224);
xor U29495 (N_29495,N_29345,N_29387);
and U29496 (N_29496,N_29364,N_29317);
xnor U29497 (N_29497,N_29356,N_29238);
nand U29498 (N_29498,N_29397,N_29146);
nand U29499 (N_29499,N_29318,N_29336);
nand U29500 (N_29500,N_29353,N_29244);
xor U29501 (N_29501,N_29103,N_29239);
nor U29502 (N_29502,N_29319,N_29242);
and U29503 (N_29503,N_29358,N_29210);
nand U29504 (N_29504,N_29333,N_29122);
and U29505 (N_29505,N_29175,N_29359);
and U29506 (N_29506,N_29189,N_29329);
or U29507 (N_29507,N_29214,N_29134);
xor U29508 (N_29508,N_29293,N_29346);
nand U29509 (N_29509,N_29154,N_29125);
nand U29510 (N_29510,N_29391,N_29126);
and U29511 (N_29511,N_29324,N_29206);
xnor U29512 (N_29512,N_29367,N_29119);
nand U29513 (N_29513,N_29357,N_29258);
xnor U29514 (N_29514,N_29330,N_29219);
nor U29515 (N_29515,N_29209,N_29277);
nand U29516 (N_29516,N_29254,N_29303);
and U29517 (N_29517,N_29156,N_29140);
or U29518 (N_29518,N_29292,N_29215);
nor U29519 (N_29519,N_29383,N_29289);
xor U29520 (N_29520,N_29399,N_29361);
and U29521 (N_29521,N_29207,N_29148);
and U29522 (N_29522,N_29130,N_29114);
xnor U29523 (N_29523,N_29147,N_29307);
xnor U29524 (N_29524,N_29158,N_29104);
or U29525 (N_29525,N_29176,N_29203);
nand U29526 (N_29526,N_29339,N_29197);
nand U29527 (N_29527,N_29183,N_29283);
and U29528 (N_29528,N_29284,N_29257);
nor U29529 (N_29529,N_29372,N_29394);
or U29530 (N_29530,N_29201,N_29216);
xor U29531 (N_29531,N_29150,N_29281);
nand U29532 (N_29532,N_29378,N_29295);
and U29533 (N_29533,N_29279,N_29386);
and U29534 (N_29534,N_29369,N_29191);
xnor U29535 (N_29535,N_29374,N_29228);
xor U29536 (N_29536,N_29350,N_29323);
nand U29537 (N_29537,N_29328,N_29178);
xnor U29538 (N_29538,N_29310,N_29225);
nand U29539 (N_29539,N_29363,N_29290);
nand U29540 (N_29540,N_29325,N_29338);
or U29541 (N_29541,N_29138,N_29124);
and U29542 (N_29542,N_29157,N_29294);
xnor U29543 (N_29543,N_29172,N_29278);
nand U29544 (N_29544,N_29211,N_29343);
or U29545 (N_29545,N_29142,N_29208);
nor U29546 (N_29546,N_29331,N_29316);
nand U29547 (N_29547,N_29133,N_29341);
nor U29548 (N_29548,N_29106,N_29217);
xor U29549 (N_29549,N_29163,N_29288);
nand U29550 (N_29550,N_29187,N_29399);
xnor U29551 (N_29551,N_29328,N_29341);
xor U29552 (N_29552,N_29330,N_29151);
or U29553 (N_29553,N_29327,N_29388);
nor U29554 (N_29554,N_29376,N_29120);
nor U29555 (N_29555,N_29364,N_29279);
and U29556 (N_29556,N_29239,N_29371);
xor U29557 (N_29557,N_29389,N_29394);
xnor U29558 (N_29558,N_29277,N_29352);
or U29559 (N_29559,N_29369,N_29372);
nand U29560 (N_29560,N_29199,N_29323);
nor U29561 (N_29561,N_29317,N_29280);
nor U29562 (N_29562,N_29365,N_29265);
and U29563 (N_29563,N_29199,N_29282);
or U29564 (N_29564,N_29389,N_29388);
nor U29565 (N_29565,N_29292,N_29272);
or U29566 (N_29566,N_29152,N_29327);
and U29567 (N_29567,N_29329,N_29246);
nand U29568 (N_29568,N_29350,N_29109);
nor U29569 (N_29569,N_29139,N_29228);
or U29570 (N_29570,N_29211,N_29333);
and U29571 (N_29571,N_29295,N_29353);
nor U29572 (N_29572,N_29158,N_29349);
nand U29573 (N_29573,N_29344,N_29141);
xor U29574 (N_29574,N_29205,N_29346);
nand U29575 (N_29575,N_29206,N_29190);
or U29576 (N_29576,N_29344,N_29289);
or U29577 (N_29577,N_29281,N_29214);
nand U29578 (N_29578,N_29359,N_29304);
or U29579 (N_29579,N_29290,N_29263);
nand U29580 (N_29580,N_29245,N_29151);
or U29581 (N_29581,N_29186,N_29276);
xor U29582 (N_29582,N_29308,N_29288);
and U29583 (N_29583,N_29237,N_29355);
xnor U29584 (N_29584,N_29309,N_29391);
nand U29585 (N_29585,N_29160,N_29359);
nor U29586 (N_29586,N_29230,N_29302);
xnor U29587 (N_29587,N_29367,N_29347);
nor U29588 (N_29588,N_29361,N_29172);
nor U29589 (N_29589,N_29327,N_29106);
or U29590 (N_29590,N_29137,N_29346);
nor U29591 (N_29591,N_29269,N_29175);
or U29592 (N_29592,N_29228,N_29158);
nor U29593 (N_29593,N_29336,N_29373);
xnor U29594 (N_29594,N_29386,N_29376);
and U29595 (N_29595,N_29179,N_29307);
or U29596 (N_29596,N_29310,N_29151);
xor U29597 (N_29597,N_29175,N_29361);
or U29598 (N_29598,N_29143,N_29160);
nand U29599 (N_29599,N_29232,N_29285);
xor U29600 (N_29600,N_29224,N_29283);
and U29601 (N_29601,N_29361,N_29290);
nand U29602 (N_29602,N_29240,N_29300);
nand U29603 (N_29603,N_29236,N_29174);
and U29604 (N_29604,N_29233,N_29211);
nor U29605 (N_29605,N_29226,N_29349);
xnor U29606 (N_29606,N_29389,N_29237);
nand U29607 (N_29607,N_29299,N_29277);
nor U29608 (N_29608,N_29162,N_29184);
nand U29609 (N_29609,N_29359,N_29390);
nand U29610 (N_29610,N_29190,N_29384);
xor U29611 (N_29611,N_29107,N_29117);
nand U29612 (N_29612,N_29184,N_29219);
nor U29613 (N_29613,N_29171,N_29187);
xor U29614 (N_29614,N_29203,N_29159);
nand U29615 (N_29615,N_29332,N_29330);
and U29616 (N_29616,N_29132,N_29120);
nor U29617 (N_29617,N_29216,N_29206);
and U29618 (N_29618,N_29367,N_29212);
nand U29619 (N_29619,N_29104,N_29129);
and U29620 (N_29620,N_29102,N_29374);
and U29621 (N_29621,N_29208,N_29233);
nand U29622 (N_29622,N_29366,N_29142);
and U29623 (N_29623,N_29333,N_29256);
and U29624 (N_29624,N_29192,N_29153);
xor U29625 (N_29625,N_29103,N_29234);
xor U29626 (N_29626,N_29367,N_29165);
xnor U29627 (N_29627,N_29155,N_29246);
or U29628 (N_29628,N_29293,N_29396);
nor U29629 (N_29629,N_29196,N_29398);
xnor U29630 (N_29630,N_29104,N_29124);
nand U29631 (N_29631,N_29228,N_29281);
nor U29632 (N_29632,N_29216,N_29120);
and U29633 (N_29633,N_29132,N_29364);
nand U29634 (N_29634,N_29317,N_29363);
xnor U29635 (N_29635,N_29201,N_29312);
or U29636 (N_29636,N_29283,N_29138);
or U29637 (N_29637,N_29169,N_29339);
xor U29638 (N_29638,N_29196,N_29371);
xnor U29639 (N_29639,N_29299,N_29230);
nand U29640 (N_29640,N_29253,N_29290);
and U29641 (N_29641,N_29320,N_29188);
nor U29642 (N_29642,N_29391,N_29268);
and U29643 (N_29643,N_29342,N_29163);
and U29644 (N_29644,N_29388,N_29165);
xor U29645 (N_29645,N_29228,N_29283);
and U29646 (N_29646,N_29315,N_29350);
nor U29647 (N_29647,N_29150,N_29342);
nor U29648 (N_29648,N_29324,N_29219);
or U29649 (N_29649,N_29341,N_29124);
xor U29650 (N_29650,N_29305,N_29213);
or U29651 (N_29651,N_29171,N_29163);
and U29652 (N_29652,N_29159,N_29251);
nand U29653 (N_29653,N_29245,N_29383);
nand U29654 (N_29654,N_29215,N_29319);
nand U29655 (N_29655,N_29188,N_29144);
nand U29656 (N_29656,N_29109,N_29385);
and U29657 (N_29657,N_29356,N_29294);
or U29658 (N_29658,N_29372,N_29186);
nand U29659 (N_29659,N_29115,N_29301);
xnor U29660 (N_29660,N_29264,N_29245);
or U29661 (N_29661,N_29115,N_29117);
and U29662 (N_29662,N_29183,N_29361);
nor U29663 (N_29663,N_29144,N_29175);
or U29664 (N_29664,N_29236,N_29358);
xor U29665 (N_29665,N_29318,N_29253);
and U29666 (N_29666,N_29289,N_29208);
nor U29667 (N_29667,N_29288,N_29184);
nor U29668 (N_29668,N_29375,N_29314);
nand U29669 (N_29669,N_29245,N_29323);
nand U29670 (N_29670,N_29210,N_29142);
xor U29671 (N_29671,N_29288,N_29277);
or U29672 (N_29672,N_29198,N_29342);
xnor U29673 (N_29673,N_29370,N_29338);
or U29674 (N_29674,N_29178,N_29126);
nor U29675 (N_29675,N_29185,N_29196);
nand U29676 (N_29676,N_29214,N_29186);
and U29677 (N_29677,N_29166,N_29385);
and U29678 (N_29678,N_29214,N_29336);
and U29679 (N_29679,N_29366,N_29391);
and U29680 (N_29680,N_29212,N_29296);
and U29681 (N_29681,N_29182,N_29269);
xnor U29682 (N_29682,N_29312,N_29256);
nand U29683 (N_29683,N_29164,N_29257);
and U29684 (N_29684,N_29341,N_29305);
nor U29685 (N_29685,N_29173,N_29363);
or U29686 (N_29686,N_29354,N_29143);
or U29687 (N_29687,N_29260,N_29388);
and U29688 (N_29688,N_29394,N_29293);
xor U29689 (N_29689,N_29206,N_29385);
and U29690 (N_29690,N_29328,N_29167);
or U29691 (N_29691,N_29217,N_29134);
xnor U29692 (N_29692,N_29337,N_29244);
xnor U29693 (N_29693,N_29193,N_29267);
nor U29694 (N_29694,N_29167,N_29206);
nor U29695 (N_29695,N_29279,N_29345);
nor U29696 (N_29696,N_29308,N_29291);
nand U29697 (N_29697,N_29257,N_29340);
nand U29698 (N_29698,N_29360,N_29311);
or U29699 (N_29699,N_29225,N_29125);
and U29700 (N_29700,N_29657,N_29426);
nor U29701 (N_29701,N_29655,N_29465);
or U29702 (N_29702,N_29549,N_29524);
or U29703 (N_29703,N_29659,N_29632);
or U29704 (N_29704,N_29403,N_29439);
xor U29705 (N_29705,N_29413,N_29679);
and U29706 (N_29706,N_29479,N_29622);
and U29707 (N_29707,N_29447,N_29402);
or U29708 (N_29708,N_29652,N_29411);
nor U29709 (N_29709,N_29563,N_29467);
nand U29710 (N_29710,N_29612,N_29500);
and U29711 (N_29711,N_29685,N_29562);
xnor U29712 (N_29712,N_29627,N_29519);
xnor U29713 (N_29713,N_29607,N_29570);
and U29714 (N_29714,N_29538,N_29459);
or U29715 (N_29715,N_29661,N_29412);
or U29716 (N_29716,N_29489,N_29573);
nand U29717 (N_29717,N_29673,N_29421);
or U29718 (N_29718,N_29584,N_29490);
or U29719 (N_29719,N_29417,N_29531);
xnor U29720 (N_29720,N_29525,N_29469);
nand U29721 (N_29721,N_29414,N_29553);
and U29722 (N_29722,N_29437,N_29491);
nand U29723 (N_29723,N_29484,N_29556);
nand U29724 (N_29724,N_29463,N_29405);
and U29725 (N_29725,N_29492,N_29532);
xor U29726 (N_29726,N_29611,N_29577);
xnor U29727 (N_29727,N_29448,N_29669);
nand U29728 (N_29728,N_29460,N_29445);
nand U29729 (N_29729,N_29610,N_29505);
xor U29730 (N_29730,N_29664,N_29662);
nand U29731 (N_29731,N_29475,N_29616);
nand U29732 (N_29732,N_29508,N_29647);
nand U29733 (N_29733,N_29651,N_29520);
and U29734 (N_29734,N_29546,N_29594);
nor U29735 (N_29735,N_29613,N_29663);
and U29736 (N_29736,N_29602,N_29453);
or U29737 (N_29737,N_29540,N_29634);
and U29738 (N_29738,N_29514,N_29511);
nor U29739 (N_29739,N_29515,N_29609);
nor U29740 (N_29740,N_29404,N_29461);
nor U29741 (N_29741,N_29644,N_29588);
and U29742 (N_29742,N_29415,N_29424);
xnor U29743 (N_29743,N_29565,N_29486);
or U29744 (N_29744,N_29560,N_29471);
and U29745 (N_29745,N_29579,N_29539);
nor U29746 (N_29746,N_29686,N_29595);
nor U29747 (N_29747,N_29599,N_29674);
nor U29748 (N_29748,N_29407,N_29528);
nand U29749 (N_29749,N_29653,N_29454);
and U29750 (N_29750,N_29541,N_29537);
or U29751 (N_29751,N_29680,N_29526);
xor U29752 (N_29752,N_29433,N_29558);
or U29753 (N_29753,N_29431,N_29438);
and U29754 (N_29754,N_29681,N_29493);
and U29755 (N_29755,N_29694,N_29658);
xor U29756 (N_29756,N_29483,N_29690);
nor U29757 (N_29757,N_29498,N_29543);
and U29758 (N_29758,N_29446,N_29472);
and U29759 (N_29759,N_29585,N_29625);
and U29760 (N_29760,N_29533,N_29406);
or U29761 (N_29761,N_29614,N_29530);
nand U29762 (N_29762,N_29677,N_29555);
nand U29763 (N_29763,N_29665,N_29682);
nor U29764 (N_29764,N_29458,N_29578);
xor U29765 (N_29765,N_29637,N_29695);
and U29766 (N_29766,N_29497,N_29568);
nor U29767 (N_29767,N_29440,N_29451);
or U29768 (N_29768,N_29697,N_29518);
xnor U29769 (N_29769,N_29494,N_29473);
xor U29770 (N_29770,N_29517,N_29551);
nor U29771 (N_29771,N_29605,N_29635);
nand U29772 (N_29772,N_29660,N_29422);
and U29773 (N_29773,N_29516,N_29423);
nand U29774 (N_29774,N_29485,N_29512);
nand U29775 (N_29775,N_29425,N_29400);
and U29776 (N_29776,N_29435,N_29429);
and U29777 (N_29777,N_29643,N_29409);
or U29778 (N_29778,N_29444,N_29509);
nand U29779 (N_29779,N_29693,N_29561);
xor U29780 (N_29780,N_29496,N_29698);
or U29781 (N_29781,N_29636,N_29600);
xor U29782 (N_29782,N_29623,N_29544);
or U29783 (N_29783,N_29419,N_29676);
or U29784 (N_29784,N_29503,N_29668);
nand U29785 (N_29785,N_29615,N_29488);
and U29786 (N_29786,N_29688,N_29442);
xor U29787 (N_29787,N_29640,N_29527);
and U29788 (N_29788,N_29513,N_29649);
nand U29789 (N_29789,N_29574,N_29521);
xnor U29790 (N_29790,N_29656,N_29523);
or U29791 (N_29791,N_29645,N_29629);
and U29792 (N_29792,N_29401,N_29542);
nor U29793 (N_29793,N_29624,N_29678);
xor U29794 (N_29794,N_29481,N_29478);
nor U29795 (N_29795,N_29552,N_29443);
or U29796 (N_29796,N_29474,N_29567);
xor U29797 (N_29797,N_29672,N_29507);
nor U29798 (N_29798,N_29495,N_29621);
xor U29799 (N_29799,N_29499,N_29476);
and U29800 (N_29800,N_29452,N_29631);
nor U29801 (N_29801,N_29418,N_29432);
and U29802 (N_29802,N_29699,N_29620);
and U29803 (N_29803,N_29683,N_29482);
xnor U29804 (N_29804,N_29536,N_29641);
or U29805 (N_29805,N_29592,N_29566);
nor U29806 (N_29806,N_29630,N_29608);
nor U29807 (N_29807,N_29571,N_29687);
nor U29808 (N_29808,N_29587,N_29598);
nand U29809 (N_29809,N_29547,N_29441);
nor U29810 (N_29810,N_29572,N_29477);
xor U29811 (N_29811,N_29597,N_29638);
and U29812 (N_29812,N_29480,N_29606);
nor U29813 (N_29813,N_29589,N_29449);
xnor U29814 (N_29814,N_29675,N_29582);
or U29815 (N_29815,N_29470,N_29581);
nand U29816 (N_29816,N_29646,N_29504);
xnor U29817 (N_29817,N_29464,N_29642);
and U29818 (N_29818,N_29416,N_29569);
nor U29819 (N_29819,N_29601,N_29502);
nand U29820 (N_29820,N_29603,N_29684);
nor U29821 (N_29821,N_29576,N_29689);
nor U29822 (N_29822,N_29654,N_29466);
xor U29823 (N_29823,N_29529,N_29457);
and U29824 (N_29824,N_29639,N_29670);
xnor U29825 (N_29825,N_29691,N_29535);
xnor U29826 (N_29826,N_29450,N_29434);
and U29827 (N_29827,N_29666,N_29436);
xnor U29828 (N_29828,N_29522,N_29548);
and U29829 (N_29829,N_29667,N_29593);
nor U29830 (N_29830,N_29618,N_29408);
nor U29831 (N_29831,N_29590,N_29462);
nor U29832 (N_29832,N_29575,N_29671);
xor U29833 (N_29833,N_29510,N_29410);
or U29834 (N_29834,N_29420,N_29559);
nand U29835 (N_29835,N_29580,N_29487);
and U29836 (N_29836,N_29455,N_29648);
nor U29837 (N_29837,N_29619,N_29564);
xnor U29838 (N_29838,N_29692,N_29428);
or U29839 (N_29839,N_29545,N_29626);
nand U29840 (N_29840,N_29554,N_29583);
nor U29841 (N_29841,N_29591,N_29633);
and U29842 (N_29842,N_29650,N_29550);
nor U29843 (N_29843,N_29604,N_29534);
or U29844 (N_29844,N_29696,N_29628);
or U29845 (N_29845,N_29501,N_29557);
xnor U29846 (N_29846,N_29596,N_29427);
xnor U29847 (N_29847,N_29506,N_29468);
xnor U29848 (N_29848,N_29430,N_29586);
and U29849 (N_29849,N_29617,N_29456);
or U29850 (N_29850,N_29454,N_29548);
nor U29851 (N_29851,N_29512,N_29621);
xor U29852 (N_29852,N_29439,N_29663);
nand U29853 (N_29853,N_29645,N_29558);
nor U29854 (N_29854,N_29485,N_29460);
or U29855 (N_29855,N_29443,N_29422);
and U29856 (N_29856,N_29679,N_29509);
nor U29857 (N_29857,N_29584,N_29528);
nand U29858 (N_29858,N_29667,N_29431);
xnor U29859 (N_29859,N_29607,N_29434);
nor U29860 (N_29860,N_29456,N_29620);
or U29861 (N_29861,N_29542,N_29474);
or U29862 (N_29862,N_29623,N_29511);
or U29863 (N_29863,N_29606,N_29602);
and U29864 (N_29864,N_29670,N_29581);
xor U29865 (N_29865,N_29552,N_29534);
or U29866 (N_29866,N_29499,N_29562);
nand U29867 (N_29867,N_29452,N_29546);
nand U29868 (N_29868,N_29512,N_29490);
and U29869 (N_29869,N_29467,N_29591);
xor U29870 (N_29870,N_29620,N_29471);
or U29871 (N_29871,N_29410,N_29662);
xnor U29872 (N_29872,N_29659,N_29638);
and U29873 (N_29873,N_29417,N_29641);
nand U29874 (N_29874,N_29568,N_29493);
or U29875 (N_29875,N_29639,N_29619);
nand U29876 (N_29876,N_29429,N_29614);
or U29877 (N_29877,N_29686,N_29488);
nor U29878 (N_29878,N_29529,N_29404);
or U29879 (N_29879,N_29413,N_29602);
xnor U29880 (N_29880,N_29658,N_29415);
and U29881 (N_29881,N_29678,N_29413);
nor U29882 (N_29882,N_29477,N_29548);
or U29883 (N_29883,N_29658,N_29513);
and U29884 (N_29884,N_29436,N_29421);
nor U29885 (N_29885,N_29593,N_29572);
and U29886 (N_29886,N_29679,N_29665);
nand U29887 (N_29887,N_29426,N_29667);
nand U29888 (N_29888,N_29642,N_29623);
or U29889 (N_29889,N_29595,N_29612);
nand U29890 (N_29890,N_29477,N_29411);
nand U29891 (N_29891,N_29549,N_29633);
and U29892 (N_29892,N_29405,N_29495);
or U29893 (N_29893,N_29480,N_29436);
xnor U29894 (N_29894,N_29407,N_29643);
nor U29895 (N_29895,N_29436,N_29598);
and U29896 (N_29896,N_29662,N_29538);
xor U29897 (N_29897,N_29551,N_29651);
or U29898 (N_29898,N_29533,N_29412);
nor U29899 (N_29899,N_29587,N_29538);
nand U29900 (N_29900,N_29549,N_29459);
nand U29901 (N_29901,N_29407,N_29693);
nor U29902 (N_29902,N_29641,N_29412);
nor U29903 (N_29903,N_29499,N_29418);
xor U29904 (N_29904,N_29601,N_29665);
nor U29905 (N_29905,N_29671,N_29494);
nand U29906 (N_29906,N_29407,N_29478);
or U29907 (N_29907,N_29509,N_29664);
nand U29908 (N_29908,N_29598,N_29507);
xor U29909 (N_29909,N_29657,N_29455);
nand U29910 (N_29910,N_29471,N_29497);
nor U29911 (N_29911,N_29459,N_29601);
nand U29912 (N_29912,N_29683,N_29571);
or U29913 (N_29913,N_29676,N_29588);
nand U29914 (N_29914,N_29460,N_29680);
and U29915 (N_29915,N_29576,N_29634);
and U29916 (N_29916,N_29593,N_29458);
and U29917 (N_29917,N_29530,N_29499);
and U29918 (N_29918,N_29470,N_29516);
xnor U29919 (N_29919,N_29441,N_29420);
xnor U29920 (N_29920,N_29433,N_29544);
xor U29921 (N_29921,N_29610,N_29680);
and U29922 (N_29922,N_29653,N_29499);
and U29923 (N_29923,N_29587,N_29629);
nand U29924 (N_29924,N_29613,N_29558);
nor U29925 (N_29925,N_29594,N_29595);
nor U29926 (N_29926,N_29664,N_29408);
and U29927 (N_29927,N_29672,N_29511);
or U29928 (N_29928,N_29537,N_29678);
xor U29929 (N_29929,N_29503,N_29491);
and U29930 (N_29930,N_29655,N_29539);
nor U29931 (N_29931,N_29469,N_29635);
nand U29932 (N_29932,N_29451,N_29691);
nand U29933 (N_29933,N_29413,N_29616);
and U29934 (N_29934,N_29503,N_29580);
xor U29935 (N_29935,N_29585,N_29565);
nand U29936 (N_29936,N_29407,N_29672);
and U29937 (N_29937,N_29604,N_29653);
or U29938 (N_29938,N_29594,N_29538);
and U29939 (N_29939,N_29541,N_29548);
xnor U29940 (N_29940,N_29532,N_29645);
xor U29941 (N_29941,N_29647,N_29541);
nand U29942 (N_29942,N_29615,N_29618);
xor U29943 (N_29943,N_29457,N_29548);
and U29944 (N_29944,N_29487,N_29515);
xor U29945 (N_29945,N_29489,N_29599);
nor U29946 (N_29946,N_29452,N_29470);
nor U29947 (N_29947,N_29538,N_29656);
and U29948 (N_29948,N_29481,N_29413);
xor U29949 (N_29949,N_29501,N_29462);
or U29950 (N_29950,N_29560,N_29456);
and U29951 (N_29951,N_29420,N_29447);
xor U29952 (N_29952,N_29621,N_29433);
nand U29953 (N_29953,N_29447,N_29623);
nand U29954 (N_29954,N_29506,N_29679);
xnor U29955 (N_29955,N_29644,N_29685);
and U29956 (N_29956,N_29495,N_29575);
xor U29957 (N_29957,N_29536,N_29437);
and U29958 (N_29958,N_29553,N_29673);
or U29959 (N_29959,N_29575,N_29423);
and U29960 (N_29960,N_29606,N_29637);
nand U29961 (N_29961,N_29508,N_29597);
or U29962 (N_29962,N_29606,N_29641);
xnor U29963 (N_29963,N_29480,N_29657);
nor U29964 (N_29964,N_29501,N_29450);
and U29965 (N_29965,N_29440,N_29643);
nand U29966 (N_29966,N_29601,N_29667);
nor U29967 (N_29967,N_29438,N_29430);
or U29968 (N_29968,N_29632,N_29531);
xnor U29969 (N_29969,N_29465,N_29563);
and U29970 (N_29970,N_29491,N_29623);
and U29971 (N_29971,N_29456,N_29669);
or U29972 (N_29972,N_29509,N_29576);
nand U29973 (N_29973,N_29584,N_29549);
and U29974 (N_29974,N_29687,N_29517);
xor U29975 (N_29975,N_29482,N_29425);
nand U29976 (N_29976,N_29443,N_29650);
and U29977 (N_29977,N_29536,N_29697);
or U29978 (N_29978,N_29448,N_29414);
or U29979 (N_29979,N_29492,N_29677);
or U29980 (N_29980,N_29439,N_29656);
xnor U29981 (N_29981,N_29485,N_29544);
and U29982 (N_29982,N_29409,N_29644);
or U29983 (N_29983,N_29575,N_29428);
nor U29984 (N_29984,N_29636,N_29575);
nor U29985 (N_29985,N_29431,N_29467);
or U29986 (N_29986,N_29484,N_29657);
and U29987 (N_29987,N_29464,N_29692);
xnor U29988 (N_29988,N_29432,N_29498);
xnor U29989 (N_29989,N_29420,N_29692);
nand U29990 (N_29990,N_29422,N_29500);
nor U29991 (N_29991,N_29474,N_29539);
or U29992 (N_29992,N_29669,N_29466);
or U29993 (N_29993,N_29525,N_29688);
or U29994 (N_29994,N_29486,N_29620);
nor U29995 (N_29995,N_29531,N_29658);
xor U29996 (N_29996,N_29473,N_29698);
nand U29997 (N_29997,N_29681,N_29581);
or U29998 (N_29998,N_29473,N_29633);
nand U29999 (N_29999,N_29584,N_29681);
xnor UO_0 (O_0,N_29913,N_29800);
nor UO_1 (O_1,N_29790,N_29880);
or UO_2 (O_2,N_29817,N_29806);
and UO_3 (O_3,N_29979,N_29931);
nand UO_4 (O_4,N_29751,N_29706);
or UO_5 (O_5,N_29703,N_29992);
xor UO_6 (O_6,N_29912,N_29918);
or UO_7 (O_7,N_29968,N_29782);
nor UO_8 (O_8,N_29711,N_29948);
nand UO_9 (O_9,N_29940,N_29828);
and UO_10 (O_10,N_29971,N_29887);
nor UO_11 (O_11,N_29893,N_29783);
nand UO_12 (O_12,N_29795,N_29770);
or UO_13 (O_13,N_29883,N_29830);
nand UO_14 (O_14,N_29869,N_29856);
nand UO_15 (O_15,N_29753,N_29889);
and UO_16 (O_16,N_29901,N_29841);
nand UO_17 (O_17,N_29779,N_29728);
nand UO_18 (O_18,N_29888,N_29808);
xor UO_19 (O_19,N_29758,N_29951);
and UO_20 (O_20,N_29952,N_29861);
or UO_21 (O_21,N_29851,N_29941);
and UO_22 (O_22,N_29932,N_29936);
nand UO_23 (O_23,N_29812,N_29911);
nor UO_24 (O_24,N_29700,N_29917);
and UO_25 (O_25,N_29972,N_29966);
nand UO_26 (O_26,N_29881,N_29767);
and UO_27 (O_27,N_29985,N_29738);
or UO_28 (O_28,N_29787,N_29963);
and UO_29 (O_29,N_29723,N_29839);
or UO_30 (O_30,N_29866,N_29965);
nand UO_31 (O_31,N_29848,N_29857);
or UO_32 (O_32,N_29704,N_29772);
and UO_33 (O_33,N_29759,N_29914);
or UO_34 (O_34,N_29967,N_29879);
or UO_35 (O_35,N_29983,N_29908);
nand UO_36 (O_36,N_29986,N_29742);
and UO_37 (O_37,N_29850,N_29944);
nand UO_38 (O_38,N_29764,N_29873);
xnor UO_39 (O_39,N_29720,N_29902);
xnor UO_40 (O_40,N_29892,N_29988);
or UO_41 (O_41,N_29993,N_29752);
and UO_42 (O_42,N_29962,N_29803);
nand UO_43 (O_43,N_29835,N_29785);
xor UO_44 (O_44,N_29725,N_29786);
or UO_45 (O_45,N_29845,N_29766);
xor UO_46 (O_46,N_29981,N_29847);
or UO_47 (O_47,N_29721,N_29777);
nor UO_48 (O_48,N_29707,N_29836);
and UO_49 (O_49,N_29823,N_29815);
nor UO_50 (O_50,N_29862,N_29852);
nor UO_51 (O_51,N_29921,N_29860);
xor UO_52 (O_52,N_29942,N_29740);
xor UO_53 (O_53,N_29778,N_29977);
xnor UO_54 (O_54,N_29957,N_29891);
xor UO_55 (O_55,N_29953,N_29833);
and UO_56 (O_56,N_29987,N_29905);
or UO_57 (O_57,N_29925,N_29959);
and UO_58 (O_58,N_29810,N_29727);
xnor UO_59 (O_59,N_29820,N_29804);
and UO_60 (O_60,N_29989,N_29747);
or UO_61 (O_61,N_29995,N_29716);
or UO_62 (O_62,N_29710,N_29745);
xnor UO_63 (O_63,N_29754,N_29875);
nor UO_64 (O_64,N_29784,N_29762);
or UO_65 (O_65,N_29884,N_29943);
or UO_66 (O_66,N_29749,N_29975);
and UO_67 (O_67,N_29739,N_29829);
nor UO_68 (O_68,N_29882,N_29874);
and UO_69 (O_69,N_29909,N_29982);
xnor UO_70 (O_70,N_29964,N_29724);
xor UO_71 (O_71,N_29717,N_29990);
or UO_72 (O_72,N_29868,N_29791);
and UO_73 (O_73,N_29765,N_29726);
nor UO_74 (O_74,N_29924,N_29744);
nor UO_75 (O_75,N_29736,N_29781);
nand UO_76 (O_76,N_29886,N_29872);
or UO_77 (O_77,N_29788,N_29903);
xor UO_78 (O_78,N_29870,N_29926);
xnor UO_79 (O_79,N_29928,N_29761);
or UO_80 (O_80,N_29947,N_29796);
and UO_81 (O_81,N_29984,N_29970);
or UO_82 (O_82,N_29755,N_29929);
and UO_83 (O_83,N_29709,N_29712);
nor UO_84 (O_84,N_29974,N_29865);
and UO_85 (O_85,N_29999,N_29771);
or UO_86 (O_86,N_29818,N_29780);
and UO_87 (O_87,N_29821,N_29976);
nor UO_88 (O_88,N_29853,N_29877);
or UO_89 (O_89,N_29998,N_29774);
nor UO_90 (O_90,N_29705,N_29846);
nand UO_91 (O_91,N_29816,N_29714);
nand UO_92 (O_92,N_29991,N_29960);
nand UO_93 (O_93,N_29849,N_29937);
and UO_94 (O_94,N_29916,N_29878);
or UO_95 (O_95,N_29825,N_29819);
xnor UO_96 (O_96,N_29933,N_29867);
xor UO_97 (O_97,N_29732,N_29797);
nand UO_98 (O_98,N_29813,N_29843);
nand UO_99 (O_99,N_29980,N_29743);
and UO_100 (O_100,N_29805,N_29904);
nand UO_101 (O_101,N_29834,N_29831);
nor UO_102 (O_102,N_29954,N_29713);
or UO_103 (O_103,N_29827,N_29802);
xor UO_104 (O_104,N_29708,N_29915);
nor UO_105 (O_105,N_29961,N_29876);
xnor UO_106 (O_106,N_29792,N_29773);
and UO_107 (O_107,N_29899,N_29768);
nand UO_108 (O_108,N_29859,N_29927);
or UO_109 (O_109,N_29840,N_29898);
xor UO_110 (O_110,N_29956,N_29864);
nor UO_111 (O_111,N_29934,N_29730);
nor UO_112 (O_112,N_29731,N_29789);
xor UO_113 (O_113,N_29939,N_29997);
nand UO_114 (O_114,N_29969,N_29793);
nor UO_115 (O_115,N_29894,N_29702);
xor UO_116 (O_116,N_29734,N_29896);
xnor UO_117 (O_117,N_29842,N_29871);
xor UO_118 (O_118,N_29798,N_29920);
nor UO_119 (O_119,N_29973,N_29722);
or UO_120 (O_120,N_29855,N_29701);
xnor UO_121 (O_121,N_29776,N_29822);
and UO_122 (O_122,N_29757,N_29919);
and UO_123 (O_123,N_29946,N_29938);
and UO_124 (O_124,N_29824,N_29885);
or UO_125 (O_125,N_29814,N_29923);
nand UO_126 (O_126,N_29719,N_29858);
xnor UO_127 (O_127,N_29958,N_29763);
xnor UO_128 (O_128,N_29729,N_29832);
nand UO_129 (O_129,N_29950,N_29996);
xnor UO_130 (O_130,N_29733,N_29854);
or UO_131 (O_131,N_29741,N_29801);
nor UO_132 (O_132,N_29863,N_29922);
nand UO_133 (O_133,N_29907,N_29735);
or UO_134 (O_134,N_29978,N_29750);
xnor UO_135 (O_135,N_29910,N_29844);
or UO_136 (O_136,N_29811,N_29715);
or UO_137 (O_137,N_29897,N_29769);
nor UO_138 (O_138,N_29994,N_29838);
xor UO_139 (O_139,N_29746,N_29930);
nor UO_140 (O_140,N_29826,N_29748);
nand UO_141 (O_141,N_29890,N_29807);
xor UO_142 (O_142,N_29945,N_29949);
and UO_143 (O_143,N_29718,N_29809);
nand UO_144 (O_144,N_29895,N_29760);
xnor UO_145 (O_145,N_29900,N_29955);
xnor UO_146 (O_146,N_29794,N_29775);
nor UO_147 (O_147,N_29799,N_29756);
and UO_148 (O_148,N_29935,N_29837);
and UO_149 (O_149,N_29906,N_29737);
nand UO_150 (O_150,N_29874,N_29819);
or UO_151 (O_151,N_29722,N_29962);
nand UO_152 (O_152,N_29883,N_29820);
and UO_153 (O_153,N_29757,N_29819);
nor UO_154 (O_154,N_29734,N_29938);
xnor UO_155 (O_155,N_29759,N_29794);
or UO_156 (O_156,N_29941,N_29944);
and UO_157 (O_157,N_29783,N_29845);
nor UO_158 (O_158,N_29803,N_29880);
xnor UO_159 (O_159,N_29730,N_29770);
xor UO_160 (O_160,N_29919,N_29855);
xnor UO_161 (O_161,N_29793,N_29840);
or UO_162 (O_162,N_29856,N_29798);
xor UO_163 (O_163,N_29828,N_29705);
nor UO_164 (O_164,N_29793,N_29855);
xor UO_165 (O_165,N_29907,N_29714);
xnor UO_166 (O_166,N_29941,N_29959);
nor UO_167 (O_167,N_29832,N_29919);
or UO_168 (O_168,N_29808,N_29877);
nand UO_169 (O_169,N_29877,N_29865);
xnor UO_170 (O_170,N_29991,N_29961);
and UO_171 (O_171,N_29844,N_29799);
and UO_172 (O_172,N_29723,N_29712);
nor UO_173 (O_173,N_29777,N_29999);
xor UO_174 (O_174,N_29957,N_29860);
xor UO_175 (O_175,N_29779,N_29924);
or UO_176 (O_176,N_29792,N_29767);
nand UO_177 (O_177,N_29989,N_29746);
xnor UO_178 (O_178,N_29946,N_29953);
nor UO_179 (O_179,N_29714,N_29954);
and UO_180 (O_180,N_29864,N_29822);
and UO_181 (O_181,N_29925,N_29845);
xor UO_182 (O_182,N_29927,N_29940);
and UO_183 (O_183,N_29907,N_29956);
or UO_184 (O_184,N_29972,N_29810);
nand UO_185 (O_185,N_29815,N_29897);
nor UO_186 (O_186,N_29955,N_29945);
xor UO_187 (O_187,N_29944,N_29758);
xor UO_188 (O_188,N_29858,N_29986);
nor UO_189 (O_189,N_29915,N_29948);
and UO_190 (O_190,N_29844,N_29725);
xnor UO_191 (O_191,N_29799,N_29859);
nand UO_192 (O_192,N_29837,N_29744);
or UO_193 (O_193,N_29733,N_29873);
nand UO_194 (O_194,N_29974,N_29774);
and UO_195 (O_195,N_29958,N_29971);
and UO_196 (O_196,N_29946,N_29812);
xor UO_197 (O_197,N_29761,N_29944);
nor UO_198 (O_198,N_29925,N_29835);
xnor UO_199 (O_199,N_29998,N_29777);
and UO_200 (O_200,N_29943,N_29767);
xor UO_201 (O_201,N_29728,N_29864);
or UO_202 (O_202,N_29765,N_29782);
nand UO_203 (O_203,N_29931,N_29973);
nand UO_204 (O_204,N_29841,N_29731);
and UO_205 (O_205,N_29943,N_29950);
or UO_206 (O_206,N_29720,N_29741);
and UO_207 (O_207,N_29985,N_29974);
and UO_208 (O_208,N_29894,N_29965);
nand UO_209 (O_209,N_29998,N_29817);
or UO_210 (O_210,N_29956,N_29838);
and UO_211 (O_211,N_29981,N_29839);
and UO_212 (O_212,N_29728,N_29756);
nor UO_213 (O_213,N_29945,N_29805);
and UO_214 (O_214,N_29820,N_29939);
or UO_215 (O_215,N_29969,N_29999);
nand UO_216 (O_216,N_29869,N_29803);
and UO_217 (O_217,N_29729,N_29815);
xnor UO_218 (O_218,N_29900,N_29843);
nor UO_219 (O_219,N_29707,N_29813);
or UO_220 (O_220,N_29895,N_29733);
nand UO_221 (O_221,N_29851,N_29791);
nor UO_222 (O_222,N_29889,N_29830);
nor UO_223 (O_223,N_29957,N_29806);
nand UO_224 (O_224,N_29760,N_29833);
and UO_225 (O_225,N_29823,N_29808);
xnor UO_226 (O_226,N_29741,N_29952);
and UO_227 (O_227,N_29726,N_29719);
xor UO_228 (O_228,N_29841,N_29851);
nand UO_229 (O_229,N_29968,N_29766);
nand UO_230 (O_230,N_29786,N_29911);
nand UO_231 (O_231,N_29886,N_29875);
or UO_232 (O_232,N_29979,N_29901);
xnor UO_233 (O_233,N_29847,N_29701);
nand UO_234 (O_234,N_29942,N_29744);
nand UO_235 (O_235,N_29849,N_29719);
xnor UO_236 (O_236,N_29823,N_29909);
nor UO_237 (O_237,N_29785,N_29932);
nor UO_238 (O_238,N_29911,N_29731);
xnor UO_239 (O_239,N_29996,N_29983);
nand UO_240 (O_240,N_29890,N_29832);
nor UO_241 (O_241,N_29946,N_29860);
and UO_242 (O_242,N_29773,N_29946);
nand UO_243 (O_243,N_29732,N_29891);
or UO_244 (O_244,N_29731,N_29774);
nor UO_245 (O_245,N_29922,N_29902);
nand UO_246 (O_246,N_29916,N_29780);
nand UO_247 (O_247,N_29790,N_29828);
xnor UO_248 (O_248,N_29848,N_29821);
nand UO_249 (O_249,N_29948,N_29782);
and UO_250 (O_250,N_29762,N_29763);
or UO_251 (O_251,N_29871,N_29911);
nor UO_252 (O_252,N_29885,N_29805);
or UO_253 (O_253,N_29855,N_29972);
nand UO_254 (O_254,N_29921,N_29854);
nand UO_255 (O_255,N_29820,N_29863);
nor UO_256 (O_256,N_29988,N_29910);
or UO_257 (O_257,N_29831,N_29960);
and UO_258 (O_258,N_29980,N_29761);
and UO_259 (O_259,N_29793,N_29873);
xor UO_260 (O_260,N_29707,N_29802);
xor UO_261 (O_261,N_29834,N_29842);
or UO_262 (O_262,N_29807,N_29787);
and UO_263 (O_263,N_29900,N_29817);
or UO_264 (O_264,N_29775,N_29822);
and UO_265 (O_265,N_29877,N_29763);
and UO_266 (O_266,N_29908,N_29701);
xnor UO_267 (O_267,N_29791,N_29993);
nor UO_268 (O_268,N_29979,N_29875);
nand UO_269 (O_269,N_29994,N_29839);
and UO_270 (O_270,N_29717,N_29904);
nand UO_271 (O_271,N_29722,N_29834);
and UO_272 (O_272,N_29906,N_29893);
nor UO_273 (O_273,N_29897,N_29882);
xnor UO_274 (O_274,N_29754,N_29925);
nand UO_275 (O_275,N_29845,N_29765);
xor UO_276 (O_276,N_29866,N_29843);
xor UO_277 (O_277,N_29853,N_29807);
or UO_278 (O_278,N_29973,N_29846);
nor UO_279 (O_279,N_29724,N_29750);
xnor UO_280 (O_280,N_29992,N_29883);
nand UO_281 (O_281,N_29931,N_29937);
xor UO_282 (O_282,N_29888,N_29906);
nor UO_283 (O_283,N_29933,N_29888);
nor UO_284 (O_284,N_29833,N_29863);
nor UO_285 (O_285,N_29779,N_29787);
nor UO_286 (O_286,N_29939,N_29709);
nor UO_287 (O_287,N_29965,N_29760);
nor UO_288 (O_288,N_29913,N_29909);
or UO_289 (O_289,N_29738,N_29934);
xnor UO_290 (O_290,N_29975,N_29805);
or UO_291 (O_291,N_29873,N_29772);
nand UO_292 (O_292,N_29825,N_29971);
nand UO_293 (O_293,N_29915,N_29791);
nand UO_294 (O_294,N_29737,N_29948);
nor UO_295 (O_295,N_29730,N_29817);
or UO_296 (O_296,N_29765,N_29853);
nor UO_297 (O_297,N_29928,N_29856);
nand UO_298 (O_298,N_29784,N_29772);
and UO_299 (O_299,N_29792,N_29887);
xnor UO_300 (O_300,N_29966,N_29934);
nand UO_301 (O_301,N_29884,N_29923);
nand UO_302 (O_302,N_29880,N_29984);
xor UO_303 (O_303,N_29881,N_29751);
nor UO_304 (O_304,N_29983,N_29749);
or UO_305 (O_305,N_29955,N_29811);
xor UO_306 (O_306,N_29813,N_29947);
nand UO_307 (O_307,N_29929,N_29971);
or UO_308 (O_308,N_29820,N_29813);
xnor UO_309 (O_309,N_29782,N_29716);
nand UO_310 (O_310,N_29778,N_29861);
and UO_311 (O_311,N_29889,N_29874);
nand UO_312 (O_312,N_29928,N_29727);
nand UO_313 (O_313,N_29730,N_29859);
or UO_314 (O_314,N_29972,N_29981);
nand UO_315 (O_315,N_29959,N_29817);
and UO_316 (O_316,N_29984,N_29886);
or UO_317 (O_317,N_29910,N_29904);
nand UO_318 (O_318,N_29946,N_29961);
or UO_319 (O_319,N_29749,N_29967);
nand UO_320 (O_320,N_29811,N_29872);
nand UO_321 (O_321,N_29940,N_29990);
or UO_322 (O_322,N_29815,N_29940);
and UO_323 (O_323,N_29782,N_29996);
xor UO_324 (O_324,N_29829,N_29868);
xnor UO_325 (O_325,N_29823,N_29705);
and UO_326 (O_326,N_29970,N_29783);
and UO_327 (O_327,N_29960,N_29939);
nor UO_328 (O_328,N_29748,N_29739);
or UO_329 (O_329,N_29701,N_29831);
or UO_330 (O_330,N_29706,N_29869);
nand UO_331 (O_331,N_29823,N_29864);
nor UO_332 (O_332,N_29969,N_29888);
or UO_333 (O_333,N_29853,N_29968);
xor UO_334 (O_334,N_29844,N_29868);
nand UO_335 (O_335,N_29865,N_29976);
xor UO_336 (O_336,N_29775,N_29998);
or UO_337 (O_337,N_29932,N_29755);
and UO_338 (O_338,N_29750,N_29893);
xnor UO_339 (O_339,N_29894,N_29713);
xnor UO_340 (O_340,N_29751,N_29754);
nand UO_341 (O_341,N_29870,N_29906);
and UO_342 (O_342,N_29875,N_29739);
and UO_343 (O_343,N_29771,N_29868);
nor UO_344 (O_344,N_29875,N_29930);
nor UO_345 (O_345,N_29950,N_29972);
nor UO_346 (O_346,N_29898,N_29757);
nand UO_347 (O_347,N_29964,N_29820);
nand UO_348 (O_348,N_29787,N_29861);
or UO_349 (O_349,N_29709,N_29784);
nand UO_350 (O_350,N_29789,N_29849);
xnor UO_351 (O_351,N_29945,N_29975);
and UO_352 (O_352,N_29983,N_29948);
or UO_353 (O_353,N_29705,N_29840);
nand UO_354 (O_354,N_29829,N_29978);
and UO_355 (O_355,N_29888,N_29767);
nand UO_356 (O_356,N_29852,N_29908);
or UO_357 (O_357,N_29910,N_29838);
nand UO_358 (O_358,N_29774,N_29892);
or UO_359 (O_359,N_29936,N_29715);
or UO_360 (O_360,N_29730,N_29768);
nor UO_361 (O_361,N_29702,N_29782);
nor UO_362 (O_362,N_29995,N_29815);
nand UO_363 (O_363,N_29883,N_29807);
nor UO_364 (O_364,N_29918,N_29789);
xor UO_365 (O_365,N_29809,N_29864);
xor UO_366 (O_366,N_29895,N_29804);
nor UO_367 (O_367,N_29953,N_29784);
or UO_368 (O_368,N_29820,N_29938);
or UO_369 (O_369,N_29768,N_29771);
xor UO_370 (O_370,N_29952,N_29715);
and UO_371 (O_371,N_29913,N_29898);
nand UO_372 (O_372,N_29798,N_29796);
and UO_373 (O_373,N_29993,N_29772);
nor UO_374 (O_374,N_29947,N_29938);
or UO_375 (O_375,N_29837,N_29832);
xnor UO_376 (O_376,N_29812,N_29823);
xor UO_377 (O_377,N_29923,N_29813);
or UO_378 (O_378,N_29774,N_29770);
nor UO_379 (O_379,N_29982,N_29877);
and UO_380 (O_380,N_29912,N_29929);
nand UO_381 (O_381,N_29839,N_29961);
xor UO_382 (O_382,N_29747,N_29981);
or UO_383 (O_383,N_29815,N_29727);
nor UO_384 (O_384,N_29971,N_29864);
and UO_385 (O_385,N_29946,N_29838);
or UO_386 (O_386,N_29719,N_29707);
xor UO_387 (O_387,N_29919,N_29836);
nand UO_388 (O_388,N_29996,N_29846);
and UO_389 (O_389,N_29876,N_29725);
nor UO_390 (O_390,N_29779,N_29869);
nand UO_391 (O_391,N_29747,N_29979);
nor UO_392 (O_392,N_29992,N_29813);
nor UO_393 (O_393,N_29811,N_29880);
and UO_394 (O_394,N_29910,N_29901);
or UO_395 (O_395,N_29740,N_29916);
and UO_396 (O_396,N_29749,N_29968);
or UO_397 (O_397,N_29759,N_29885);
or UO_398 (O_398,N_29956,N_29798);
nor UO_399 (O_399,N_29919,N_29871);
nor UO_400 (O_400,N_29941,N_29805);
nand UO_401 (O_401,N_29917,N_29719);
nor UO_402 (O_402,N_29853,N_29710);
and UO_403 (O_403,N_29886,N_29817);
and UO_404 (O_404,N_29870,N_29947);
nand UO_405 (O_405,N_29831,N_29956);
nor UO_406 (O_406,N_29791,N_29711);
xor UO_407 (O_407,N_29966,N_29775);
nand UO_408 (O_408,N_29873,N_29816);
and UO_409 (O_409,N_29817,N_29706);
or UO_410 (O_410,N_29792,N_29831);
xnor UO_411 (O_411,N_29779,N_29912);
xor UO_412 (O_412,N_29712,N_29896);
xor UO_413 (O_413,N_29884,N_29914);
nor UO_414 (O_414,N_29791,N_29710);
xor UO_415 (O_415,N_29873,N_29875);
and UO_416 (O_416,N_29858,N_29941);
xnor UO_417 (O_417,N_29825,N_29723);
xnor UO_418 (O_418,N_29807,N_29849);
xor UO_419 (O_419,N_29711,N_29734);
xor UO_420 (O_420,N_29826,N_29779);
nor UO_421 (O_421,N_29720,N_29796);
nor UO_422 (O_422,N_29771,N_29916);
or UO_423 (O_423,N_29785,N_29950);
nand UO_424 (O_424,N_29783,N_29924);
nor UO_425 (O_425,N_29899,N_29808);
or UO_426 (O_426,N_29859,N_29865);
or UO_427 (O_427,N_29841,N_29934);
nand UO_428 (O_428,N_29801,N_29735);
or UO_429 (O_429,N_29962,N_29791);
nor UO_430 (O_430,N_29895,N_29975);
and UO_431 (O_431,N_29867,N_29786);
xnor UO_432 (O_432,N_29956,N_29915);
nand UO_433 (O_433,N_29780,N_29883);
xnor UO_434 (O_434,N_29830,N_29810);
nand UO_435 (O_435,N_29722,N_29737);
xnor UO_436 (O_436,N_29804,N_29798);
or UO_437 (O_437,N_29940,N_29757);
xnor UO_438 (O_438,N_29960,N_29812);
nor UO_439 (O_439,N_29728,N_29751);
xor UO_440 (O_440,N_29990,N_29762);
xnor UO_441 (O_441,N_29949,N_29990);
and UO_442 (O_442,N_29706,N_29875);
and UO_443 (O_443,N_29738,N_29987);
or UO_444 (O_444,N_29724,N_29834);
and UO_445 (O_445,N_29771,N_29971);
xnor UO_446 (O_446,N_29770,N_29959);
nand UO_447 (O_447,N_29925,N_29876);
nand UO_448 (O_448,N_29885,N_29979);
xor UO_449 (O_449,N_29856,N_29988);
nand UO_450 (O_450,N_29971,N_29723);
nand UO_451 (O_451,N_29885,N_29949);
or UO_452 (O_452,N_29986,N_29934);
nor UO_453 (O_453,N_29877,N_29934);
and UO_454 (O_454,N_29880,N_29787);
nand UO_455 (O_455,N_29903,N_29923);
and UO_456 (O_456,N_29781,N_29959);
or UO_457 (O_457,N_29793,N_29806);
and UO_458 (O_458,N_29716,N_29899);
nand UO_459 (O_459,N_29848,N_29814);
nand UO_460 (O_460,N_29933,N_29884);
xnor UO_461 (O_461,N_29831,N_29802);
nand UO_462 (O_462,N_29907,N_29870);
or UO_463 (O_463,N_29729,N_29998);
nor UO_464 (O_464,N_29817,N_29958);
and UO_465 (O_465,N_29954,N_29765);
nand UO_466 (O_466,N_29924,N_29900);
and UO_467 (O_467,N_29837,N_29700);
nand UO_468 (O_468,N_29716,N_29717);
nor UO_469 (O_469,N_29857,N_29741);
nand UO_470 (O_470,N_29739,N_29971);
and UO_471 (O_471,N_29917,N_29918);
nand UO_472 (O_472,N_29744,N_29804);
and UO_473 (O_473,N_29772,N_29999);
xnor UO_474 (O_474,N_29917,N_29973);
nor UO_475 (O_475,N_29901,N_29774);
or UO_476 (O_476,N_29952,N_29883);
and UO_477 (O_477,N_29890,N_29764);
nor UO_478 (O_478,N_29935,N_29876);
or UO_479 (O_479,N_29822,N_29914);
nand UO_480 (O_480,N_29900,N_29785);
nand UO_481 (O_481,N_29801,N_29922);
xor UO_482 (O_482,N_29869,N_29916);
and UO_483 (O_483,N_29968,N_29841);
and UO_484 (O_484,N_29776,N_29849);
or UO_485 (O_485,N_29768,N_29936);
or UO_486 (O_486,N_29780,N_29972);
or UO_487 (O_487,N_29809,N_29837);
nand UO_488 (O_488,N_29718,N_29858);
nor UO_489 (O_489,N_29703,N_29769);
nand UO_490 (O_490,N_29925,N_29729);
nor UO_491 (O_491,N_29869,N_29757);
and UO_492 (O_492,N_29888,N_29974);
or UO_493 (O_493,N_29709,N_29868);
nand UO_494 (O_494,N_29822,N_29998);
nand UO_495 (O_495,N_29762,N_29720);
or UO_496 (O_496,N_29976,N_29757);
or UO_497 (O_497,N_29748,N_29753);
xnor UO_498 (O_498,N_29969,N_29802);
or UO_499 (O_499,N_29768,N_29974);
and UO_500 (O_500,N_29981,N_29730);
nor UO_501 (O_501,N_29909,N_29760);
or UO_502 (O_502,N_29791,N_29809);
nor UO_503 (O_503,N_29980,N_29925);
or UO_504 (O_504,N_29784,N_29764);
and UO_505 (O_505,N_29817,N_29722);
nor UO_506 (O_506,N_29987,N_29759);
or UO_507 (O_507,N_29725,N_29957);
nor UO_508 (O_508,N_29924,N_29748);
xor UO_509 (O_509,N_29769,N_29927);
xor UO_510 (O_510,N_29749,N_29978);
and UO_511 (O_511,N_29988,N_29768);
and UO_512 (O_512,N_29929,N_29722);
nand UO_513 (O_513,N_29930,N_29781);
nor UO_514 (O_514,N_29771,N_29841);
xnor UO_515 (O_515,N_29749,N_29865);
nand UO_516 (O_516,N_29758,N_29957);
and UO_517 (O_517,N_29777,N_29765);
and UO_518 (O_518,N_29778,N_29892);
or UO_519 (O_519,N_29743,N_29737);
xor UO_520 (O_520,N_29878,N_29827);
nor UO_521 (O_521,N_29712,N_29773);
xor UO_522 (O_522,N_29848,N_29884);
nand UO_523 (O_523,N_29805,N_29893);
nor UO_524 (O_524,N_29974,N_29837);
nand UO_525 (O_525,N_29876,N_29948);
nand UO_526 (O_526,N_29890,N_29802);
nand UO_527 (O_527,N_29952,N_29734);
nor UO_528 (O_528,N_29889,N_29747);
and UO_529 (O_529,N_29813,N_29980);
nor UO_530 (O_530,N_29782,N_29933);
or UO_531 (O_531,N_29874,N_29778);
and UO_532 (O_532,N_29784,N_29797);
xnor UO_533 (O_533,N_29821,N_29994);
and UO_534 (O_534,N_29854,N_29887);
nand UO_535 (O_535,N_29874,N_29918);
nand UO_536 (O_536,N_29841,N_29774);
nand UO_537 (O_537,N_29866,N_29768);
and UO_538 (O_538,N_29700,N_29775);
xnor UO_539 (O_539,N_29916,N_29986);
xnor UO_540 (O_540,N_29903,N_29830);
nor UO_541 (O_541,N_29937,N_29846);
nor UO_542 (O_542,N_29748,N_29716);
xor UO_543 (O_543,N_29726,N_29976);
nor UO_544 (O_544,N_29780,N_29821);
xor UO_545 (O_545,N_29730,N_29928);
or UO_546 (O_546,N_29764,N_29957);
and UO_547 (O_547,N_29813,N_29826);
xnor UO_548 (O_548,N_29769,N_29809);
or UO_549 (O_549,N_29774,N_29793);
or UO_550 (O_550,N_29904,N_29937);
xor UO_551 (O_551,N_29942,N_29947);
or UO_552 (O_552,N_29719,N_29922);
or UO_553 (O_553,N_29858,N_29927);
nor UO_554 (O_554,N_29764,N_29999);
nand UO_555 (O_555,N_29848,N_29762);
xor UO_556 (O_556,N_29864,N_29803);
or UO_557 (O_557,N_29890,N_29817);
and UO_558 (O_558,N_29989,N_29972);
or UO_559 (O_559,N_29801,N_29854);
nand UO_560 (O_560,N_29934,N_29987);
xor UO_561 (O_561,N_29940,N_29974);
or UO_562 (O_562,N_29845,N_29917);
and UO_563 (O_563,N_29997,N_29768);
nand UO_564 (O_564,N_29763,N_29820);
and UO_565 (O_565,N_29894,N_29845);
nor UO_566 (O_566,N_29841,N_29756);
xnor UO_567 (O_567,N_29821,N_29729);
or UO_568 (O_568,N_29839,N_29857);
and UO_569 (O_569,N_29980,N_29836);
xnor UO_570 (O_570,N_29745,N_29828);
or UO_571 (O_571,N_29784,N_29750);
nor UO_572 (O_572,N_29915,N_29707);
xnor UO_573 (O_573,N_29952,N_29913);
nor UO_574 (O_574,N_29897,N_29845);
nor UO_575 (O_575,N_29853,N_29871);
or UO_576 (O_576,N_29867,N_29951);
and UO_577 (O_577,N_29746,N_29908);
and UO_578 (O_578,N_29924,N_29797);
nor UO_579 (O_579,N_29875,N_29701);
nand UO_580 (O_580,N_29835,N_29853);
or UO_581 (O_581,N_29767,N_29721);
nor UO_582 (O_582,N_29765,N_29701);
nand UO_583 (O_583,N_29796,N_29819);
nand UO_584 (O_584,N_29979,N_29751);
or UO_585 (O_585,N_29705,N_29876);
nand UO_586 (O_586,N_29720,N_29869);
or UO_587 (O_587,N_29938,N_29928);
nand UO_588 (O_588,N_29941,N_29890);
or UO_589 (O_589,N_29921,N_29718);
or UO_590 (O_590,N_29730,N_29719);
nor UO_591 (O_591,N_29891,N_29777);
nand UO_592 (O_592,N_29778,N_29891);
nor UO_593 (O_593,N_29941,N_29916);
xnor UO_594 (O_594,N_29741,N_29824);
or UO_595 (O_595,N_29883,N_29758);
nand UO_596 (O_596,N_29728,N_29950);
or UO_597 (O_597,N_29887,N_29893);
and UO_598 (O_598,N_29984,N_29885);
or UO_599 (O_599,N_29734,N_29866);
and UO_600 (O_600,N_29835,N_29900);
nand UO_601 (O_601,N_29807,N_29873);
or UO_602 (O_602,N_29849,N_29894);
and UO_603 (O_603,N_29782,N_29706);
nor UO_604 (O_604,N_29765,N_29950);
or UO_605 (O_605,N_29828,N_29916);
and UO_606 (O_606,N_29717,N_29903);
or UO_607 (O_607,N_29865,N_29824);
nor UO_608 (O_608,N_29884,N_29954);
xor UO_609 (O_609,N_29916,N_29775);
nor UO_610 (O_610,N_29902,N_29844);
nor UO_611 (O_611,N_29823,N_29926);
nor UO_612 (O_612,N_29718,N_29739);
nor UO_613 (O_613,N_29957,N_29920);
nor UO_614 (O_614,N_29963,N_29964);
and UO_615 (O_615,N_29897,N_29758);
nand UO_616 (O_616,N_29799,N_29735);
or UO_617 (O_617,N_29917,N_29741);
xnor UO_618 (O_618,N_29913,N_29702);
and UO_619 (O_619,N_29993,N_29716);
xor UO_620 (O_620,N_29917,N_29711);
nor UO_621 (O_621,N_29885,N_29742);
and UO_622 (O_622,N_29741,N_29919);
xor UO_623 (O_623,N_29873,N_29717);
xor UO_624 (O_624,N_29967,N_29838);
and UO_625 (O_625,N_29992,N_29834);
nor UO_626 (O_626,N_29715,N_29765);
xnor UO_627 (O_627,N_29738,N_29790);
nand UO_628 (O_628,N_29714,N_29887);
nor UO_629 (O_629,N_29858,N_29717);
xor UO_630 (O_630,N_29785,N_29844);
xnor UO_631 (O_631,N_29790,N_29903);
or UO_632 (O_632,N_29732,N_29769);
xor UO_633 (O_633,N_29907,N_29822);
or UO_634 (O_634,N_29931,N_29955);
nor UO_635 (O_635,N_29813,N_29961);
xnor UO_636 (O_636,N_29893,N_29734);
nand UO_637 (O_637,N_29813,N_29878);
and UO_638 (O_638,N_29850,N_29856);
nand UO_639 (O_639,N_29958,N_29832);
or UO_640 (O_640,N_29874,N_29996);
or UO_641 (O_641,N_29710,N_29938);
nand UO_642 (O_642,N_29794,N_29929);
xor UO_643 (O_643,N_29829,N_29814);
nand UO_644 (O_644,N_29995,N_29824);
and UO_645 (O_645,N_29878,N_29730);
nand UO_646 (O_646,N_29768,N_29762);
nand UO_647 (O_647,N_29770,N_29717);
and UO_648 (O_648,N_29892,N_29752);
nor UO_649 (O_649,N_29885,N_29856);
or UO_650 (O_650,N_29841,N_29883);
xor UO_651 (O_651,N_29859,N_29982);
nor UO_652 (O_652,N_29806,N_29893);
and UO_653 (O_653,N_29935,N_29999);
nor UO_654 (O_654,N_29978,N_29777);
nor UO_655 (O_655,N_29756,N_29824);
nand UO_656 (O_656,N_29843,N_29881);
nor UO_657 (O_657,N_29900,N_29858);
nor UO_658 (O_658,N_29965,N_29780);
and UO_659 (O_659,N_29986,N_29765);
xnor UO_660 (O_660,N_29762,N_29718);
nor UO_661 (O_661,N_29741,N_29851);
nand UO_662 (O_662,N_29728,N_29980);
nor UO_663 (O_663,N_29801,N_29894);
or UO_664 (O_664,N_29777,N_29798);
xor UO_665 (O_665,N_29744,N_29956);
and UO_666 (O_666,N_29703,N_29756);
or UO_667 (O_667,N_29979,N_29965);
nor UO_668 (O_668,N_29831,N_29945);
nor UO_669 (O_669,N_29900,N_29897);
nand UO_670 (O_670,N_29932,N_29899);
xnor UO_671 (O_671,N_29960,N_29867);
and UO_672 (O_672,N_29898,N_29704);
and UO_673 (O_673,N_29867,N_29875);
xor UO_674 (O_674,N_29958,N_29800);
nor UO_675 (O_675,N_29725,N_29920);
or UO_676 (O_676,N_29955,N_29957);
nand UO_677 (O_677,N_29868,N_29720);
xor UO_678 (O_678,N_29808,N_29831);
nand UO_679 (O_679,N_29852,N_29914);
xor UO_680 (O_680,N_29929,N_29726);
nor UO_681 (O_681,N_29787,N_29902);
and UO_682 (O_682,N_29734,N_29821);
nor UO_683 (O_683,N_29935,N_29952);
and UO_684 (O_684,N_29991,N_29898);
xnor UO_685 (O_685,N_29707,N_29925);
and UO_686 (O_686,N_29805,N_29879);
and UO_687 (O_687,N_29744,N_29896);
or UO_688 (O_688,N_29880,N_29756);
nor UO_689 (O_689,N_29999,N_29784);
nand UO_690 (O_690,N_29883,N_29808);
xor UO_691 (O_691,N_29789,N_29772);
and UO_692 (O_692,N_29944,N_29976);
nor UO_693 (O_693,N_29796,N_29704);
nor UO_694 (O_694,N_29736,N_29883);
or UO_695 (O_695,N_29972,N_29875);
nand UO_696 (O_696,N_29840,N_29855);
or UO_697 (O_697,N_29727,N_29960);
nor UO_698 (O_698,N_29763,N_29919);
or UO_699 (O_699,N_29950,N_29775);
nand UO_700 (O_700,N_29809,N_29710);
xnor UO_701 (O_701,N_29783,N_29934);
xor UO_702 (O_702,N_29817,N_29742);
nor UO_703 (O_703,N_29862,N_29953);
nor UO_704 (O_704,N_29726,N_29872);
nand UO_705 (O_705,N_29711,N_29901);
nand UO_706 (O_706,N_29737,N_29922);
xor UO_707 (O_707,N_29862,N_29708);
and UO_708 (O_708,N_29750,N_29830);
xor UO_709 (O_709,N_29769,N_29902);
nor UO_710 (O_710,N_29899,N_29827);
or UO_711 (O_711,N_29964,N_29928);
nor UO_712 (O_712,N_29945,N_29936);
and UO_713 (O_713,N_29881,N_29787);
or UO_714 (O_714,N_29998,N_29804);
nor UO_715 (O_715,N_29791,N_29764);
nor UO_716 (O_716,N_29837,N_29954);
xor UO_717 (O_717,N_29701,N_29929);
and UO_718 (O_718,N_29877,N_29993);
nor UO_719 (O_719,N_29992,N_29863);
nor UO_720 (O_720,N_29802,N_29767);
nor UO_721 (O_721,N_29932,N_29723);
or UO_722 (O_722,N_29863,N_29971);
xnor UO_723 (O_723,N_29908,N_29929);
nand UO_724 (O_724,N_29909,N_29858);
or UO_725 (O_725,N_29992,N_29848);
and UO_726 (O_726,N_29750,N_29884);
xnor UO_727 (O_727,N_29954,N_29921);
or UO_728 (O_728,N_29831,N_29729);
and UO_729 (O_729,N_29790,N_29731);
nor UO_730 (O_730,N_29831,N_29852);
xor UO_731 (O_731,N_29866,N_29716);
or UO_732 (O_732,N_29949,N_29725);
and UO_733 (O_733,N_29991,N_29904);
or UO_734 (O_734,N_29776,N_29834);
xnor UO_735 (O_735,N_29892,N_29887);
xor UO_736 (O_736,N_29880,N_29805);
xnor UO_737 (O_737,N_29863,N_29905);
xnor UO_738 (O_738,N_29954,N_29818);
xnor UO_739 (O_739,N_29800,N_29916);
or UO_740 (O_740,N_29974,N_29781);
or UO_741 (O_741,N_29792,N_29788);
and UO_742 (O_742,N_29865,N_29732);
xnor UO_743 (O_743,N_29934,N_29784);
nand UO_744 (O_744,N_29964,N_29706);
xor UO_745 (O_745,N_29889,N_29725);
and UO_746 (O_746,N_29958,N_29815);
and UO_747 (O_747,N_29856,N_29906);
and UO_748 (O_748,N_29702,N_29753);
or UO_749 (O_749,N_29958,N_29730);
nor UO_750 (O_750,N_29989,N_29859);
nand UO_751 (O_751,N_29840,N_29906);
nand UO_752 (O_752,N_29968,N_29865);
and UO_753 (O_753,N_29947,N_29726);
nand UO_754 (O_754,N_29817,N_29915);
xor UO_755 (O_755,N_29987,N_29856);
or UO_756 (O_756,N_29763,N_29968);
or UO_757 (O_757,N_29968,N_29813);
nor UO_758 (O_758,N_29901,N_29725);
nor UO_759 (O_759,N_29967,N_29738);
xnor UO_760 (O_760,N_29990,N_29701);
xor UO_761 (O_761,N_29909,N_29774);
nand UO_762 (O_762,N_29743,N_29969);
and UO_763 (O_763,N_29830,N_29717);
xor UO_764 (O_764,N_29853,N_29928);
xnor UO_765 (O_765,N_29949,N_29800);
nor UO_766 (O_766,N_29970,N_29945);
or UO_767 (O_767,N_29804,N_29870);
nor UO_768 (O_768,N_29927,N_29736);
nor UO_769 (O_769,N_29979,N_29841);
xnor UO_770 (O_770,N_29728,N_29739);
nand UO_771 (O_771,N_29702,N_29889);
or UO_772 (O_772,N_29829,N_29965);
xnor UO_773 (O_773,N_29993,N_29830);
or UO_774 (O_774,N_29797,N_29744);
nand UO_775 (O_775,N_29719,N_29995);
nor UO_776 (O_776,N_29830,N_29867);
or UO_777 (O_777,N_29963,N_29745);
nor UO_778 (O_778,N_29746,N_29727);
nand UO_779 (O_779,N_29746,N_29843);
nand UO_780 (O_780,N_29899,N_29809);
nand UO_781 (O_781,N_29752,N_29706);
or UO_782 (O_782,N_29892,N_29890);
nor UO_783 (O_783,N_29831,N_29997);
or UO_784 (O_784,N_29958,N_29752);
nor UO_785 (O_785,N_29964,N_29708);
and UO_786 (O_786,N_29953,N_29873);
and UO_787 (O_787,N_29709,N_29825);
and UO_788 (O_788,N_29962,N_29970);
nand UO_789 (O_789,N_29834,N_29840);
and UO_790 (O_790,N_29950,N_29936);
and UO_791 (O_791,N_29927,N_29850);
nor UO_792 (O_792,N_29997,N_29917);
and UO_793 (O_793,N_29729,N_29949);
or UO_794 (O_794,N_29965,N_29926);
nand UO_795 (O_795,N_29780,N_29753);
xor UO_796 (O_796,N_29788,N_29703);
or UO_797 (O_797,N_29987,N_29750);
and UO_798 (O_798,N_29852,N_29896);
and UO_799 (O_799,N_29804,N_29838);
and UO_800 (O_800,N_29985,N_29707);
nand UO_801 (O_801,N_29784,N_29759);
and UO_802 (O_802,N_29987,N_29926);
and UO_803 (O_803,N_29847,N_29888);
xor UO_804 (O_804,N_29886,N_29827);
nor UO_805 (O_805,N_29939,N_29830);
xor UO_806 (O_806,N_29752,N_29709);
xnor UO_807 (O_807,N_29865,N_29947);
xor UO_808 (O_808,N_29752,N_29972);
xor UO_809 (O_809,N_29790,N_29964);
nor UO_810 (O_810,N_29749,N_29818);
and UO_811 (O_811,N_29760,N_29798);
and UO_812 (O_812,N_29794,N_29767);
xnor UO_813 (O_813,N_29727,N_29745);
nor UO_814 (O_814,N_29926,N_29711);
xnor UO_815 (O_815,N_29759,N_29875);
or UO_816 (O_816,N_29956,N_29778);
or UO_817 (O_817,N_29980,N_29945);
nor UO_818 (O_818,N_29848,N_29878);
or UO_819 (O_819,N_29976,N_29706);
nand UO_820 (O_820,N_29977,N_29888);
xor UO_821 (O_821,N_29953,N_29872);
xnor UO_822 (O_822,N_29912,N_29716);
and UO_823 (O_823,N_29858,N_29852);
nand UO_824 (O_824,N_29864,N_29908);
nand UO_825 (O_825,N_29949,N_29749);
xnor UO_826 (O_826,N_29726,N_29709);
xor UO_827 (O_827,N_29877,N_29784);
or UO_828 (O_828,N_29957,N_29927);
and UO_829 (O_829,N_29782,N_29946);
or UO_830 (O_830,N_29790,N_29784);
nor UO_831 (O_831,N_29967,N_29998);
and UO_832 (O_832,N_29807,N_29718);
xor UO_833 (O_833,N_29702,N_29709);
nand UO_834 (O_834,N_29842,N_29787);
and UO_835 (O_835,N_29851,N_29962);
nor UO_836 (O_836,N_29743,N_29859);
and UO_837 (O_837,N_29959,N_29754);
xor UO_838 (O_838,N_29908,N_29801);
or UO_839 (O_839,N_29717,N_29992);
nand UO_840 (O_840,N_29974,N_29894);
nand UO_841 (O_841,N_29713,N_29808);
xor UO_842 (O_842,N_29976,N_29940);
xor UO_843 (O_843,N_29741,N_29784);
nand UO_844 (O_844,N_29996,N_29892);
nand UO_845 (O_845,N_29912,N_29944);
nor UO_846 (O_846,N_29907,N_29933);
and UO_847 (O_847,N_29826,N_29746);
and UO_848 (O_848,N_29827,N_29888);
nor UO_849 (O_849,N_29771,N_29847);
nor UO_850 (O_850,N_29891,N_29887);
nand UO_851 (O_851,N_29971,N_29872);
xor UO_852 (O_852,N_29882,N_29887);
nand UO_853 (O_853,N_29807,N_29886);
nand UO_854 (O_854,N_29890,N_29827);
and UO_855 (O_855,N_29929,N_29876);
xor UO_856 (O_856,N_29898,N_29993);
or UO_857 (O_857,N_29810,N_29994);
nor UO_858 (O_858,N_29784,N_29899);
nor UO_859 (O_859,N_29817,N_29832);
and UO_860 (O_860,N_29761,N_29837);
nand UO_861 (O_861,N_29780,N_29824);
or UO_862 (O_862,N_29977,N_29803);
and UO_863 (O_863,N_29711,N_29841);
or UO_864 (O_864,N_29896,N_29834);
nor UO_865 (O_865,N_29748,N_29742);
and UO_866 (O_866,N_29834,N_29756);
nor UO_867 (O_867,N_29710,N_29937);
and UO_868 (O_868,N_29924,N_29716);
and UO_869 (O_869,N_29850,N_29928);
nand UO_870 (O_870,N_29882,N_29791);
or UO_871 (O_871,N_29865,N_29860);
xnor UO_872 (O_872,N_29709,N_29927);
xnor UO_873 (O_873,N_29700,N_29740);
or UO_874 (O_874,N_29790,N_29855);
xor UO_875 (O_875,N_29811,N_29799);
nor UO_876 (O_876,N_29875,N_29981);
nor UO_877 (O_877,N_29849,N_29785);
nor UO_878 (O_878,N_29887,N_29777);
xor UO_879 (O_879,N_29794,N_29916);
nand UO_880 (O_880,N_29912,N_29840);
and UO_881 (O_881,N_29890,N_29762);
xor UO_882 (O_882,N_29776,N_29739);
and UO_883 (O_883,N_29766,N_29792);
nor UO_884 (O_884,N_29799,N_29909);
xor UO_885 (O_885,N_29711,N_29784);
and UO_886 (O_886,N_29751,N_29756);
or UO_887 (O_887,N_29988,N_29747);
nor UO_888 (O_888,N_29890,N_29889);
or UO_889 (O_889,N_29875,N_29885);
and UO_890 (O_890,N_29990,N_29856);
and UO_891 (O_891,N_29754,N_29952);
nand UO_892 (O_892,N_29737,N_29823);
or UO_893 (O_893,N_29932,N_29801);
or UO_894 (O_894,N_29849,N_29715);
nand UO_895 (O_895,N_29915,N_29889);
xnor UO_896 (O_896,N_29815,N_29719);
nor UO_897 (O_897,N_29959,N_29724);
or UO_898 (O_898,N_29779,N_29839);
or UO_899 (O_899,N_29992,N_29732);
nor UO_900 (O_900,N_29898,N_29837);
or UO_901 (O_901,N_29777,N_29785);
nand UO_902 (O_902,N_29918,N_29755);
nand UO_903 (O_903,N_29871,N_29762);
and UO_904 (O_904,N_29905,N_29807);
or UO_905 (O_905,N_29948,N_29934);
or UO_906 (O_906,N_29973,N_29796);
nor UO_907 (O_907,N_29927,N_29979);
and UO_908 (O_908,N_29758,N_29874);
nor UO_909 (O_909,N_29872,N_29938);
nor UO_910 (O_910,N_29936,N_29820);
xnor UO_911 (O_911,N_29856,N_29881);
nor UO_912 (O_912,N_29910,N_29764);
or UO_913 (O_913,N_29930,N_29952);
or UO_914 (O_914,N_29925,N_29741);
xnor UO_915 (O_915,N_29954,N_29860);
nand UO_916 (O_916,N_29708,N_29879);
nand UO_917 (O_917,N_29865,N_29925);
nand UO_918 (O_918,N_29960,N_29719);
and UO_919 (O_919,N_29754,N_29811);
and UO_920 (O_920,N_29774,N_29859);
or UO_921 (O_921,N_29992,N_29786);
nor UO_922 (O_922,N_29848,N_29998);
nand UO_923 (O_923,N_29706,N_29912);
or UO_924 (O_924,N_29845,N_29891);
nor UO_925 (O_925,N_29897,N_29807);
nand UO_926 (O_926,N_29752,N_29700);
nand UO_927 (O_927,N_29910,N_29754);
or UO_928 (O_928,N_29789,N_29955);
and UO_929 (O_929,N_29895,N_29793);
xnor UO_930 (O_930,N_29823,N_29898);
and UO_931 (O_931,N_29933,N_29812);
xor UO_932 (O_932,N_29963,N_29744);
or UO_933 (O_933,N_29871,N_29953);
or UO_934 (O_934,N_29812,N_29899);
or UO_935 (O_935,N_29705,N_29748);
and UO_936 (O_936,N_29784,N_29846);
nand UO_937 (O_937,N_29765,N_29970);
and UO_938 (O_938,N_29728,N_29771);
nand UO_939 (O_939,N_29778,N_29905);
nor UO_940 (O_940,N_29927,N_29800);
nor UO_941 (O_941,N_29912,N_29838);
or UO_942 (O_942,N_29887,N_29982);
nor UO_943 (O_943,N_29909,N_29874);
and UO_944 (O_944,N_29851,N_29749);
xnor UO_945 (O_945,N_29757,N_29917);
and UO_946 (O_946,N_29923,N_29761);
and UO_947 (O_947,N_29758,N_29956);
and UO_948 (O_948,N_29938,N_29825);
nand UO_949 (O_949,N_29825,N_29718);
xnor UO_950 (O_950,N_29947,N_29802);
nor UO_951 (O_951,N_29965,N_29752);
nor UO_952 (O_952,N_29892,N_29708);
nand UO_953 (O_953,N_29938,N_29766);
xor UO_954 (O_954,N_29796,N_29837);
xnor UO_955 (O_955,N_29853,N_29976);
nor UO_956 (O_956,N_29774,N_29883);
nor UO_957 (O_957,N_29898,N_29975);
xor UO_958 (O_958,N_29803,N_29805);
xor UO_959 (O_959,N_29778,N_29909);
nand UO_960 (O_960,N_29942,N_29741);
nand UO_961 (O_961,N_29892,N_29702);
and UO_962 (O_962,N_29836,N_29753);
nand UO_963 (O_963,N_29764,N_29962);
nor UO_964 (O_964,N_29856,N_29763);
or UO_965 (O_965,N_29938,N_29822);
xnor UO_966 (O_966,N_29800,N_29806);
or UO_967 (O_967,N_29823,N_29760);
nor UO_968 (O_968,N_29796,N_29897);
xnor UO_969 (O_969,N_29829,N_29768);
nor UO_970 (O_970,N_29912,N_29834);
xor UO_971 (O_971,N_29970,N_29728);
nor UO_972 (O_972,N_29886,N_29889);
and UO_973 (O_973,N_29700,N_29954);
nor UO_974 (O_974,N_29842,N_29789);
or UO_975 (O_975,N_29950,N_29934);
xnor UO_976 (O_976,N_29751,N_29735);
xor UO_977 (O_977,N_29781,N_29829);
nor UO_978 (O_978,N_29811,N_29746);
xnor UO_979 (O_979,N_29731,N_29827);
xnor UO_980 (O_980,N_29977,N_29784);
nand UO_981 (O_981,N_29878,N_29984);
xnor UO_982 (O_982,N_29750,N_29747);
xnor UO_983 (O_983,N_29900,N_29973);
or UO_984 (O_984,N_29836,N_29756);
xor UO_985 (O_985,N_29737,N_29827);
and UO_986 (O_986,N_29771,N_29938);
and UO_987 (O_987,N_29715,N_29863);
nand UO_988 (O_988,N_29831,N_29898);
nand UO_989 (O_989,N_29895,N_29875);
and UO_990 (O_990,N_29817,N_29922);
or UO_991 (O_991,N_29751,N_29982);
xor UO_992 (O_992,N_29701,N_29986);
nor UO_993 (O_993,N_29706,N_29899);
and UO_994 (O_994,N_29944,N_29784);
or UO_995 (O_995,N_29777,N_29717);
and UO_996 (O_996,N_29860,N_29711);
xnor UO_997 (O_997,N_29892,N_29850);
or UO_998 (O_998,N_29709,N_29881);
nor UO_999 (O_999,N_29970,N_29906);
and UO_1000 (O_1000,N_29993,N_29730);
and UO_1001 (O_1001,N_29878,N_29883);
xor UO_1002 (O_1002,N_29771,N_29866);
nor UO_1003 (O_1003,N_29947,N_29789);
xnor UO_1004 (O_1004,N_29938,N_29877);
or UO_1005 (O_1005,N_29885,N_29804);
or UO_1006 (O_1006,N_29766,N_29789);
and UO_1007 (O_1007,N_29759,N_29919);
or UO_1008 (O_1008,N_29773,N_29847);
and UO_1009 (O_1009,N_29978,N_29944);
and UO_1010 (O_1010,N_29781,N_29991);
or UO_1011 (O_1011,N_29783,N_29762);
xnor UO_1012 (O_1012,N_29732,N_29960);
xor UO_1013 (O_1013,N_29928,N_29818);
or UO_1014 (O_1014,N_29792,N_29990);
xnor UO_1015 (O_1015,N_29908,N_29803);
or UO_1016 (O_1016,N_29928,N_29722);
nor UO_1017 (O_1017,N_29749,N_29727);
nand UO_1018 (O_1018,N_29815,N_29807);
and UO_1019 (O_1019,N_29728,N_29883);
xor UO_1020 (O_1020,N_29964,N_29893);
nand UO_1021 (O_1021,N_29832,N_29703);
nor UO_1022 (O_1022,N_29799,N_29796);
nor UO_1023 (O_1023,N_29976,N_29785);
or UO_1024 (O_1024,N_29816,N_29894);
and UO_1025 (O_1025,N_29793,N_29771);
xor UO_1026 (O_1026,N_29893,N_29986);
and UO_1027 (O_1027,N_29956,N_29857);
and UO_1028 (O_1028,N_29779,N_29961);
nor UO_1029 (O_1029,N_29859,N_29778);
nor UO_1030 (O_1030,N_29855,N_29764);
xnor UO_1031 (O_1031,N_29743,N_29890);
nand UO_1032 (O_1032,N_29703,N_29911);
nand UO_1033 (O_1033,N_29779,N_29823);
nand UO_1034 (O_1034,N_29894,N_29977);
and UO_1035 (O_1035,N_29718,N_29787);
or UO_1036 (O_1036,N_29778,N_29735);
nor UO_1037 (O_1037,N_29809,N_29740);
xor UO_1038 (O_1038,N_29906,N_29866);
and UO_1039 (O_1039,N_29804,N_29994);
xor UO_1040 (O_1040,N_29966,N_29919);
and UO_1041 (O_1041,N_29860,N_29745);
nand UO_1042 (O_1042,N_29849,N_29708);
xnor UO_1043 (O_1043,N_29945,N_29973);
or UO_1044 (O_1044,N_29893,N_29995);
and UO_1045 (O_1045,N_29987,N_29932);
and UO_1046 (O_1046,N_29853,N_29940);
nor UO_1047 (O_1047,N_29788,N_29784);
nor UO_1048 (O_1048,N_29930,N_29895);
xnor UO_1049 (O_1049,N_29811,N_29998);
xnor UO_1050 (O_1050,N_29922,N_29755);
xor UO_1051 (O_1051,N_29914,N_29973);
or UO_1052 (O_1052,N_29830,N_29756);
or UO_1053 (O_1053,N_29832,N_29775);
or UO_1054 (O_1054,N_29940,N_29900);
nand UO_1055 (O_1055,N_29818,N_29967);
and UO_1056 (O_1056,N_29718,N_29841);
nand UO_1057 (O_1057,N_29950,N_29973);
and UO_1058 (O_1058,N_29747,N_29795);
xnor UO_1059 (O_1059,N_29870,N_29837);
xnor UO_1060 (O_1060,N_29707,N_29880);
nand UO_1061 (O_1061,N_29823,N_29701);
and UO_1062 (O_1062,N_29923,N_29947);
xor UO_1063 (O_1063,N_29714,N_29773);
and UO_1064 (O_1064,N_29989,N_29749);
nand UO_1065 (O_1065,N_29775,N_29933);
xor UO_1066 (O_1066,N_29967,N_29861);
nand UO_1067 (O_1067,N_29982,N_29849);
and UO_1068 (O_1068,N_29947,N_29937);
and UO_1069 (O_1069,N_29814,N_29936);
xnor UO_1070 (O_1070,N_29838,N_29908);
nand UO_1071 (O_1071,N_29744,N_29860);
xor UO_1072 (O_1072,N_29955,N_29915);
nor UO_1073 (O_1073,N_29958,N_29795);
nor UO_1074 (O_1074,N_29966,N_29710);
and UO_1075 (O_1075,N_29809,N_29828);
and UO_1076 (O_1076,N_29777,N_29903);
nor UO_1077 (O_1077,N_29845,N_29938);
nand UO_1078 (O_1078,N_29820,N_29954);
xor UO_1079 (O_1079,N_29912,N_29713);
or UO_1080 (O_1080,N_29811,N_29702);
and UO_1081 (O_1081,N_29791,N_29736);
or UO_1082 (O_1082,N_29827,N_29847);
and UO_1083 (O_1083,N_29966,N_29848);
nor UO_1084 (O_1084,N_29910,N_29997);
xnor UO_1085 (O_1085,N_29909,N_29906);
nand UO_1086 (O_1086,N_29800,N_29818);
xnor UO_1087 (O_1087,N_29870,N_29973);
nand UO_1088 (O_1088,N_29848,N_29775);
xor UO_1089 (O_1089,N_29808,N_29848);
nand UO_1090 (O_1090,N_29894,N_29762);
or UO_1091 (O_1091,N_29955,N_29800);
and UO_1092 (O_1092,N_29878,N_29823);
or UO_1093 (O_1093,N_29810,N_29834);
or UO_1094 (O_1094,N_29779,N_29865);
xor UO_1095 (O_1095,N_29819,N_29810);
nor UO_1096 (O_1096,N_29932,N_29706);
and UO_1097 (O_1097,N_29767,N_29755);
xor UO_1098 (O_1098,N_29755,N_29730);
nor UO_1099 (O_1099,N_29788,N_29998);
and UO_1100 (O_1100,N_29802,N_29957);
xor UO_1101 (O_1101,N_29960,N_29840);
nor UO_1102 (O_1102,N_29899,N_29880);
nor UO_1103 (O_1103,N_29905,N_29811);
nor UO_1104 (O_1104,N_29909,N_29902);
xnor UO_1105 (O_1105,N_29811,N_29986);
nor UO_1106 (O_1106,N_29969,N_29735);
or UO_1107 (O_1107,N_29924,N_29927);
and UO_1108 (O_1108,N_29889,N_29836);
nand UO_1109 (O_1109,N_29725,N_29732);
xnor UO_1110 (O_1110,N_29853,N_29849);
and UO_1111 (O_1111,N_29744,N_29781);
nor UO_1112 (O_1112,N_29828,N_29869);
nand UO_1113 (O_1113,N_29947,N_29829);
and UO_1114 (O_1114,N_29818,N_29875);
or UO_1115 (O_1115,N_29755,N_29867);
nand UO_1116 (O_1116,N_29911,N_29990);
xor UO_1117 (O_1117,N_29956,N_29998);
nor UO_1118 (O_1118,N_29949,N_29837);
and UO_1119 (O_1119,N_29801,N_29739);
nand UO_1120 (O_1120,N_29884,N_29798);
nand UO_1121 (O_1121,N_29981,N_29729);
nand UO_1122 (O_1122,N_29959,N_29837);
and UO_1123 (O_1123,N_29877,N_29791);
xor UO_1124 (O_1124,N_29818,N_29998);
and UO_1125 (O_1125,N_29851,N_29923);
xor UO_1126 (O_1126,N_29768,N_29864);
xor UO_1127 (O_1127,N_29750,N_29727);
and UO_1128 (O_1128,N_29945,N_29891);
xnor UO_1129 (O_1129,N_29919,N_29862);
and UO_1130 (O_1130,N_29706,N_29797);
and UO_1131 (O_1131,N_29754,N_29940);
and UO_1132 (O_1132,N_29725,N_29982);
nand UO_1133 (O_1133,N_29719,N_29983);
or UO_1134 (O_1134,N_29931,N_29718);
nor UO_1135 (O_1135,N_29710,N_29703);
or UO_1136 (O_1136,N_29991,N_29833);
nand UO_1137 (O_1137,N_29895,N_29963);
xnor UO_1138 (O_1138,N_29997,N_29795);
nand UO_1139 (O_1139,N_29794,N_29730);
or UO_1140 (O_1140,N_29799,N_29971);
nor UO_1141 (O_1141,N_29893,N_29882);
nand UO_1142 (O_1142,N_29911,N_29796);
and UO_1143 (O_1143,N_29789,N_29833);
or UO_1144 (O_1144,N_29842,N_29858);
xor UO_1145 (O_1145,N_29824,N_29787);
nand UO_1146 (O_1146,N_29918,N_29985);
xnor UO_1147 (O_1147,N_29960,N_29927);
xnor UO_1148 (O_1148,N_29996,N_29711);
xor UO_1149 (O_1149,N_29742,N_29760);
xnor UO_1150 (O_1150,N_29938,N_29779);
or UO_1151 (O_1151,N_29876,N_29986);
or UO_1152 (O_1152,N_29938,N_29783);
nand UO_1153 (O_1153,N_29813,N_29766);
nand UO_1154 (O_1154,N_29841,N_29864);
nor UO_1155 (O_1155,N_29929,N_29959);
nor UO_1156 (O_1156,N_29764,N_29763);
nor UO_1157 (O_1157,N_29815,N_29775);
and UO_1158 (O_1158,N_29969,N_29989);
and UO_1159 (O_1159,N_29862,N_29827);
nand UO_1160 (O_1160,N_29939,N_29795);
or UO_1161 (O_1161,N_29845,N_29777);
xor UO_1162 (O_1162,N_29701,N_29989);
nand UO_1163 (O_1163,N_29759,N_29971);
xor UO_1164 (O_1164,N_29877,N_29896);
and UO_1165 (O_1165,N_29935,N_29833);
nand UO_1166 (O_1166,N_29961,N_29919);
nand UO_1167 (O_1167,N_29891,N_29763);
or UO_1168 (O_1168,N_29744,N_29768);
and UO_1169 (O_1169,N_29711,N_29842);
and UO_1170 (O_1170,N_29807,N_29800);
or UO_1171 (O_1171,N_29846,N_29813);
nand UO_1172 (O_1172,N_29908,N_29783);
and UO_1173 (O_1173,N_29772,N_29978);
and UO_1174 (O_1174,N_29867,N_29859);
nor UO_1175 (O_1175,N_29942,N_29833);
and UO_1176 (O_1176,N_29706,N_29930);
nor UO_1177 (O_1177,N_29811,N_29766);
nand UO_1178 (O_1178,N_29939,N_29776);
nor UO_1179 (O_1179,N_29792,N_29875);
nor UO_1180 (O_1180,N_29984,N_29774);
or UO_1181 (O_1181,N_29776,N_29926);
and UO_1182 (O_1182,N_29712,N_29941);
and UO_1183 (O_1183,N_29901,N_29938);
and UO_1184 (O_1184,N_29804,N_29837);
nand UO_1185 (O_1185,N_29962,N_29945);
xnor UO_1186 (O_1186,N_29762,N_29927);
nor UO_1187 (O_1187,N_29703,N_29859);
nand UO_1188 (O_1188,N_29906,N_29756);
nor UO_1189 (O_1189,N_29704,N_29869);
xnor UO_1190 (O_1190,N_29738,N_29804);
xnor UO_1191 (O_1191,N_29780,N_29971);
or UO_1192 (O_1192,N_29787,N_29839);
xor UO_1193 (O_1193,N_29701,N_29802);
and UO_1194 (O_1194,N_29823,N_29973);
xnor UO_1195 (O_1195,N_29815,N_29708);
or UO_1196 (O_1196,N_29997,N_29931);
xor UO_1197 (O_1197,N_29989,N_29795);
xor UO_1198 (O_1198,N_29830,N_29910);
nor UO_1199 (O_1199,N_29706,N_29916);
or UO_1200 (O_1200,N_29748,N_29994);
nand UO_1201 (O_1201,N_29880,N_29848);
xor UO_1202 (O_1202,N_29733,N_29976);
and UO_1203 (O_1203,N_29918,N_29708);
or UO_1204 (O_1204,N_29733,N_29701);
nand UO_1205 (O_1205,N_29838,N_29872);
nor UO_1206 (O_1206,N_29922,N_29943);
nand UO_1207 (O_1207,N_29721,N_29738);
nand UO_1208 (O_1208,N_29887,N_29769);
and UO_1209 (O_1209,N_29988,N_29776);
or UO_1210 (O_1210,N_29850,N_29744);
or UO_1211 (O_1211,N_29969,N_29741);
nor UO_1212 (O_1212,N_29929,N_29963);
xnor UO_1213 (O_1213,N_29913,N_29774);
nand UO_1214 (O_1214,N_29916,N_29805);
or UO_1215 (O_1215,N_29813,N_29835);
nor UO_1216 (O_1216,N_29773,N_29729);
xor UO_1217 (O_1217,N_29749,N_29934);
and UO_1218 (O_1218,N_29947,N_29929);
nand UO_1219 (O_1219,N_29728,N_29908);
or UO_1220 (O_1220,N_29882,N_29916);
nor UO_1221 (O_1221,N_29958,N_29903);
or UO_1222 (O_1222,N_29798,N_29733);
xnor UO_1223 (O_1223,N_29726,N_29870);
xnor UO_1224 (O_1224,N_29973,N_29995);
nand UO_1225 (O_1225,N_29758,N_29991);
nand UO_1226 (O_1226,N_29764,N_29790);
nor UO_1227 (O_1227,N_29913,N_29847);
or UO_1228 (O_1228,N_29853,N_29703);
and UO_1229 (O_1229,N_29958,N_29937);
and UO_1230 (O_1230,N_29723,N_29899);
xor UO_1231 (O_1231,N_29990,N_29944);
and UO_1232 (O_1232,N_29784,N_29716);
or UO_1233 (O_1233,N_29752,N_29990);
and UO_1234 (O_1234,N_29847,N_29737);
nor UO_1235 (O_1235,N_29720,N_29881);
nor UO_1236 (O_1236,N_29766,N_29916);
or UO_1237 (O_1237,N_29998,N_29992);
nand UO_1238 (O_1238,N_29767,N_29951);
nand UO_1239 (O_1239,N_29954,N_29845);
nor UO_1240 (O_1240,N_29702,N_29844);
nand UO_1241 (O_1241,N_29819,N_29927);
nand UO_1242 (O_1242,N_29956,N_29951);
or UO_1243 (O_1243,N_29843,N_29935);
nand UO_1244 (O_1244,N_29801,N_29826);
and UO_1245 (O_1245,N_29713,N_29868);
nand UO_1246 (O_1246,N_29958,N_29862);
nand UO_1247 (O_1247,N_29811,N_29728);
and UO_1248 (O_1248,N_29879,N_29798);
xnor UO_1249 (O_1249,N_29912,N_29856);
nand UO_1250 (O_1250,N_29705,N_29977);
nor UO_1251 (O_1251,N_29780,N_29738);
nor UO_1252 (O_1252,N_29917,N_29796);
and UO_1253 (O_1253,N_29933,N_29727);
nor UO_1254 (O_1254,N_29710,N_29750);
nand UO_1255 (O_1255,N_29747,N_29991);
and UO_1256 (O_1256,N_29969,N_29796);
and UO_1257 (O_1257,N_29773,N_29886);
or UO_1258 (O_1258,N_29884,N_29765);
xor UO_1259 (O_1259,N_29857,N_29715);
xnor UO_1260 (O_1260,N_29874,N_29867);
nor UO_1261 (O_1261,N_29735,N_29983);
nor UO_1262 (O_1262,N_29742,N_29985);
nand UO_1263 (O_1263,N_29907,N_29743);
nand UO_1264 (O_1264,N_29947,N_29936);
xnor UO_1265 (O_1265,N_29747,N_29882);
and UO_1266 (O_1266,N_29822,N_29990);
nor UO_1267 (O_1267,N_29904,N_29905);
or UO_1268 (O_1268,N_29721,N_29796);
nand UO_1269 (O_1269,N_29745,N_29746);
nand UO_1270 (O_1270,N_29822,N_29737);
and UO_1271 (O_1271,N_29827,N_29735);
or UO_1272 (O_1272,N_29828,N_29773);
or UO_1273 (O_1273,N_29808,N_29964);
nand UO_1274 (O_1274,N_29801,N_29872);
nor UO_1275 (O_1275,N_29702,N_29904);
and UO_1276 (O_1276,N_29850,N_29891);
nand UO_1277 (O_1277,N_29971,N_29950);
nor UO_1278 (O_1278,N_29884,N_29976);
nor UO_1279 (O_1279,N_29733,N_29742);
and UO_1280 (O_1280,N_29775,N_29925);
nand UO_1281 (O_1281,N_29847,N_29907);
or UO_1282 (O_1282,N_29848,N_29709);
and UO_1283 (O_1283,N_29987,N_29904);
nor UO_1284 (O_1284,N_29889,N_29768);
nand UO_1285 (O_1285,N_29740,N_29832);
and UO_1286 (O_1286,N_29995,N_29891);
or UO_1287 (O_1287,N_29987,N_29901);
nor UO_1288 (O_1288,N_29743,N_29884);
xor UO_1289 (O_1289,N_29898,N_29791);
nand UO_1290 (O_1290,N_29988,N_29986);
xnor UO_1291 (O_1291,N_29752,N_29925);
and UO_1292 (O_1292,N_29724,N_29742);
nor UO_1293 (O_1293,N_29729,N_29719);
or UO_1294 (O_1294,N_29739,N_29757);
nor UO_1295 (O_1295,N_29782,N_29903);
or UO_1296 (O_1296,N_29728,N_29948);
and UO_1297 (O_1297,N_29998,N_29946);
nand UO_1298 (O_1298,N_29944,N_29865);
and UO_1299 (O_1299,N_29764,N_29708);
xor UO_1300 (O_1300,N_29933,N_29850);
and UO_1301 (O_1301,N_29752,N_29967);
nor UO_1302 (O_1302,N_29703,N_29903);
nor UO_1303 (O_1303,N_29842,N_29862);
nand UO_1304 (O_1304,N_29842,N_29760);
or UO_1305 (O_1305,N_29809,N_29797);
nand UO_1306 (O_1306,N_29876,N_29715);
xor UO_1307 (O_1307,N_29734,N_29852);
nand UO_1308 (O_1308,N_29746,N_29737);
xnor UO_1309 (O_1309,N_29779,N_29928);
nor UO_1310 (O_1310,N_29905,N_29927);
or UO_1311 (O_1311,N_29910,N_29857);
nor UO_1312 (O_1312,N_29935,N_29945);
nand UO_1313 (O_1313,N_29881,N_29930);
or UO_1314 (O_1314,N_29758,N_29824);
and UO_1315 (O_1315,N_29744,N_29826);
nand UO_1316 (O_1316,N_29858,N_29828);
nor UO_1317 (O_1317,N_29714,N_29851);
xor UO_1318 (O_1318,N_29777,N_29804);
nor UO_1319 (O_1319,N_29819,N_29868);
nand UO_1320 (O_1320,N_29930,N_29864);
or UO_1321 (O_1321,N_29944,N_29969);
nor UO_1322 (O_1322,N_29770,N_29783);
or UO_1323 (O_1323,N_29917,N_29742);
nor UO_1324 (O_1324,N_29832,N_29930);
nand UO_1325 (O_1325,N_29771,N_29702);
and UO_1326 (O_1326,N_29887,N_29823);
nand UO_1327 (O_1327,N_29923,N_29876);
xnor UO_1328 (O_1328,N_29918,N_29944);
nor UO_1329 (O_1329,N_29951,N_29906);
or UO_1330 (O_1330,N_29925,N_29911);
and UO_1331 (O_1331,N_29973,N_29890);
nor UO_1332 (O_1332,N_29833,N_29952);
nor UO_1333 (O_1333,N_29801,N_29888);
or UO_1334 (O_1334,N_29739,N_29838);
nor UO_1335 (O_1335,N_29939,N_29703);
and UO_1336 (O_1336,N_29824,N_29855);
and UO_1337 (O_1337,N_29974,N_29785);
xor UO_1338 (O_1338,N_29852,N_29985);
nor UO_1339 (O_1339,N_29848,N_29859);
and UO_1340 (O_1340,N_29926,N_29999);
nand UO_1341 (O_1341,N_29920,N_29810);
nor UO_1342 (O_1342,N_29992,N_29779);
and UO_1343 (O_1343,N_29738,N_29731);
nor UO_1344 (O_1344,N_29985,N_29851);
nor UO_1345 (O_1345,N_29733,N_29744);
or UO_1346 (O_1346,N_29888,N_29821);
or UO_1347 (O_1347,N_29771,N_29717);
or UO_1348 (O_1348,N_29972,N_29941);
xor UO_1349 (O_1349,N_29763,N_29721);
xnor UO_1350 (O_1350,N_29985,N_29901);
nor UO_1351 (O_1351,N_29882,N_29925);
and UO_1352 (O_1352,N_29915,N_29810);
and UO_1353 (O_1353,N_29845,N_29764);
nor UO_1354 (O_1354,N_29922,N_29771);
and UO_1355 (O_1355,N_29733,N_29765);
nor UO_1356 (O_1356,N_29754,N_29865);
or UO_1357 (O_1357,N_29832,N_29784);
xnor UO_1358 (O_1358,N_29706,N_29870);
xor UO_1359 (O_1359,N_29873,N_29852);
or UO_1360 (O_1360,N_29724,N_29854);
and UO_1361 (O_1361,N_29899,N_29859);
and UO_1362 (O_1362,N_29849,N_29919);
and UO_1363 (O_1363,N_29908,N_29788);
and UO_1364 (O_1364,N_29874,N_29854);
nand UO_1365 (O_1365,N_29730,N_29706);
nor UO_1366 (O_1366,N_29784,N_29983);
or UO_1367 (O_1367,N_29854,N_29911);
nand UO_1368 (O_1368,N_29886,N_29918);
nand UO_1369 (O_1369,N_29851,N_29944);
nor UO_1370 (O_1370,N_29874,N_29905);
or UO_1371 (O_1371,N_29700,N_29756);
or UO_1372 (O_1372,N_29870,N_29868);
xor UO_1373 (O_1373,N_29747,N_29846);
nor UO_1374 (O_1374,N_29732,N_29968);
and UO_1375 (O_1375,N_29789,N_29883);
nor UO_1376 (O_1376,N_29819,N_29842);
and UO_1377 (O_1377,N_29935,N_29867);
nor UO_1378 (O_1378,N_29768,N_29732);
or UO_1379 (O_1379,N_29796,N_29941);
nor UO_1380 (O_1380,N_29721,N_29843);
nor UO_1381 (O_1381,N_29789,N_29776);
nor UO_1382 (O_1382,N_29731,N_29755);
nor UO_1383 (O_1383,N_29881,N_29927);
nor UO_1384 (O_1384,N_29777,N_29788);
nand UO_1385 (O_1385,N_29816,N_29957);
or UO_1386 (O_1386,N_29824,N_29825);
nor UO_1387 (O_1387,N_29892,N_29792);
and UO_1388 (O_1388,N_29832,N_29822);
or UO_1389 (O_1389,N_29939,N_29802);
xor UO_1390 (O_1390,N_29972,N_29963);
or UO_1391 (O_1391,N_29940,N_29891);
or UO_1392 (O_1392,N_29929,N_29883);
and UO_1393 (O_1393,N_29890,N_29835);
nand UO_1394 (O_1394,N_29721,N_29969);
nand UO_1395 (O_1395,N_29986,N_29709);
or UO_1396 (O_1396,N_29831,N_29812);
xor UO_1397 (O_1397,N_29732,N_29895);
or UO_1398 (O_1398,N_29974,N_29705);
or UO_1399 (O_1399,N_29822,N_29935);
or UO_1400 (O_1400,N_29776,N_29968);
or UO_1401 (O_1401,N_29917,N_29859);
nand UO_1402 (O_1402,N_29780,N_29851);
and UO_1403 (O_1403,N_29784,N_29754);
and UO_1404 (O_1404,N_29737,N_29811);
or UO_1405 (O_1405,N_29741,N_29961);
xnor UO_1406 (O_1406,N_29765,N_29889);
and UO_1407 (O_1407,N_29848,N_29736);
or UO_1408 (O_1408,N_29901,N_29857);
nor UO_1409 (O_1409,N_29861,N_29710);
nor UO_1410 (O_1410,N_29799,N_29918);
and UO_1411 (O_1411,N_29719,N_29933);
nand UO_1412 (O_1412,N_29995,N_29713);
or UO_1413 (O_1413,N_29853,N_29720);
xnor UO_1414 (O_1414,N_29939,N_29908);
and UO_1415 (O_1415,N_29968,N_29820);
xor UO_1416 (O_1416,N_29975,N_29731);
nor UO_1417 (O_1417,N_29739,N_29797);
xnor UO_1418 (O_1418,N_29849,N_29973);
and UO_1419 (O_1419,N_29706,N_29903);
xnor UO_1420 (O_1420,N_29924,N_29765);
nand UO_1421 (O_1421,N_29976,N_29734);
and UO_1422 (O_1422,N_29946,N_29855);
nor UO_1423 (O_1423,N_29842,N_29791);
and UO_1424 (O_1424,N_29852,N_29820);
nand UO_1425 (O_1425,N_29766,N_29877);
nor UO_1426 (O_1426,N_29796,N_29776);
or UO_1427 (O_1427,N_29885,N_29901);
or UO_1428 (O_1428,N_29756,N_29910);
nor UO_1429 (O_1429,N_29853,N_29737);
xnor UO_1430 (O_1430,N_29830,N_29753);
nand UO_1431 (O_1431,N_29836,N_29906);
xnor UO_1432 (O_1432,N_29969,N_29889);
and UO_1433 (O_1433,N_29727,N_29935);
nand UO_1434 (O_1434,N_29750,N_29822);
and UO_1435 (O_1435,N_29708,N_29825);
nand UO_1436 (O_1436,N_29741,N_29806);
or UO_1437 (O_1437,N_29911,N_29883);
nor UO_1438 (O_1438,N_29890,N_29815);
nand UO_1439 (O_1439,N_29763,N_29773);
xnor UO_1440 (O_1440,N_29972,N_29802);
nand UO_1441 (O_1441,N_29797,N_29927);
nor UO_1442 (O_1442,N_29832,N_29710);
or UO_1443 (O_1443,N_29809,N_29708);
or UO_1444 (O_1444,N_29853,N_29925);
xnor UO_1445 (O_1445,N_29829,N_29840);
nand UO_1446 (O_1446,N_29970,N_29839);
or UO_1447 (O_1447,N_29780,N_29764);
nor UO_1448 (O_1448,N_29988,N_29982);
xnor UO_1449 (O_1449,N_29739,N_29925);
nand UO_1450 (O_1450,N_29814,N_29957);
xor UO_1451 (O_1451,N_29960,N_29920);
and UO_1452 (O_1452,N_29907,N_29940);
or UO_1453 (O_1453,N_29741,N_29953);
nand UO_1454 (O_1454,N_29985,N_29801);
nand UO_1455 (O_1455,N_29719,N_29846);
nor UO_1456 (O_1456,N_29826,N_29964);
nand UO_1457 (O_1457,N_29703,N_29980);
and UO_1458 (O_1458,N_29734,N_29977);
nor UO_1459 (O_1459,N_29874,N_29805);
and UO_1460 (O_1460,N_29959,N_29866);
nand UO_1461 (O_1461,N_29753,N_29747);
and UO_1462 (O_1462,N_29851,N_29983);
xnor UO_1463 (O_1463,N_29730,N_29991);
and UO_1464 (O_1464,N_29880,N_29973);
nand UO_1465 (O_1465,N_29742,N_29989);
or UO_1466 (O_1466,N_29888,N_29903);
nor UO_1467 (O_1467,N_29778,N_29796);
or UO_1468 (O_1468,N_29804,N_29929);
nor UO_1469 (O_1469,N_29706,N_29859);
nand UO_1470 (O_1470,N_29926,N_29860);
nor UO_1471 (O_1471,N_29986,N_29965);
xor UO_1472 (O_1472,N_29776,N_29801);
nor UO_1473 (O_1473,N_29886,N_29787);
and UO_1474 (O_1474,N_29894,N_29717);
nand UO_1475 (O_1475,N_29903,N_29954);
xor UO_1476 (O_1476,N_29721,N_29734);
xor UO_1477 (O_1477,N_29956,N_29835);
and UO_1478 (O_1478,N_29818,N_29817);
and UO_1479 (O_1479,N_29769,N_29817);
nor UO_1480 (O_1480,N_29890,N_29924);
xnor UO_1481 (O_1481,N_29912,N_29904);
nand UO_1482 (O_1482,N_29931,N_29784);
nor UO_1483 (O_1483,N_29905,N_29768);
xnor UO_1484 (O_1484,N_29894,N_29826);
nand UO_1485 (O_1485,N_29988,N_29831);
nor UO_1486 (O_1486,N_29883,N_29706);
nand UO_1487 (O_1487,N_29799,N_29961);
xor UO_1488 (O_1488,N_29971,N_29728);
nand UO_1489 (O_1489,N_29792,N_29843);
nand UO_1490 (O_1490,N_29708,N_29787);
nand UO_1491 (O_1491,N_29797,N_29877);
xnor UO_1492 (O_1492,N_29761,N_29869);
and UO_1493 (O_1493,N_29988,N_29841);
nor UO_1494 (O_1494,N_29727,N_29711);
or UO_1495 (O_1495,N_29819,N_29736);
or UO_1496 (O_1496,N_29761,N_29899);
nor UO_1497 (O_1497,N_29813,N_29911);
or UO_1498 (O_1498,N_29728,N_29700);
xor UO_1499 (O_1499,N_29768,N_29926);
nand UO_1500 (O_1500,N_29930,N_29815);
and UO_1501 (O_1501,N_29945,N_29981);
xor UO_1502 (O_1502,N_29836,N_29967);
and UO_1503 (O_1503,N_29728,N_29775);
nor UO_1504 (O_1504,N_29970,N_29829);
or UO_1505 (O_1505,N_29890,N_29703);
xnor UO_1506 (O_1506,N_29735,N_29968);
nand UO_1507 (O_1507,N_29957,N_29800);
nand UO_1508 (O_1508,N_29716,N_29780);
and UO_1509 (O_1509,N_29962,N_29771);
nand UO_1510 (O_1510,N_29909,N_29700);
or UO_1511 (O_1511,N_29765,N_29792);
nor UO_1512 (O_1512,N_29874,N_29965);
and UO_1513 (O_1513,N_29705,N_29769);
nand UO_1514 (O_1514,N_29830,N_29844);
nor UO_1515 (O_1515,N_29705,N_29975);
nand UO_1516 (O_1516,N_29961,N_29744);
and UO_1517 (O_1517,N_29970,N_29871);
xnor UO_1518 (O_1518,N_29815,N_29923);
nand UO_1519 (O_1519,N_29985,N_29798);
nor UO_1520 (O_1520,N_29992,N_29749);
nor UO_1521 (O_1521,N_29913,N_29773);
and UO_1522 (O_1522,N_29881,N_29826);
nand UO_1523 (O_1523,N_29949,N_29756);
nand UO_1524 (O_1524,N_29870,N_29766);
xor UO_1525 (O_1525,N_29945,N_29863);
nor UO_1526 (O_1526,N_29785,N_29944);
and UO_1527 (O_1527,N_29741,N_29836);
and UO_1528 (O_1528,N_29720,N_29884);
or UO_1529 (O_1529,N_29710,N_29949);
or UO_1530 (O_1530,N_29852,N_29976);
xor UO_1531 (O_1531,N_29927,N_29705);
nor UO_1532 (O_1532,N_29875,N_29954);
nand UO_1533 (O_1533,N_29943,N_29941);
nand UO_1534 (O_1534,N_29853,N_29867);
or UO_1535 (O_1535,N_29983,N_29835);
and UO_1536 (O_1536,N_29786,N_29840);
nand UO_1537 (O_1537,N_29886,N_29761);
and UO_1538 (O_1538,N_29941,N_29769);
nor UO_1539 (O_1539,N_29704,N_29965);
nor UO_1540 (O_1540,N_29859,N_29700);
and UO_1541 (O_1541,N_29767,N_29844);
nor UO_1542 (O_1542,N_29876,N_29860);
nor UO_1543 (O_1543,N_29779,N_29725);
xor UO_1544 (O_1544,N_29894,N_29913);
and UO_1545 (O_1545,N_29828,N_29862);
nor UO_1546 (O_1546,N_29955,N_29759);
nand UO_1547 (O_1547,N_29981,N_29879);
and UO_1548 (O_1548,N_29935,N_29825);
or UO_1549 (O_1549,N_29982,N_29850);
nand UO_1550 (O_1550,N_29814,N_29928);
and UO_1551 (O_1551,N_29940,N_29755);
xnor UO_1552 (O_1552,N_29907,N_29913);
nand UO_1553 (O_1553,N_29909,N_29703);
nor UO_1554 (O_1554,N_29748,N_29960);
or UO_1555 (O_1555,N_29882,N_29841);
xor UO_1556 (O_1556,N_29937,N_29889);
nor UO_1557 (O_1557,N_29989,N_29923);
or UO_1558 (O_1558,N_29790,N_29895);
nor UO_1559 (O_1559,N_29724,N_29736);
xor UO_1560 (O_1560,N_29841,N_29950);
nand UO_1561 (O_1561,N_29899,N_29749);
or UO_1562 (O_1562,N_29904,N_29920);
and UO_1563 (O_1563,N_29812,N_29810);
nand UO_1564 (O_1564,N_29929,N_29844);
xnor UO_1565 (O_1565,N_29849,N_29834);
nor UO_1566 (O_1566,N_29726,N_29832);
and UO_1567 (O_1567,N_29859,N_29824);
and UO_1568 (O_1568,N_29935,N_29923);
xor UO_1569 (O_1569,N_29740,N_29979);
xor UO_1570 (O_1570,N_29933,N_29908);
nand UO_1571 (O_1571,N_29830,N_29967);
xnor UO_1572 (O_1572,N_29988,N_29970);
or UO_1573 (O_1573,N_29998,N_29713);
nor UO_1574 (O_1574,N_29851,N_29931);
nor UO_1575 (O_1575,N_29758,N_29819);
nand UO_1576 (O_1576,N_29845,N_29959);
nor UO_1577 (O_1577,N_29941,N_29794);
nor UO_1578 (O_1578,N_29964,N_29807);
and UO_1579 (O_1579,N_29876,N_29723);
or UO_1580 (O_1580,N_29895,N_29808);
nand UO_1581 (O_1581,N_29924,N_29821);
nand UO_1582 (O_1582,N_29907,N_29752);
xnor UO_1583 (O_1583,N_29939,N_29729);
and UO_1584 (O_1584,N_29921,N_29738);
xnor UO_1585 (O_1585,N_29856,N_29938);
xor UO_1586 (O_1586,N_29898,N_29723);
nand UO_1587 (O_1587,N_29708,N_29882);
or UO_1588 (O_1588,N_29763,N_29908);
xnor UO_1589 (O_1589,N_29731,N_29945);
nand UO_1590 (O_1590,N_29815,N_29798);
xnor UO_1591 (O_1591,N_29940,N_29713);
and UO_1592 (O_1592,N_29706,N_29775);
nor UO_1593 (O_1593,N_29799,N_29828);
xnor UO_1594 (O_1594,N_29886,N_29905);
xor UO_1595 (O_1595,N_29932,N_29780);
nor UO_1596 (O_1596,N_29909,N_29936);
and UO_1597 (O_1597,N_29743,N_29782);
or UO_1598 (O_1598,N_29720,N_29984);
xor UO_1599 (O_1599,N_29750,N_29988);
xor UO_1600 (O_1600,N_29940,N_29772);
nand UO_1601 (O_1601,N_29823,N_29723);
nor UO_1602 (O_1602,N_29707,N_29795);
nor UO_1603 (O_1603,N_29904,N_29948);
nor UO_1604 (O_1604,N_29783,N_29978);
or UO_1605 (O_1605,N_29905,N_29893);
and UO_1606 (O_1606,N_29907,N_29928);
nand UO_1607 (O_1607,N_29753,N_29983);
nand UO_1608 (O_1608,N_29899,N_29783);
nand UO_1609 (O_1609,N_29933,N_29773);
nor UO_1610 (O_1610,N_29759,N_29795);
nand UO_1611 (O_1611,N_29955,N_29719);
and UO_1612 (O_1612,N_29748,N_29992);
or UO_1613 (O_1613,N_29865,N_29740);
nand UO_1614 (O_1614,N_29707,N_29987);
nand UO_1615 (O_1615,N_29732,N_29777);
xor UO_1616 (O_1616,N_29875,N_29704);
or UO_1617 (O_1617,N_29872,N_29863);
or UO_1618 (O_1618,N_29764,N_29828);
or UO_1619 (O_1619,N_29937,N_29807);
and UO_1620 (O_1620,N_29710,N_29701);
nand UO_1621 (O_1621,N_29945,N_29750);
or UO_1622 (O_1622,N_29708,N_29998);
and UO_1623 (O_1623,N_29803,N_29989);
xnor UO_1624 (O_1624,N_29828,N_29842);
nor UO_1625 (O_1625,N_29750,N_29785);
xor UO_1626 (O_1626,N_29811,N_29987);
and UO_1627 (O_1627,N_29798,N_29857);
or UO_1628 (O_1628,N_29958,N_29938);
nand UO_1629 (O_1629,N_29933,N_29876);
xnor UO_1630 (O_1630,N_29856,N_29719);
nor UO_1631 (O_1631,N_29703,N_29882);
and UO_1632 (O_1632,N_29809,N_29823);
nor UO_1633 (O_1633,N_29811,N_29711);
or UO_1634 (O_1634,N_29851,N_29913);
or UO_1635 (O_1635,N_29806,N_29864);
nor UO_1636 (O_1636,N_29775,N_29838);
nor UO_1637 (O_1637,N_29775,N_29981);
or UO_1638 (O_1638,N_29710,N_29904);
xor UO_1639 (O_1639,N_29897,N_29973);
or UO_1640 (O_1640,N_29925,N_29906);
or UO_1641 (O_1641,N_29998,N_29756);
and UO_1642 (O_1642,N_29926,N_29773);
nor UO_1643 (O_1643,N_29913,N_29957);
and UO_1644 (O_1644,N_29903,N_29802);
nand UO_1645 (O_1645,N_29971,N_29804);
and UO_1646 (O_1646,N_29735,N_29743);
nand UO_1647 (O_1647,N_29980,N_29876);
or UO_1648 (O_1648,N_29708,N_29734);
xnor UO_1649 (O_1649,N_29854,N_29879);
or UO_1650 (O_1650,N_29781,N_29718);
nor UO_1651 (O_1651,N_29819,N_29932);
nand UO_1652 (O_1652,N_29935,N_29812);
or UO_1653 (O_1653,N_29783,N_29904);
nor UO_1654 (O_1654,N_29860,N_29893);
nand UO_1655 (O_1655,N_29959,N_29716);
or UO_1656 (O_1656,N_29954,N_29989);
nand UO_1657 (O_1657,N_29912,N_29772);
or UO_1658 (O_1658,N_29939,N_29748);
nor UO_1659 (O_1659,N_29788,N_29870);
nand UO_1660 (O_1660,N_29953,N_29772);
nand UO_1661 (O_1661,N_29736,N_29961);
xnor UO_1662 (O_1662,N_29991,N_29858);
or UO_1663 (O_1663,N_29893,N_29867);
nor UO_1664 (O_1664,N_29977,N_29852);
nor UO_1665 (O_1665,N_29795,N_29723);
or UO_1666 (O_1666,N_29869,N_29983);
xnor UO_1667 (O_1667,N_29767,N_29872);
nand UO_1668 (O_1668,N_29967,N_29918);
or UO_1669 (O_1669,N_29932,N_29846);
and UO_1670 (O_1670,N_29831,N_29840);
and UO_1671 (O_1671,N_29742,N_29721);
nor UO_1672 (O_1672,N_29824,N_29754);
nand UO_1673 (O_1673,N_29956,N_29813);
and UO_1674 (O_1674,N_29924,N_29870);
nand UO_1675 (O_1675,N_29899,N_29945);
nor UO_1676 (O_1676,N_29758,N_29710);
or UO_1677 (O_1677,N_29975,N_29713);
nand UO_1678 (O_1678,N_29831,N_29752);
xor UO_1679 (O_1679,N_29894,N_29918);
or UO_1680 (O_1680,N_29875,N_29956);
and UO_1681 (O_1681,N_29815,N_29860);
xnor UO_1682 (O_1682,N_29970,N_29857);
nor UO_1683 (O_1683,N_29734,N_29971);
xor UO_1684 (O_1684,N_29730,N_29890);
and UO_1685 (O_1685,N_29965,N_29721);
or UO_1686 (O_1686,N_29787,N_29806);
nand UO_1687 (O_1687,N_29885,N_29728);
or UO_1688 (O_1688,N_29756,N_29816);
or UO_1689 (O_1689,N_29814,N_29709);
xor UO_1690 (O_1690,N_29843,N_29716);
or UO_1691 (O_1691,N_29879,N_29903);
nor UO_1692 (O_1692,N_29995,N_29797);
xnor UO_1693 (O_1693,N_29903,N_29996);
nand UO_1694 (O_1694,N_29948,N_29873);
xor UO_1695 (O_1695,N_29781,N_29747);
xor UO_1696 (O_1696,N_29715,N_29934);
or UO_1697 (O_1697,N_29871,N_29829);
or UO_1698 (O_1698,N_29714,N_29843);
and UO_1699 (O_1699,N_29814,N_29706);
or UO_1700 (O_1700,N_29755,N_29776);
and UO_1701 (O_1701,N_29994,N_29746);
xor UO_1702 (O_1702,N_29704,N_29881);
or UO_1703 (O_1703,N_29983,N_29992);
and UO_1704 (O_1704,N_29827,N_29997);
or UO_1705 (O_1705,N_29904,N_29880);
or UO_1706 (O_1706,N_29987,N_29749);
and UO_1707 (O_1707,N_29760,N_29724);
or UO_1708 (O_1708,N_29753,N_29902);
and UO_1709 (O_1709,N_29811,N_29988);
and UO_1710 (O_1710,N_29858,N_29910);
nor UO_1711 (O_1711,N_29945,N_29719);
xor UO_1712 (O_1712,N_29892,N_29935);
xnor UO_1713 (O_1713,N_29992,N_29707);
xor UO_1714 (O_1714,N_29835,N_29934);
and UO_1715 (O_1715,N_29989,N_29708);
or UO_1716 (O_1716,N_29740,N_29773);
and UO_1717 (O_1717,N_29782,N_29723);
nor UO_1718 (O_1718,N_29701,N_29832);
xor UO_1719 (O_1719,N_29859,N_29791);
and UO_1720 (O_1720,N_29824,N_29923);
nor UO_1721 (O_1721,N_29991,N_29713);
xnor UO_1722 (O_1722,N_29869,N_29802);
and UO_1723 (O_1723,N_29914,N_29970);
xor UO_1724 (O_1724,N_29815,N_29888);
xor UO_1725 (O_1725,N_29984,N_29937);
and UO_1726 (O_1726,N_29723,N_29908);
and UO_1727 (O_1727,N_29851,N_29754);
nor UO_1728 (O_1728,N_29735,N_29949);
xnor UO_1729 (O_1729,N_29765,N_29793);
nor UO_1730 (O_1730,N_29987,N_29842);
nor UO_1731 (O_1731,N_29714,N_29738);
nor UO_1732 (O_1732,N_29993,N_29805);
xor UO_1733 (O_1733,N_29984,N_29889);
nor UO_1734 (O_1734,N_29851,N_29900);
or UO_1735 (O_1735,N_29955,N_29838);
and UO_1736 (O_1736,N_29868,N_29768);
and UO_1737 (O_1737,N_29805,N_29980);
xor UO_1738 (O_1738,N_29892,N_29977);
nand UO_1739 (O_1739,N_29926,N_29804);
or UO_1740 (O_1740,N_29814,N_29739);
xnor UO_1741 (O_1741,N_29809,N_29982);
and UO_1742 (O_1742,N_29988,N_29932);
nand UO_1743 (O_1743,N_29736,N_29934);
and UO_1744 (O_1744,N_29865,N_29869);
or UO_1745 (O_1745,N_29882,N_29902);
nand UO_1746 (O_1746,N_29831,N_29819);
and UO_1747 (O_1747,N_29908,N_29966);
nor UO_1748 (O_1748,N_29807,N_29947);
and UO_1749 (O_1749,N_29870,N_29987);
or UO_1750 (O_1750,N_29975,N_29773);
nand UO_1751 (O_1751,N_29947,N_29856);
and UO_1752 (O_1752,N_29740,N_29733);
xor UO_1753 (O_1753,N_29723,N_29917);
or UO_1754 (O_1754,N_29814,N_29822);
and UO_1755 (O_1755,N_29895,N_29862);
nor UO_1756 (O_1756,N_29871,N_29858);
and UO_1757 (O_1757,N_29713,N_29720);
xor UO_1758 (O_1758,N_29710,N_29978);
xor UO_1759 (O_1759,N_29984,N_29888);
nand UO_1760 (O_1760,N_29989,N_29898);
and UO_1761 (O_1761,N_29775,N_29957);
or UO_1762 (O_1762,N_29903,N_29849);
nand UO_1763 (O_1763,N_29876,N_29884);
and UO_1764 (O_1764,N_29716,N_29720);
nand UO_1765 (O_1765,N_29906,N_29882);
nor UO_1766 (O_1766,N_29856,N_29986);
and UO_1767 (O_1767,N_29961,N_29852);
xnor UO_1768 (O_1768,N_29899,N_29709);
xor UO_1769 (O_1769,N_29944,N_29996);
xnor UO_1770 (O_1770,N_29811,N_29902);
nor UO_1771 (O_1771,N_29858,N_29708);
nand UO_1772 (O_1772,N_29813,N_29963);
nand UO_1773 (O_1773,N_29711,N_29920);
and UO_1774 (O_1774,N_29991,N_29954);
nor UO_1775 (O_1775,N_29800,N_29802);
nand UO_1776 (O_1776,N_29768,N_29717);
or UO_1777 (O_1777,N_29945,N_29847);
xnor UO_1778 (O_1778,N_29957,N_29834);
and UO_1779 (O_1779,N_29716,N_29768);
xor UO_1780 (O_1780,N_29939,N_29894);
nand UO_1781 (O_1781,N_29941,N_29744);
nor UO_1782 (O_1782,N_29991,N_29956);
nor UO_1783 (O_1783,N_29756,N_29819);
and UO_1784 (O_1784,N_29880,N_29719);
nand UO_1785 (O_1785,N_29981,N_29978);
and UO_1786 (O_1786,N_29861,N_29867);
or UO_1787 (O_1787,N_29931,N_29757);
or UO_1788 (O_1788,N_29769,N_29727);
nand UO_1789 (O_1789,N_29982,N_29705);
nand UO_1790 (O_1790,N_29881,N_29719);
xnor UO_1791 (O_1791,N_29832,N_29986);
xnor UO_1792 (O_1792,N_29776,N_29716);
and UO_1793 (O_1793,N_29780,N_29719);
nand UO_1794 (O_1794,N_29922,N_29871);
or UO_1795 (O_1795,N_29971,N_29849);
nor UO_1796 (O_1796,N_29849,N_29765);
xnor UO_1797 (O_1797,N_29780,N_29830);
and UO_1798 (O_1798,N_29901,N_29761);
xnor UO_1799 (O_1799,N_29927,N_29825);
nor UO_1800 (O_1800,N_29893,N_29962);
nand UO_1801 (O_1801,N_29887,N_29917);
and UO_1802 (O_1802,N_29767,N_29837);
xor UO_1803 (O_1803,N_29962,N_29772);
or UO_1804 (O_1804,N_29963,N_29861);
xnor UO_1805 (O_1805,N_29841,N_29754);
nand UO_1806 (O_1806,N_29813,N_29964);
and UO_1807 (O_1807,N_29884,N_29880);
or UO_1808 (O_1808,N_29972,N_29834);
or UO_1809 (O_1809,N_29718,N_29964);
and UO_1810 (O_1810,N_29855,N_29963);
nand UO_1811 (O_1811,N_29879,N_29836);
or UO_1812 (O_1812,N_29764,N_29937);
nand UO_1813 (O_1813,N_29998,N_29765);
nor UO_1814 (O_1814,N_29877,N_29705);
or UO_1815 (O_1815,N_29902,N_29741);
nand UO_1816 (O_1816,N_29841,N_29964);
or UO_1817 (O_1817,N_29839,N_29761);
nand UO_1818 (O_1818,N_29825,N_29872);
nand UO_1819 (O_1819,N_29966,N_29976);
nor UO_1820 (O_1820,N_29815,N_29768);
nor UO_1821 (O_1821,N_29985,N_29774);
and UO_1822 (O_1822,N_29889,N_29767);
xor UO_1823 (O_1823,N_29774,N_29925);
and UO_1824 (O_1824,N_29857,N_29986);
nor UO_1825 (O_1825,N_29737,N_29937);
xnor UO_1826 (O_1826,N_29761,N_29912);
xnor UO_1827 (O_1827,N_29839,N_29977);
and UO_1828 (O_1828,N_29855,N_29786);
nand UO_1829 (O_1829,N_29948,N_29741);
xnor UO_1830 (O_1830,N_29722,N_29988);
nand UO_1831 (O_1831,N_29959,N_29899);
xor UO_1832 (O_1832,N_29758,N_29924);
nand UO_1833 (O_1833,N_29922,N_29999);
xnor UO_1834 (O_1834,N_29940,N_29875);
xor UO_1835 (O_1835,N_29770,N_29992);
or UO_1836 (O_1836,N_29732,N_29981);
nor UO_1837 (O_1837,N_29824,N_29819);
nand UO_1838 (O_1838,N_29774,N_29871);
and UO_1839 (O_1839,N_29906,N_29743);
xor UO_1840 (O_1840,N_29918,N_29807);
xnor UO_1841 (O_1841,N_29814,N_29778);
nand UO_1842 (O_1842,N_29864,N_29970);
xor UO_1843 (O_1843,N_29761,N_29885);
and UO_1844 (O_1844,N_29798,N_29976);
nor UO_1845 (O_1845,N_29725,N_29747);
and UO_1846 (O_1846,N_29812,N_29914);
nand UO_1847 (O_1847,N_29833,N_29941);
nand UO_1848 (O_1848,N_29959,N_29927);
and UO_1849 (O_1849,N_29836,N_29856);
and UO_1850 (O_1850,N_29706,N_29767);
nand UO_1851 (O_1851,N_29759,N_29805);
or UO_1852 (O_1852,N_29884,N_29748);
or UO_1853 (O_1853,N_29846,N_29701);
xnor UO_1854 (O_1854,N_29943,N_29857);
nand UO_1855 (O_1855,N_29856,N_29939);
nor UO_1856 (O_1856,N_29743,N_29959);
nor UO_1857 (O_1857,N_29799,N_29959);
or UO_1858 (O_1858,N_29964,N_29821);
nand UO_1859 (O_1859,N_29740,N_29709);
or UO_1860 (O_1860,N_29825,N_29917);
and UO_1861 (O_1861,N_29941,N_29933);
xnor UO_1862 (O_1862,N_29843,N_29986);
nor UO_1863 (O_1863,N_29846,N_29866);
xnor UO_1864 (O_1864,N_29910,N_29939);
or UO_1865 (O_1865,N_29825,N_29823);
and UO_1866 (O_1866,N_29819,N_29826);
xnor UO_1867 (O_1867,N_29827,N_29945);
nor UO_1868 (O_1868,N_29880,N_29796);
or UO_1869 (O_1869,N_29987,N_29978);
nor UO_1870 (O_1870,N_29835,N_29861);
xnor UO_1871 (O_1871,N_29882,N_29733);
nand UO_1872 (O_1872,N_29934,N_29811);
and UO_1873 (O_1873,N_29866,N_29794);
nor UO_1874 (O_1874,N_29717,N_29836);
nor UO_1875 (O_1875,N_29911,N_29837);
nand UO_1876 (O_1876,N_29981,N_29721);
nor UO_1877 (O_1877,N_29740,N_29850);
or UO_1878 (O_1878,N_29899,N_29815);
xor UO_1879 (O_1879,N_29870,N_29972);
nor UO_1880 (O_1880,N_29867,N_29881);
nor UO_1881 (O_1881,N_29971,N_29886);
nor UO_1882 (O_1882,N_29885,N_29747);
xnor UO_1883 (O_1883,N_29767,N_29762);
and UO_1884 (O_1884,N_29740,N_29983);
or UO_1885 (O_1885,N_29973,N_29744);
nor UO_1886 (O_1886,N_29882,N_29705);
or UO_1887 (O_1887,N_29979,N_29953);
or UO_1888 (O_1888,N_29781,N_29872);
or UO_1889 (O_1889,N_29794,N_29704);
or UO_1890 (O_1890,N_29863,N_29984);
nor UO_1891 (O_1891,N_29788,N_29936);
or UO_1892 (O_1892,N_29713,N_29966);
xnor UO_1893 (O_1893,N_29918,N_29749);
or UO_1894 (O_1894,N_29953,N_29751);
nor UO_1895 (O_1895,N_29908,N_29950);
xor UO_1896 (O_1896,N_29717,N_29994);
nand UO_1897 (O_1897,N_29977,N_29978);
or UO_1898 (O_1898,N_29774,N_29911);
nand UO_1899 (O_1899,N_29926,N_29723);
xor UO_1900 (O_1900,N_29806,N_29980);
or UO_1901 (O_1901,N_29927,N_29757);
nand UO_1902 (O_1902,N_29806,N_29863);
nor UO_1903 (O_1903,N_29948,N_29726);
or UO_1904 (O_1904,N_29895,N_29708);
xor UO_1905 (O_1905,N_29948,N_29747);
nand UO_1906 (O_1906,N_29966,N_29828);
nand UO_1907 (O_1907,N_29971,N_29912);
nand UO_1908 (O_1908,N_29820,N_29906);
nor UO_1909 (O_1909,N_29912,N_29943);
nor UO_1910 (O_1910,N_29716,N_29996);
or UO_1911 (O_1911,N_29970,N_29920);
and UO_1912 (O_1912,N_29818,N_29769);
and UO_1913 (O_1913,N_29925,N_29715);
or UO_1914 (O_1914,N_29753,N_29915);
or UO_1915 (O_1915,N_29958,N_29944);
and UO_1916 (O_1916,N_29969,N_29700);
nor UO_1917 (O_1917,N_29989,N_29990);
nor UO_1918 (O_1918,N_29758,N_29714);
nand UO_1919 (O_1919,N_29994,N_29812);
nand UO_1920 (O_1920,N_29795,N_29751);
nand UO_1921 (O_1921,N_29770,N_29809);
and UO_1922 (O_1922,N_29723,N_29755);
xnor UO_1923 (O_1923,N_29844,N_29832);
nor UO_1924 (O_1924,N_29949,N_29906);
nand UO_1925 (O_1925,N_29727,N_29794);
and UO_1926 (O_1926,N_29791,N_29987);
and UO_1927 (O_1927,N_29801,N_29912);
nand UO_1928 (O_1928,N_29929,N_29834);
or UO_1929 (O_1929,N_29867,N_29765);
xnor UO_1930 (O_1930,N_29931,N_29983);
nor UO_1931 (O_1931,N_29752,N_29984);
nand UO_1932 (O_1932,N_29771,N_29813);
or UO_1933 (O_1933,N_29844,N_29878);
and UO_1934 (O_1934,N_29901,N_29752);
or UO_1935 (O_1935,N_29943,N_29751);
nor UO_1936 (O_1936,N_29798,N_29738);
or UO_1937 (O_1937,N_29964,N_29758);
xor UO_1938 (O_1938,N_29927,N_29846);
xor UO_1939 (O_1939,N_29713,N_29990);
and UO_1940 (O_1940,N_29834,N_29915);
or UO_1941 (O_1941,N_29901,N_29904);
nor UO_1942 (O_1942,N_29841,N_29808);
nor UO_1943 (O_1943,N_29974,N_29971);
nand UO_1944 (O_1944,N_29867,N_29702);
xnor UO_1945 (O_1945,N_29827,N_29745);
and UO_1946 (O_1946,N_29849,N_29968);
nor UO_1947 (O_1947,N_29792,N_29911);
nand UO_1948 (O_1948,N_29764,N_29902);
nand UO_1949 (O_1949,N_29984,N_29728);
or UO_1950 (O_1950,N_29886,N_29713);
or UO_1951 (O_1951,N_29907,N_29781);
nand UO_1952 (O_1952,N_29760,N_29929);
or UO_1953 (O_1953,N_29814,N_29929);
nand UO_1954 (O_1954,N_29843,N_29787);
nor UO_1955 (O_1955,N_29905,N_29943);
xor UO_1956 (O_1956,N_29915,N_29809);
xor UO_1957 (O_1957,N_29784,N_29964);
and UO_1958 (O_1958,N_29756,N_29930);
nand UO_1959 (O_1959,N_29820,N_29909);
xnor UO_1960 (O_1960,N_29956,N_29773);
xnor UO_1961 (O_1961,N_29775,N_29991);
nor UO_1962 (O_1962,N_29972,N_29778);
nand UO_1963 (O_1963,N_29849,N_29935);
nor UO_1964 (O_1964,N_29956,N_29828);
and UO_1965 (O_1965,N_29899,N_29744);
nand UO_1966 (O_1966,N_29887,N_29964);
and UO_1967 (O_1967,N_29942,N_29789);
and UO_1968 (O_1968,N_29740,N_29813);
nand UO_1969 (O_1969,N_29824,N_29897);
nand UO_1970 (O_1970,N_29909,N_29794);
xnor UO_1971 (O_1971,N_29992,N_29957);
or UO_1972 (O_1972,N_29703,N_29889);
and UO_1973 (O_1973,N_29901,N_29756);
and UO_1974 (O_1974,N_29917,N_29839);
nand UO_1975 (O_1975,N_29708,N_29759);
nand UO_1976 (O_1976,N_29947,N_29718);
and UO_1977 (O_1977,N_29817,N_29792);
nand UO_1978 (O_1978,N_29704,N_29812);
xnor UO_1979 (O_1979,N_29862,N_29936);
and UO_1980 (O_1980,N_29779,N_29726);
xnor UO_1981 (O_1981,N_29764,N_29969);
nor UO_1982 (O_1982,N_29849,N_29885);
or UO_1983 (O_1983,N_29775,N_29829);
or UO_1984 (O_1984,N_29859,N_29722);
or UO_1985 (O_1985,N_29952,N_29922);
nand UO_1986 (O_1986,N_29707,N_29831);
xnor UO_1987 (O_1987,N_29704,N_29963);
nor UO_1988 (O_1988,N_29983,N_29923);
nand UO_1989 (O_1989,N_29765,N_29851);
nand UO_1990 (O_1990,N_29855,N_29757);
nor UO_1991 (O_1991,N_29827,N_29895);
nand UO_1992 (O_1992,N_29824,N_29856);
nor UO_1993 (O_1993,N_29771,N_29816);
and UO_1994 (O_1994,N_29786,N_29792);
xnor UO_1995 (O_1995,N_29937,N_29815);
nor UO_1996 (O_1996,N_29731,N_29775);
xnor UO_1997 (O_1997,N_29828,N_29914);
and UO_1998 (O_1998,N_29891,N_29828);
and UO_1999 (O_1999,N_29777,N_29715);
nand UO_2000 (O_2000,N_29732,N_29701);
nor UO_2001 (O_2001,N_29859,N_29863);
and UO_2002 (O_2002,N_29903,N_29714);
nor UO_2003 (O_2003,N_29747,N_29760);
xnor UO_2004 (O_2004,N_29778,N_29932);
xor UO_2005 (O_2005,N_29851,N_29920);
nand UO_2006 (O_2006,N_29813,N_29853);
xnor UO_2007 (O_2007,N_29940,N_29860);
or UO_2008 (O_2008,N_29752,N_29808);
nand UO_2009 (O_2009,N_29742,N_29737);
xnor UO_2010 (O_2010,N_29834,N_29764);
or UO_2011 (O_2011,N_29712,N_29902);
xor UO_2012 (O_2012,N_29966,N_29741);
nor UO_2013 (O_2013,N_29926,N_29849);
xor UO_2014 (O_2014,N_29798,N_29783);
or UO_2015 (O_2015,N_29982,N_29796);
or UO_2016 (O_2016,N_29961,N_29875);
xor UO_2017 (O_2017,N_29813,N_29979);
nor UO_2018 (O_2018,N_29708,N_29949);
and UO_2019 (O_2019,N_29952,N_29911);
and UO_2020 (O_2020,N_29991,N_29731);
and UO_2021 (O_2021,N_29980,N_29850);
and UO_2022 (O_2022,N_29749,N_29769);
or UO_2023 (O_2023,N_29827,N_29752);
or UO_2024 (O_2024,N_29989,N_29851);
nor UO_2025 (O_2025,N_29972,N_29731);
and UO_2026 (O_2026,N_29760,N_29820);
nor UO_2027 (O_2027,N_29879,N_29852);
nor UO_2028 (O_2028,N_29760,N_29941);
nand UO_2029 (O_2029,N_29848,N_29822);
nand UO_2030 (O_2030,N_29844,N_29961);
nor UO_2031 (O_2031,N_29816,N_29868);
and UO_2032 (O_2032,N_29774,N_29824);
and UO_2033 (O_2033,N_29701,N_29835);
or UO_2034 (O_2034,N_29708,N_29778);
and UO_2035 (O_2035,N_29950,N_29723);
or UO_2036 (O_2036,N_29774,N_29991);
nand UO_2037 (O_2037,N_29964,N_29811);
or UO_2038 (O_2038,N_29919,N_29905);
nor UO_2039 (O_2039,N_29714,N_29745);
and UO_2040 (O_2040,N_29768,N_29851);
nor UO_2041 (O_2041,N_29979,N_29917);
xnor UO_2042 (O_2042,N_29820,N_29873);
or UO_2043 (O_2043,N_29849,N_29985);
xnor UO_2044 (O_2044,N_29732,N_29790);
or UO_2045 (O_2045,N_29962,N_29723);
and UO_2046 (O_2046,N_29830,N_29827);
nor UO_2047 (O_2047,N_29805,N_29908);
nor UO_2048 (O_2048,N_29849,N_29995);
or UO_2049 (O_2049,N_29968,N_29707);
nor UO_2050 (O_2050,N_29998,N_29867);
nor UO_2051 (O_2051,N_29744,N_29701);
nand UO_2052 (O_2052,N_29774,N_29776);
nand UO_2053 (O_2053,N_29963,N_29733);
nand UO_2054 (O_2054,N_29805,N_29958);
or UO_2055 (O_2055,N_29788,N_29923);
nand UO_2056 (O_2056,N_29896,N_29760);
nor UO_2057 (O_2057,N_29907,N_29975);
or UO_2058 (O_2058,N_29995,N_29771);
xnor UO_2059 (O_2059,N_29894,N_29758);
or UO_2060 (O_2060,N_29755,N_29808);
nor UO_2061 (O_2061,N_29983,N_29793);
xor UO_2062 (O_2062,N_29749,N_29896);
or UO_2063 (O_2063,N_29969,N_29765);
nor UO_2064 (O_2064,N_29953,N_29748);
nand UO_2065 (O_2065,N_29916,N_29777);
nor UO_2066 (O_2066,N_29963,N_29829);
and UO_2067 (O_2067,N_29783,N_29998);
nor UO_2068 (O_2068,N_29714,N_29805);
xor UO_2069 (O_2069,N_29838,N_29839);
nand UO_2070 (O_2070,N_29841,N_29735);
xor UO_2071 (O_2071,N_29794,N_29765);
nor UO_2072 (O_2072,N_29900,N_29820);
and UO_2073 (O_2073,N_29808,N_29759);
xor UO_2074 (O_2074,N_29859,N_29911);
and UO_2075 (O_2075,N_29857,N_29714);
and UO_2076 (O_2076,N_29970,N_29814);
and UO_2077 (O_2077,N_29735,N_29890);
nor UO_2078 (O_2078,N_29818,N_29853);
and UO_2079 (O_2079,N_29878,N_29973);
xor UO_2080 (O_2080,N_29997,N_29803);
xnor UO_2081 (O_2081,N_29863,N_29940);
nor UO_2082 (O_2082,N_29933,N_29720);
nand UO_2083 (O_2083,N_29980,N_29835);
nand UO_2084 (O_2084,N_29700,N_29972);
nand UO_2085 (O_2085,N_29989,N_29806);
nor UO_2086 (O_2086,N_29961,N_29881);
nor UO_2087 (O_2087,N_29912,N_29799);
nand UO_2088 (O_2088,N_29832,N_29988);
nand UO_2089 (O_2089,N_29818,N_29888);
xnor UO_2090 (O_2090,N_29742,N_29855);
or UO_2091 (O_2091,N_29945,N_29765);
nor UO_2092 (O_2092,N_29745,N_29723);
or UO_2093 (O_2093,N_29916,N_29939);
and UO_2094 (O_2094,N_29859,N_29806);
nor UO_2095 (O_2095,N_29931,N_29700);
xnor UO_2096 (O_2096,N_29980,N_29822);
nand UO_2097 (O_2097,N_29718,N_29894);
nand UO_2098 (O_2098,N_29898,N_29708);
xnor UO_2099 (O_2099,N_29809,N_29749);
nor UO_2100 (O_2100,N_29810,N_29968);
nand UO_2101 (O_2101,N_29802,N_29999);
nor UO_2102 (O_2102,N_29979,N_29891);
nor UO_2103 (O_2103,N_29948,N_29924);
xor UO_2104 (O_2104,N_29731,N_29848);
and UO_2105 (O_2105,N_29771,N_29799);
xor UO_2106 (O_2106,N_29702,N_29906);
nor UO_2107 (O_2107,N_29713,N_29716);
nor UO_2108 (O_2108,N_29742,N_29927);
nand UO_2109 (O_2109,N_29728,N_29902);
and UO_2110 (O_2110,N_29957,N_29864);
xnor UO_2111 (O_2111,N_29808,N_29830);
nand UO_2112 (O_2112,N_29975,N_29779);
and UO_2113 (O_2113,N_29997,N_29953);
and UO_2114 (O_2114,N_29896,N_29948);
or UO_2115 (O_2115,N_29740,N_29926);
or UO_2116 (O_2116,N_29906,N_29811);
xnor UO_2117 (O_2117,N_29736,N_29888);
and UO_2118 (O_2118,N_29771,N_29828);
and UO_2119 (O_2119,N_29701,N_29951);
nand UO_2120 (O_2120,N_29769,N_29871);
or UO_2121 (O_2121,N_29737,N_29792);
nor UO_2122 (O_2122,N_29941,N_29920);
nand UO_2123 (O_2123,N_29989,N_29788);
and UO_2124 (O_2124,N_29793,N_29792);
and UO_2125 (O_2125,N_29967,N_29720);
nand UO_2126 (O_2126,N_29986,N_29872);
xor UO_2127 (O_2127,N_29729,N_29826);
and UO_2128 (O_2128,N_29827,N_29821);
or UO_2129 (O_2129,N_29873,N_29792);
and UO_2130 (O_2130,N_29956,N_29964);
or UO_2131 (O_2131,N_29967,N_29942);
xnor UO_2132 (O_2132,N_29910,N_29793);
xor UO_2133 (O_2133,N_29819,N_29898);
or UO_2134 (O_2134,N_29796,N_29792);
or UO_2135 (O_2135,N_29931,N_29724);
nor UO_2136 (O_2136,N_29716,N_29710);
and UO_2137 (O_2137,N_29983,N_29986);
nand UO_2138 (O_2138,N_29993,N_29985);
and UO_2139 (O_2139,N_29718,N_29790);
and UO_2140 (O_2140,N_29985,N_29889);
and UO_2141 (O_2141,N_29812,N_29956);
and UO_2142 (O_2142,N_29835,N_29882);
or UO_2143 (O_2143,N_29863,N_29965);
nand UO_2144 (O_2144,N_29822,N_29851);
or UO_2145 (O_2145,N_29978,N_29942);
and UO_2146 (O_2146,N_29984,N_29874);
or UO_2147 (O_2147,N_29996,N_29721);
nand UO_2148 (O_2148,N_29968,N_29793);
nor UO_2149 (O_2149,N_29791,N_29858);
xnor UO_2150 (O_2150,N_29927,N_29832);
or UO_2151 (O_2151,N_29747,N_29895);
xor UO_2152 (O_2152,N_29923,N_29724);
and UO_2153 (O_2153,N_29955,N_29763);
xor UO_2154 (O_2154,N_29712,N_29928);
nand UO_2155 (O_2155,N_29981,N_29987);
xor UO_2156 (O_2156,N_29981,N_29726);
or UO_2157 (O_2157,N_29804,N_29899);
nor UO_2158 (O_2158,N_29984,N_29972);
nand UO_2159 (O_2159,N_29768,N_29850);
nor UO_2160 (O_2160,N_29852,N_29849);
nor UO_2161 (O_2161,N_29721,N_29729);
and UO_2162 (O_2162,N_29713,N_29933);
and UO_2163 (O_2163,N_29870,N_29760);
nor UO_2164 (O_2164,N_29820,N_29844);
or UO_2165 (O_2165,N_29952,N_29717);
xor UO_2166 (O_2166,N_29973,N_29864);
nor UO_2167 (O_2167,N_29940,N_29944);
nand UO_2168 (O_2168,N_29804,N_29898);
or UO_2169 (O_2169,N_29895,N_29999);
xnor UO_2170 (O_2170,N_29906,N_29816);
or UO_2171 (O_2171,N_29883,N_29753);
nand UO_2172 (O_2172,N_29977,N_29740);
and UO_2173 (O_2173,N_29909,N_29867);
or UO_2174 (O_2174,N_29850,N_29958);
xor UO_2175 (O_2175,N_29704,N_29919);
nand UO_2176 (O_2176,N_29785,N_29743);
nor UO_2177 (O_2177,N_29925,N_29778);
nor UO_2178 (O_2178,N_29721,N_29984);
nand UO_2179 (O_2179,N_29755,N_29975);
nand UO_2180 (O_2180,N_29994,N_29715);
or UO_2181 (O_2181,N_29972,N_29842);
or UO_2182 (O_2182,N_29739,N_29706);
nand UO_2183 (O_2183,N_29740,N_29908);
nor UO_2184 (O_2184,N_29868,N_29838);
or UO_2185 (O_2185,N_29826,N_29815);
xor UO_2186 (O_2186,N_29711,N_29856);
or UO_2187 (O_2187,N_29741,N_29802);
nand UO_2188 (O_2188,N_29981,N_29727);
and UO_2189 (O_2189,N_29894,N_29935);
nand UO_2190 (O_2190,N_29967,N_29754);
nor UO_2191 (O_2191,N_29780,N_29844);
and UO_2192 (O_2192,N_29862,N_29779);
or UO_2193 (O_2193,N_29929,N_29758);
or UO_2194 (O_2194,N_29873,N_29881);
nor UO_2195 (O_2195,N_29874,N_29743);
nand UO_2196 (O_2196,N_29854,N_29764);
nand UO_2197 (O_2197,N_29878,N_29894);
xor UO_2198 (O_2198,N_29989,N_29830);
xor UO_2199 (O_2199,N_29786,N_29740);
and UO_2200 (O_2200,N_29709,N_29834);
and UO_2201 (O_2201,N_29943,N_29733);
nand UO_2202 (O_2202,N_29741,N_29891);
nand UO_2203 (O_2203,N_29823,N_29803);
and UO_2204 (O_2204,N_29717,N_29780);
or UO_2205 (O_2205,N_29875,N_29730);
nor UO_2206 (O_2206,N_29835,N_29817);
xnor UO_2207 (O_2207,N_29719,N_29716);
nand UO_2208 (O_2208,N_29862,N_29889);
nor UO_2209 (O_2209,N_29989,N_29769);
and UO_2210 (O_2210,N_29760,N_29981);
and UO_2211 (O_2211,N_29858,N_29823);
nor UO_2212 (O_2212,N_29704,N_29810);
xnor UO_2213 (O_2213,N_29939,N_29751);
xnor UO_2214 (O_2214,N_29818,N_29871);
or UO_2215 (O_2215,N_29928,N_29924);
and UO_2216 (O_2216,N_29713,N_29797);
and UO_2217 (O_2217,N_29787,N_29831);
and UO_2218 (O_2218,N_29933,N_29953);
xnor UO_2219 (O_2219,N_29783,N_29920);
nand UO_2220 (O_2220,N_29709,N_29860);
or UO_2221 (O_2221,N_29809,N_29743);
and UO_2222 (O_2222,N_29792,N_29979);
xor UO_2223 (O_2223,N_29748,N_29957);
and UO_2224 (O_2224,N_29891,N_29924);
nor UO_2225 (O_2225,N_29835,N_29984);
or UO_2226 (O_2226,N_29842,N_29899);
xnor UO_2227 (O_2227,N_29867,N_29799);
xor UO_2228 (O_2228,N_29894,N_29921);
or UO_2229 (O_2229,N_29869,N_29938);
nand UO_2230 (O_2230,N_29869,N_29731);
nand UO_2231 (O_2231,N_29727,N_29716);
nand UO_2232 (O_2232,N_29907,N_29911);
nand UO_2233 (O_2233,N_29719,N_29761);
nor UO_2234 (O_2234,N_29818,N_29725);
nand UO_2235 (O_2235,N_29959,N_29838);
and UO_2236 (O_2236,N_29767,N_29822);
nand UO_2237 (O_2237,N_29782,N_29740);
nand UO_2238 (O_2238,N_29889,N_29947);
nor UO_2239 (O_2239,N_29950,N_29827);
and UO_2240 (O_2240,N_29845,N_29788);
or UO_2241 (O_2241,N_29717,N_29778);
nand UO_2242 (O_2242,N_29754,N_29825);
nand UO_2243 (O_2243,N_29861,N_29978);
nand UO_2244 (O_2244,N_29964,N_29950);
nand UO_2245 (O_2245,N_29829,N_29876);
nand UO_2246 (O_2246,N_29721,N_29926);
xor UO_2247 (O_2247,N_29803,N_29862);
and UO_2248 (O_2248,N_29956,N_29795);
or UO_2249 (O_2249,N_29980,N_29766);
xor UO_2250 (O_2250,N_29906,N_29707);
nand UO_2251 (O_2251,N_29809,N_29856);
xnor UO_2252 (O_2252,N_29989,N_29777);
xor UO_2253 (O_2253,N_29822,N_29934);
nor UO_2254 (O_2254,N_29808,N_29894);
and UO_2255 (O_2255,N_29750,N_29941);
nor UO_2256 (O_2256,N_29987,N_29853);
and UO_2257 (O_2257,N_29901,N_29891);
xor UO_2258 (O_2258,N_29815,N_29766);
or UO_2259 (O_2259,N_29705,N_29837);
and UO_2260 (O_2260,N_29886,N_29819);
xor UO_2261 (O_2261,N_29753,N_29744);
nand UO_2262 (O_2262,N_29950,N_29700);
or UO_2263 (O_2263,N_29898,N_29755);
nor UO_2264 (O_2264,N_29956,N_29713);
and UO_2265 (O_2265,N_29822,N_29995);
or UO_2266 (O_2266,N_29870,N_29727);
xnor UO_2267 (O_2267,N_29750,N_29703);
xor UO_2268 (O_2268,N_29991,N_29926);
nor UO_2269 (O_2269,N_29773,N_29746);
or UO_2270 (O_2270,N_29783,N_29968);
or UO_2271 (O_2271,N_29729,N_29710);
nor UO_2272 (O_2272,N_29888,N_29874);
or UO_2273 (O_2273,N_29817,N_29785);
xnor UO_2274 (O_2274,N_29920,N_29806);
and UO_2275 (O_2275,N_29782,N_29871);
xnor UO_2276 (O_2276,N_29994,N_29822);
and UO_2277 (O_2277,N_29852,N_29810);
nor UO_2278 (O_2278,N_29768,N_29810);
nor UO_2279 (O_2279,N_29843,N_29818);
nor UO_2280 (O_2280,N_29937,N_29968);
nor UO_2281 (O_2281,N_29812,N_29821);
or UO_2282 (O_2282,N_29795,N_29964);
xnor UO_2283 (O_2283,N_29941,N_29770);
and UO_2284 (O_2284,N_29991,N_29870);
xor UO_2285 (O_2285,N_29722,N_29709);
and UO_2286 (O_2286,N_29971,N_29987);
nand UO_2287 (O_2287,N_29858,N_29914);
nand UO_2288 (O_2288,N_29915,N_29912);
and UO_2289 (O_2289,N_29957,N_29746);
nand UO_2290 (O_2290,N_29807,N_29783);
nor UO_2291 (O_2291,N_29747,N_29824);
nor UO_2292 (O_2292,N_29785,N_29713);
and UO_2293 (O_2293,N_29765,N_29881);
nor UO_2294 (O_2294,N_29922,N_29811);
and UO_2295 (O_2295,N_29904,N_29979);
or UO_2296 (O_2296,N_29743,N_29918);
and UO_2297 (O_2297,N_29801,N_29880);
nor UO_2298 (O_2298,N_29890,N_29921);
nand UO_2299 (O_2299,N_29964,N_29988);
or UO_2300 (O_2300,N_29942,N_29888);
nor UO_2301 (O_2301,N_29885,N_29779);
xnor UO_2302 (O_2302,N_29746,N_29938);
xnor UO_2303 (O_2303,N_29750,N_29766);
nand UO_2304 (O_2304,N_29925,N_29912);
nor UO_2305 (O_2305,N_29950,N_29780);
xnor UO_2306 (O_2306,N_29888,N_29981);
xor UO_2307 (O_2307,N_29803,N_29868);
xnor UO_2308 (O_2308,N_29766,N_29798);
nand UO_2309 (O_2309,N_29795,N_29957);
xnor UO_2310 (O_2310,N_29977,N_29729);
and UO_2311 (O_2311,N_29866,N_29926);
and UO_2312 (O_2312,N_29928,N_29872);
or UO_2313 (O_2313,N_29771,N_29991);
xnor UO_2314 (O_2314,N_29721,N_29815);
xnor UO_2315 (O_2315,N_29807,N_29792);
and UO_2316 (O_2316,N_29755,N_29903);
nand UO_2317 (O_2317,N_29945,N_29815);
nor UO_2318 (O_2318,N_29756,N_29925);
nand UO_2319 (O_2319,N_29990,N_29795);
or UO_2320 (O_2320,N_29729,N_29751);
or UO_2321 (O_2321,N_29964,N_29938);
and UO_2322 (O_2322,N_29991,N_29811);
and UO_2323 (O_2323,N_29704,N_29962);
nor UO_2324 (O_2324,N_29766,N_29831);
xor UO_2325 (O_2325,N_29708,N_29830);
xor UO_2326 (O_2326,N_29993,N_29874);
nand UO_2327 (O_2327,N_29811,N_29775);
and UO_2328 (O_2328,N_29862,N_29857);
and UO_2329 (O_2329,N_29741,N_29959);
and UO_2330 (O_2330,N_29879,N_29871);
and UO_2331 (O_2331,N_29881,N_29891);
nand UO_2332 (O_2332,N_29853,N_29821);
xnor UO_2333 (O_2333,N_29812,N_29742);
or UO_2334 (O_2334,N_29959,N_29707);
nor UO_2335 (O_2335,N_29784,N_29727);
nor UO_2336 (O_2336,N_29796,N_29962);
nor UO_2337 (O_2337,N_29933,N_29860);
and UO_2338 (O_2338,N_29963,N_29984);
nand UO_2339 (O_2339,N_29719,N_29816);
nand UO_2340 (O_2340,N_29808,N_29702);
xor UO_2341 (O_2341,N_29745,N_29998);
nand UO_2342 (O_2342,N_29840,N_29949);
xor UO_2343 (O_2343,N_29952,N_29790);
nand UO_2344 (O_2344,N_29870,N_29762);
xnor UO_2345 (O_2345,N_29908,N_29787);
xnor UO_2346 (O_2346,N_29847,N_29870);
nand UO_2347 (O_2347,N_29839,N_29732);
nor UO_2348 (O_2348,N_29743,N_29701);
nor UO_2349 (O_2349,N_29978,N_29720);
and UO_2350 (O_2350,N_29941,N_29977);
and UO_2351 (O_2351,N_29713,N_29842);
xnor UO_2352 (O_2352,N_29769,N_29745);
or UO_2353 (O_2353,N_29753,N_29996);
nor UO_2354 (O_2354,N_29975,N_29840);
xor UO_2355 (O_2355,N_29757,N_29797);
and UO_2356 (O_2356,N_29751,N_29954);
nand UO_2357 (O_2357,N_29796,N_29790);
xor UO_2358 (O_2358,N_29939,N_29961);
or UO_2359 (O_2359,N_29907,N_29982);
nand UO_2360 (O_2360,N_29768,N_29991);
and UO_2361 (O_2361,N_29745,N_29953);
and UO_2362 (O_2362,N_29708,N_29965);
or UO_2363 (O_2363,N_29799,N_29831);
nand UO_2364 (O_2364,N_29823,N_29847);
nor UO_2365 (O_2365,N_29984,N_29870);
or UO_2366 (O_2366,N_29896,N_29890);
or UO_2367 (O_2367,N_29935,N_29967);
xnor UO_2368 (O_2368,N_29882,N_29828);
xnor UO_2369 (O_2369,N_29980,N_29918);
or UO_2370 (O_2370,N_29853,N_29960);
or UO_2371 (O_2371,N_29781,N_29920);
and UO_2372 (O_2372,N_29998,N_29934);
or UO_2373 (O_2373,N_29980,N_29826);
nor UO_2374 (O_2374,N_29956,N_29866);
and UO_2375 (O_2375,N_29988,N_29891);
and UO_2376 (O_2376,N_29811,N_29749);
and UO_2377 (O_2377,N_29919,N_29890);
nand UO_2378 (O_2378,N_29786,N_29704);
or UO_2379 (O_2379,N_29703,N_29776);
nor UO_2380 (O_2380,N_29723,N_29834);
or UO_2381 (O_2381,N_29815,N_29728);
xnor UO_2382 (O_2382,N_29952,N_29808);
and UO_2383 (O_2383,N_29833,N_29904);
xor UO_2384 (O_2384,N_29896,N_29756);
and UO_2385 (O_2385,N_29794,N_29743);
nor UO_2386 (O_2386,N_29864,N_29854);
nor UO_2387 (O_2387,N_29751,N_29942);
nor UO_2388 (O_2388,N_29930,N_29898);
nor UO_2389 (O_2389,N_29784,N_29714);
nand UO_2390 (O_2390,N_29852,N_29707);
xor UO_2391 (O_2391,N_29839,N_29995);
xor UO_2392 (O_2392,N_29775,N_29760);
and UO_2393 (O_2393,N_29929,N_29839);
nor UO_2394 (O_2394,N_29702,N_29740);
xnor UO_2395 (O_2395,N_29956,N_29909);
or UO_2396 (O_2396,N_29715,N_29911);
nand UO_2397 (O_2397,N_29837,N_29998);
nor UO_2398 (O_2398,N_29925,N_29770);
nor UO_2399 (O_2399,N_29802,N_29927);
xnor UO_2400 (O_2400,N_29803,N_29853);
nor UO_2401 (O_2401,N_29985,N_29965);
and UO_2402 (O_2402,N_29759,N_29945);
and UO_2403 (O_2403,N_29702,N_29705);
xnor UO_2404 (O_2404,N_29761,N_29953);
nand UO_2405 (O_2405,N_29944,N_29974);
and UO_2406 (O_2406,N_29798,N_29880);
and UO_2407 (O_2407,N_29735,N_29737);
nor UO_2408 (O_2408,N_29780,N_29927);
or UO_2409 (O_2409,N_29966,N_29974);
nor UO_2410 (O_2410,N_29760,N_29763);
nor UO_2411 (O_2411,N_29841,N_29782);
or UO_2412 (O_2412,N_29949,N_29926);
xnor UO_2413 (O_2413,N_29795,N_29897);
and UO_2414 (O_2414,N_29947,N_29713);
nor UO_2415 (O_2415,N_29957,N_29798);
xnor UO_2416 (O_2416,N_29956,N_29842);
xor UO_2417 (O_2417,N_29997,N_29944);
or UO_2418 (O_2418,N_29854,N_29940);
and UO_2419 (O_2419,N_29753,N_29947);
xnor UO_2420 (O_2420,N_29983,N_29702);
nand UO_2421 (O_2421,N_29755,N_29746);
nand UO_2422 (O_2422,N_29721,N_29703);
nand UO_2423 (O_2423,N_29864,N_29954);
nor UO_2424 (O_2424,N_29768,N_29713);
or UO_2425 (O_2425,N_29880,N_29744);
nor UO_2426 (O_2426,N_29755,N_29727);
nand UO_2427 (O_2427,N_29912,N_29732);
xor UO_2428 (O_2428,N_29801,N_29890);
and UO_2429 (O_2429,N_29837,N_29800);
and UO_2430 (O_2430,N_29750,N_29944);
nor UO_2431 (O_2431,N_29945,N_29851);
nand UO_2432 (O_2432,N_29785,N_29792);
and UO_2433 (O_2433,N_29981,N_29947);
xnor UO_2434 (O_2434,N_29734,N_29825);
nor UO_2435 (O_2435,N_29905,N_29950);
and UO_2436 (O_2436,N_29932,N_29865);
nor UO_2437 (O_2437,N_29938,N_29759);
and UO_2438 (O_2438,N_29759,N_29811);
nand UO_2439 (O_2439,N_29931,N_29893);
nand UO_2440 (O_2440,N_29981,N_29854);
and UO_2441 (O_2441,N_29921,N_29732);
and UO_2442 (O_2442,N_29772,N_29856);
or UO_2443 (O_2443,N_29850,N_29871);
xnor UO_2444 (O_2444,N_29875,N_29765);
or UO_2445 (O_2445,N_29761,N_29847);
nor UO_2446 (O_2446,N_29950,N_29902);
nor UO_2447 (O_2447,N_29807,N_29860);
nand UO_2448 (O_2448,N_29911,N_29906);
or UO_2449 (O_2449,N_29716,N_29831);
nor UO_2450 (O_2450,N_29963,N_29869);
xor UO_2451 (O_2451,N_29983,N_29949);
nand UO_2452 (O_2452,N_29799,N_29942);
or UO_2453 (O_2453,N_29990,N_29956);
xnor UO_2454 (O_2454,N_29860,N_29742);
xnor UO_2455 (O_2455,N_29897,N_29971);
or UO_2456 (O_2456,N_29744,N_29767);
xor UO_2457 (O_2457,N_29900,N_29833);
nand UO_2458 (O_2458,N_29965,N_29971);
and UO_2459 (O_2459,N_29737,N_29800);
xnor UO_2460 (O_2460,N_29823,N_29707);
nand UO_2461 (O_2461,N_29945,N_29723);
and UO_2462 (O_2462,N_29980,N_29943);
or UO_2463 (O_2463,N_29859,N_29943);
and UO_2464 (O_2464,N_29736,N_29706);
or UO_2465 (O_2465,N_29997,N_29908);
and UO_2466 (O_2466,N_29898,N_29877);
xor UO_2467 (O_2467,N_29927,N_29912);
nor UO_2468 (O_2468,N_29761,N_29849);
nand UO_2469 (O_2469,N_29870,N_29935);
and UO_2470 (O_2470,N_29764,N_29967);
and UO_2471 (O_2471,N_29985,N_29930);
or UO_2472 (O_2472,N_29713,N_29852);
xor UO_2473 (O_2473,N_29983,N_29832);
nor UO_2474 (O_2474,N_29754,N_29971);
xnor UO_2475 (O_2475,N_29928,N_29758);
xnor UO_2476 (O_2476,N_29797,N_29737);
nand UO_2477 (O_2477,N_29865,N_29854);
xnor UO_2478 (O_2478,N_29921,N_29948);
xnor UO_2479 (O_2479,N_29707,N_29882);
and UO_2480 (O_2480,N_29793,N_29762);
nor UO_2481 (O_2481,N_29714,N_29964);
or UO_2482 (O_2482,N_29734,N_29730);
and UO_2483 (O_2483,N_29984,N_29930);
nand UO_2484 (O_2484,N_29882,N_29954);
or UO_2485 (O_2485,N_29884,N_29984);
nand UO_2486 (O_2486,N_29933,N_29831);
or UO_2487 (O_2487,N_29934,N_29735);
nand UO_2488 (O_2488,N_29701,N_29771);
nor UO_2489 (O_2489,N_29744,N_29981);
or UO_2490 (O_2490,N_29792,N_29881);
xor UO_2491 (O_2491,N_29903,N_29822);
nor UO_2492 (O_2492,N_29767,N_29702);
or UO_2493 (O_2493,N_29894,N_29730);
nand UO_2494 (O_2494,N_29969,N_29887);
or UO_2495 (O_2495,N_29980,N_29996);
or UO_2496 (O_2496,N_29774,N_29878);
nor UO_2497 (O_2497,N_29780,N_29729);
and UO_2498 (O_2498,N_29779,N_29886);
and UO_2499 (O_2499,N_29987,N_29744);
nand UO_2500 (O_2500,N_29908,N_29851);
nand UO_2501 (O_2501,N_29915,N_29750);
or UO_2502 (O_2502,N_29833,N_29948);
or UO_2503 (O_2503,N_29700,N_29827);
nor UO_2504 (O_2504,N_29848,N_29851);
and UO_2505 (O_2505,N_29831,N_29751);
and UO_2506 (O_2506,N_29784,N_29810);
xnor UO_2507 (O_2507,N_29932,N_29953);
or UO_2508 (O_2508,N_29824,N_29942);
nand UO_2509 (O_2509,N_29923,N_29912);
nor UO_2510 (O_2510,N_29964,N_29886);
and UO_2511 (O_2511,N_29956,N_29765);
nand UO_2512 (O_2512,N_29826,N_29708);
nor UO_2513 (O_2513,N_29731,N_29734);
xnor UO_2514 (O_2514,N_29703,N_29907);
or UO_2515 (O_2515,N_29778,N_29819);
nor UO_2516 (O_2516,N_29921,N_29841);
nand UO_2517 (O_2517,N_29800,N_29774);
or UO_2518 (O_2518,N_29938,N_29702);
nor UO_2519 (O_2519,N_29924,N_29971);
xnor UO_2520 (O_2520,N_29837,N_29943);
or UO_2521 (O_2521,N_29763,N_29839);
xor UO_2522 (O_2522,N_29745,N_29967);
and UO_2523 (O_2523,N_29841,N_29998);
xor UO_2524 (O_2524,N_29927,N_29700);
and UO_2525 (O_2525,N_29894,N_29864);
xnor UO_2526 (O_2526,N_29873,N_29805);
or UO_2527 (O_2527,N_29910,N_29709);
and UO_2528 (O_2528,N_29729,N_29814);
and UO_2529 (O_2529,N_29912,N_29934);
nor UO_2530 (O_2530,N_29723,N_29864);
nand UO_2531 (O_2531,N_29712,N_29750);
and UO_2532 (O_2532,N_29925,N_29871);
nor UO_2533 (O_2533,N_29821,N_29710);
and UO_2534 (O_2534,N_29822,N_29722);
and UO_2535 (O_2535,N_29948,N_29953);
nand UO_2536 (O_2536,N_29967,N_29710);
or UO_2537 (O_2537,N_29960,N_29977);
nand UO_2538 (O_2538,N_29968,N_29915);
nand UO_2539 (O_2539,N_29826,N_29941);
or UO_2540 (O_2540,N_29906,N_29749);
nor UO_2541 (O_2541,N_29738,N_29936);
nor UO_2542 (O_2542,N_29747,N_29849);
nand UO_2543 (O_2543,N_29900,N_29705);
xor UO_2544 (O_2544,N_29843,N_29997);
nand UO_2545 (O_2545,N_29752,N_29852);
and UO_2546 (O_2546,N_29863,N_29906);
nand UO_2547 (O_2547,N_29895,N_29964);
xnor UO_2548 (O_2548,N_29840,N_29772);
or UO_2549 (O_2549,N_29804,N_29977);
nor UO_2550 (O_2550,N_29958,N_29880);
and UO_2551 (O_2551,N_29861,N_29986);
nand UO_2552 (O_2552,N_29834,N_29923);
nor UO_2553 (O_2553,N_29847,N_29873);
xnor UO_2554 (O_2554,N_29951,N_29733);
nand UO_2555 (O_2555,N_29735,N_29953);
nor UO_2556 (O_2556,N_29750,N_29829);
nor UO_2557 (O_2557,N_29885,N_29955);
nor UO_2558 (O_2558,N_29825,N_29788);
nor UO_2559 (O_2559,N_29798,N_29927);
xor UO_2560 (O_2560,N_29744,N_29986);
xor UO_2561 (O_2561,N_29900,N_29993);
xor UO_2562 (O_2562,N_29906,N_29900);
nor UO_2563 (O_2563,N_29871,N_29931);
nor UO_2564 (O_2564,N_29866,N_29949);
nand UO_2565 (O_2565,N_29936,N_29865);
xnor UO_2566 (O_2566,N_29760,N_29737);
and UO_2567 (O_2567,N_29740,N_29914);
nor UO_2568 (O_2568,N_29993,N_29735);
or UO_2569 (O_2569,N_29728,N_29801);
nand UO_2570 (O_2570,N_29740,N_29784);
and UO_2571 (O_2571,N_29779,N_29958);
or UO_2572 (O_2572,N_29757,N_29982);
nor UO_2573 (O_2573,N_29773,N_29776);
and UO_2574 (O_2574,N_29949,N_29843);
and UO_2575 (O_2575,N_29747,N_29800);
or UO_2576 (O_2576,N_29955,N_29853);
and UO_2577 (O_2577,N_29969,N_29742);
xor UO_2578 (O_2578,N_29849,N_29811);
or UO_2579 (O_2579,N_29789,N_29806);
nand UO_2580 (O_2580,N_29779,N_29714);
nand UO_2581 (O_2581,N_29750,N_29924);
xnor UO_2582 (O_2582,N_29861,N_29717);
nor UO_2583 (O_2583,N_29923,N_29785);
xnor UO_2584 (O_2584,N_29866,N_29709);
and UO_2585 (O_2585,N_29818,N_29743);
or UO_2586 (O_2586,N_29755,N_29763);
xor UO_2587 (O_2587,N_29886,N_29834);
xor UO_2588 (O_2588,N_29929,N_29868);
and UO_2589 (O_2589,N_29899,N_29926);
nand UO_2590 (O_2590,N_29855,N_29833);
and UO_2591 (O_2591,N_29730,N_29994);
nor UO_2592 (O_2592,N_29717,N_29934);
nor UO_2593 (O_2593,N_29829,N_29812);
nand UO_2594 (O_2594,N_29949,N_29794);
or UO_2595 (O_2595,N_29984,N_29758);
and UO_2596 (O_2596,N_29765,N_29807);
or UO_2597 (O_2597,N_29834,N_29953);
and UO_2598 (O_2598,N_29867,N_29985);
and UO_2599 (O_2599,N_29973,N_29841);
and UO_2600 (O_2600,N_29913,N_29836);
xnor UO_2601 (O_2601,N_29804,N_29927);
xnor UO_2602 (O_2602,N_29790,N_29891);
nand UO_2603 (O_2603,N_29924,N_29887);
and UO_2604 (O_2604,N_29896,N_29985);
nand UO_2605 (O_2605,N_29787,N_29987);
or UO_2606 (O_2606,N_29906,N_29834);
xnor UO_2607 (O_2607,N_29701,N_29848);
xor UO_2608 (O_2608,N_29878,N_29735);
or UO_2609 (O_2609,N_29732,N_29793);
nand UO_2610 (O_2610,N_29783,N_29874);
and UO_2611 (O_2611,N_29811,N_29815);
and UO_2612 (O_2612,N_29924,N_29762);
nand UO_2613 (O_2613,N_29807,N_29831);
nor UO_2614 (O_2614,N_29976,N_29742);
and UO_2615 (O_2615,N_29842,N_29998);
or UO_2616 (O_2616,N_29949,N_29733);
and UO_2617 (O_2617,N_29885,N_29900);
and UO_2618 (O_2618,N_29838,N_29737);
xor UO_2619 (O_2619,N_29710,N_29778);
xor UO_2620 (O_2620,N_29756,N_29897);
and UO_2621 (O_2621,N_29896,N_29743);
nand UO_2622 (O_2622,N_29991,N_29896);
and UO_2623 (O_2623,N_29747,N_29946);
nor UO_2624 (O_2624,N_29921,N_29875);
and UO_2625 (O_2625,N_29770,N_29948);
xnor UO_2626 (O_2626,N_29886,N_29742);
nor UO_2627 (O_2627,N_29712,N_29796);
nand UO_2628 (O_2628,N_29900,N_29700);
nand UO_2629 (O_2629,N_29858,N_29899);
or UO_2630 (O_2630,N_29953,N_29829);
and UO_2631 (O_2631,N_29856,N_29895);
nor UO_2632 (O_2632,N_29991,N_29809);
nand UO_2633 (O_2633,N_29839,N_29705);
and UO_2634 (O_2634,N_29791,N_29757);
nand UO_2635 (O_2635,N_29799,N_29919);
nand UO_2636 (O_2636,N_29876,N_29774);
and UO_2637 (O_2637,N_29890,N_29980);
nor UO_2638 (O_2638,N_29897,N_29978);
nand UO_2639 (O_2639,N_29987,N_29745);
and UO_2640 (O_2640,N_29769,N_29831);
nor UO_2641 (O_2641,N_29732,N_29818);
xor UO_2642 (O_2642,N_29931,N_29843);
or UO_2643 (O_2643,N_29835,N_29857);
and UO_2644 (O_2644,N_29950,N_29992);
and UO_2645 (O_2645,N_29793,N_29978);
nand UO_2646 (O_2646,N_29807,N_29892);
or UO_2647 (O_2647,N_29932,N_29876);
nor UO_2648 (O_2648,N_29904,N_29814);
and UO_2649 (O_2649,N_29873,N_29808);
xor UO_2650 (O_2650,N_29885,N_29928);
xor UO_2651 (O_2651,N_29703,N_29899);
xor UO_2652 (O_2652,N_29727,N_29865);
or UO_2653 (O_2653,N_29728,N_29839);
nand UO_2654 (O_2654,N_29776,N_29891);
nand UO_2655 (O_2655,N_29872,N_29796);
and UO_2656 (O_2656,N_29775,N_29982);
or UO_2657 (O_2657,N_29993,N_29816);
or UO_2658 (O_2658,N_29831,N_29814);
and UO_2659 (O_2659,N_29880,N_29746);
nor UO_2660 (O_2660,N_29735,N_29970);
and UO_2661 (O_2661,N_29885,N_29968);
xor UO_2662 (O_2662,N_29936,N_29751);
nand UO_2663 (O_2663,N_29867,N_29918);
and UO_2664 (O_2664,N_29848,N_29785);
and UO_2665 (O_2665,N_29910,N_29710);
nand UO_2666 (O_2666,N_29745,N_29829);
or UO_2667 (O_2667,N_29807,N_29935);
xor UO_2668 (O_2668,N_29728,N_29727);
nor UO_2669 (O_2669,N_29779,N_29893);
xor UO_2670 (O_2670,N_29864,N_29947);
or UO_2671 (O_2671,N_29978,N_29738);
and UO_2672 (O_2672,N_29958,N_29794);
nor UO_2673 (O_2673,N_29787,N_29934);
and UO_2674 (O_2674,N_29882,N_29905);
and UO_2675 (O_2675,N_29795,N_29838);
nor UO_2676 (O_2676,N_29742,N_29961);
nor UO_2677 (O_2677,N_29921,N_29950);
and UO_2678 (O_2678,N_29751,N_29913);
xnor UO_2679 (O_2679,N_29979,N_29943);
nor UO_2680 (O_2680,N_29877,N_29884);
nand UO_2681 (O_2681,N_29710,N_29933);
and UO_2682 (O_2682,N_29807,N_29901);
and UO_2683 (O_2683,N_29852,N_29754);
and UO_2684 (O_2684,N_29721,N_29787);
and UO_2685 (O_2685,N_29876,N_29755);
nor UO_2686 (O_2686,N_29972,N_29991);
nand UO_2687 (O_2687,N_29986,N_29837);
xor UO_2688 (O_2688,N_29771,N_29973);
or UO_2689 (O_2689,N_29996,N_29789);
nor UO_2690 (O_2690,N_29754,N_29866);
xor UO_2691 (O_2691,N_29760,N_29951);
nand UO_2692 (O_2692,N_29810,N_29825);
or UO_2693 (O_2693,N_29982,N_29764);
nand UO_2694 (O_2694,N_29846,N_29824);
nand UO_2695 (O_2695,N_29972,N_29801);
and UO_2696 (O_2696,N_29778,N_29929);
and UO_2697 (O_2697,N_29978,N_29854);
nand UO_2698 (O_2698,N_29823,N_29855);
or UO_2699 (O_2699,N_29905,N_29812);
xor UO_2700 (O_2700,N_29925,N_29888);
or UO_2701 (O_2701,N_29839,N_29788);
nor UO_2702 (O_2702,N_29997,N_29906);
xnor UO_2703 (O_2703,N_29812,N_29866);
xor UO_2704 (O_2704,N_29775,N_29830);
nor UO_2705 (O_2705,N_29868,N_29704);
xnor UO_2706 (O_2706,N_29951,N_29927);
or UO_2707 (O_2707,N_29848,N_29920);
and UO_2708 (O_2708,N_29920,N_29965);
nor UO_2709 (O_2709,N_29884,N_29713);
and UO_2710 (O_2710,N_29954,N_29808);
nand UO_2711 (O_2711,N_29939,N_29872);
nor UO_2712 (O_2712,N_29790,N_29715);
and UO_2713 (O_2713,N_29817,N_29708);
nor UO_2714 (O_2714,N_29756,N_29965);
nand UO_2715 (O_2715,N_29996,N_29880);
xnor UO_2716 (O_2716,N_29705,N_29885);
or UO_2717 (O_2717,N_29700,N_29863);
xnor UO_2718 (O_2718,N_29852,N_29903);
xor UO_2719 (O_2719,N_29852,N_29963);
nor UO_2720 (O_2720,N_29998,N_29973);
and UO_2721 (O_2721,N_29777,N_29907);
xor UO_2722 (O_2722,N_29928,N_29707);
and UO_2723 (O_2723,N_29787,N_29827);
or UO_2724 (O_2724,N_29748,N_29754);
or UO_2725 (O_2725,N_29717,N_29957);
nand UO_2726 (O_2726,N_29892,N_29730);
nand UO_2727 (O_2727,N_29771,N_29770);
nand UO_2728 (O_2728,N_29889,N_29821);
xnor UO_2729 (O_2729,N_29906,N_29887);
nor UO_2730 (O_2730,N_29891,N_29809);
nor UO_2731 (O_2731,N_29799,N_29987);
nand UO_2732 (O_2732,N_29933,N_29984);
nor UO_2733 (O_2733,N_29952,N_29941);
and UO_2734 (O_2734,N_29746,N_29978);
and UO_2735 (O_2735,N_29986,N_29729);
xor UO_2736 (O_2736,N_29953,N_29861);
nor UO_2737 (O_2737,N_29905,N_29993);
or UO_2738 (O_2738,N_29755,N_29866);
xnor UO_2739 (O_2739,N_29809,N_29726);
or UO_2740 (O_2740,N_29759,N_29901);
and UO_2741 (O_2741,N_29985,N_29716);
xnor UO_2742 (O_2742,N_29980,N_29866);
nand UO_2743 (O_2743,N_29705,N_29996);
xnor UO_2744 (O_2744,N_29924,N_29873);
and UO_2745 (O_2745,N_29769,N_29784);
nand UO_2746 (O_2746,N_29836,N_29925);
nand UO_2747 (O_2747,N_29806,N_29967);
nand UO_2748 (O_2748,N_29885,N_29976);
and UO_2749 (O_2749,N_29720,N_29711);
nand UO_2750 (O_2750,N_29835,N_29898);
nor UO_2751 (O_2751,N_29714,N_29948);
nor UO_2752 (O_2752,N_29706,N_29761);
nor UO_2753 (O_2753,N_29935,N_29809);
or UO_2754 (O_2754,N_29750,N_29994);
and UO_2755 (O_2755,N_29951,N_29784);
and UO_2756 (O_2756,N_29731,N_29794);
xnor UO_2757 (O_2757,N_29804,N_29827);
or UO_2758 (O_2758,N_29981,N_29709);
or UO_2759 (O_2759,N_29802,N_29912);
nor UO_2760 (O_2760,N_29754,N_29768);
nand UO_2761 (O_2761,N_29986,N_29936);
and UO_2762 (O_2762,N_29743,N_29934);
xnor UO_2763 (O_2763,N_29833,N_29712);
nand UO_2764 (O_2764,N_29770,N_29844);
xor UO_2765 (O_2765,N_29759,N_29735);
nand UO_2766 (O_2766,N_29982,N_29839);
and UO_2767 (O_2767,N_29983,N_29822);
and UO_2768 (O_2768,N_29850,N_29720);
nand UO_2769 (O_2769,N_29951,N_29878);
nor UO_2770 (O_2770,N_29832,N_29935);
nor UO_2771 (O_2771,N_29762,N_29771);
nand UO_2772 (O_2772,N_29993,N_29978);
or UO_2773 (O_2773,N_29720,N_29749);
nand UO_2774 (O_2774,N_29961,N_29820);
nand UO_2775 (O_2775,N_29813,N_29962);
or UO_2776 (O_2776,N_29958,N_29967);
nor UO_2777 (O_2777,N_29770,N_29837);
and UO_2778 (O_2778,N_29882,N_29898);
nor UO_2779 (O_2779,N_29815,N_29750);
and UO_2780 (O_2780,N_29816,N_29852);
xor UO_2781 (O_2781,N_29814,N_29953);
xnor UO_2782 (O_2782,N_29749,N_29837);
xnor UO_2783 (O_2783,N_29717,N_29935);
nor UO_2784 (O_2784,N_29811,N_29976);
or UO_2785 (O_2785,N_29974,N_29928);
nor UO_2786 (O_2786,N_29807,N_29708);
nand UO_2787 (O_2787,N_29717,N_29871);
nand UO_2788 (O_2788,N_29858,N_29821);
xnor UO_2789 (O_2789,N_29825,N_29768);
nand UO_2790 (O_2790,N_29829,N_29759);
or UO_2791 (O_2791,N_29723,N_29973);
and UO_2792 (O_2792,N_29869,N_29752);
and UO_2793 (O_2793,N_29874,N_29999);
or UO_2794 (O_2794,N_29929,N_29901);
and UO_2795 (O_2795,N_29994,N_29910);
or UO_2796 (O_2796,N_29814,N_29967);
xnor UO_2797 (O_2797,N_29917,N_29798);
or UO_2798 (O_2798,N_29714,N_29821);
xnor UO_2799 (O_2799,N_29712,N_29799);
and UO_2800 (O_2800,N_29892,N_29975);
nand UO_2801 (O_2801,N_29810,N_29781);
xor UO_2802 (O_2802,N_29932,N_29818);
and UO_2803 (O_2803,N_29921,N_29782);
and UO_2804 (O_2804,N_29727,N_29899);
nand UO_2805 (O_2805,N_29810,N_29777);
xor UO_2806 (O_2806,N_29892,N_29932);
nor UO_2807 (O_2807,N_29916,N_29968);
and UO_2808 (O_2808,N_29828,N_29759);
or UO_2809 (O_2809,N_29769,N_29960);
or UO_2810 (O_2810,N_29744,N_29808);
or UO_2811 (O_2811,N_29936,N_29968);
nand UO_2812 (O_2812,N_29935,N_29926);
nand UO_2813 (O_2813,N_29737,N_29994);
nand UO_2814 (O_2814,N_29919,N_29967);
xnor UO_2815 (O_2815,N_29794,N_29888);
xor UO_2816 (O_2816,N_29998,N_29755);
and UO_2817 (O_2817,N_29843,N_29908);
and UO_2818 (O_2818,N_29921,N_29803);
nand UO_2819 (O_2819,N_29709,N_29974);
and UO_2820 (O_2820,N_29885,N_29924);
xnor UO_2821 (O_2821,N_29871,N_29884);
nor UO_2822 (O_2822,N_29792,N_29891);
and UO_2823 (O_2823,N_29909,N_29836);
or UO_2824 (O_2824,N_29799,N_29783);
nor UO_2825 (O_2825,N_29768,N_29875);
or UO_2826 (O_2826,N_29895,N_29830);
nor UO_2827 (O_2827,N_29934,N_29728);
nand UO_2828 (O_2828,N_29988,N_29760);
or UO_2829 (O_2829,N_29868,N_29830);
or UO_2830 (O_2830,N_29837,N_29819);
or UO_2831 (O_2831,N_29773,N_29717);
and UO_2832 (O_2832,N_29884,N_29989);
nand UO_2833 (O_2833,N_29978,N_29769);
nand UO_2834 (O_2834,N_29891,N_29868);
or UO_2835 (O_2835,N_29839,N_29913);
nor UO_2836 (O_2836,N_29858,N_29848);
nor UO_2837 (O_2837,N_29853,N_29724);
or UO_2838 (O_2838,N_29900,N_29962);
or UO_2839 (O_2839,N_29947,N_29746);
nand UO_2840 (O_2840,N_29839,N_29925);
or UO_2841 (O_2841,N_29744,N_29723);
xnor UO_2842 (O_2842,N_29749,N_29785);
and UO_2843 (O_2843,N_29781,N_29976);
or UO_2844 (O_2844,N_29835,N_29779);
nor UO_2845 (O_2845,N_29914,N_29855);
nand UO_2846 (O_2846,N_29904,N_29736);
xnor UO_2847 (O_2847,N_29962,N_29776);
and UO_2848 (O_2848,N_29732,N_29903);
and UO_2849 (O_2849,N_29860,N_29848);
xnor UO_2850 (O_2850,N_29764,N_29756);
or UO_2851 (O_2851,N_29724,N_29842);
nand UO_2852 (O_2852,N_29943,N_29876);
xnor UO_2853 (O_2853,N_29930,N_29823);
xnor UO_2854 (O_2854,N_29722,N_29783);
xor UO_2855 (O_2855,N_29830,N_29988);
nor UO_2856 (O_2856,N_29840,N_29930);
and UO_2857 (O_2857,N_29927,N_29837);
and UO_2858 (O_2858,N_29787,N_29852);
xor UO_2859 (O_2859,N_29813,N_29922);
nand UO_2860 (O_2860,N_29821,N_29986);
nand UO_2861 (O_2861,N_29778,N_29943);
xnor UO_2862 (O_2862,N_29876,N_29709);
xnor UO_2863 (O_2863,N_29768,N_29882);
xnor UO_2864 (O_2864,N_29772,N_29907);
nor UO_2865 (O_2865,N_29984,N_29773);
nand UO_2866 (O_2866,N_29820,N_29732);
or UO_2867 (O_2867,N_29905,N_29818);
or UO_2868 (O_2868,N_29876,N_29878);
nand UO_2869 (O_2869,N_29935,N_29746);
xor UO_2870 (O_2870,N_29968,N_29921);
and UO_2871 (O_2871,N_29965,N_29974);
xnor UO_2872 (O_2872,N_29755,N_29882);
xor UO_2873 (O_2873,N_29724,N_29705);
and UO_2874 (O_2874,N_29829,N_29944);
nand UO_2875 (O_2875,N_29717,N_29971);
and UO_2876 (O_2876,N_29728,N_29861);
nand UO_2877 (O_2877,N_29733,N_29938);
nand UO_2878 (O_2878,N_29937,N_29935);
or UO_2879 (O_2879,N_29911,N_29757);
nand UO_2880 (O_2880,N_29783,N_29873);
nor UO_2881 (O_2881,N_29951,N_29823);
nor UO_2882 (O_2882,N_29922,N_29867);
nor UO_2883 (O_2883,N_29932,N_29765);
nor UO_2884 (O_2884,N_29889,N_29851);
nor UO_2885 (O_2885,N_29865,N_29821);
nand UO_2886 (O_2886,N_29756,N_29945);
or UO_2887 (O_2887,N_29973,N_29816);
or UO_2888 (O_2888,N_29842,N_29825);
nor UO_2889 (O_2889,N_29720,N_29766);
xnor UO_2890 (O_2890,N_29956,N_29960);
nand UO_2891 (O_2891,N_29821,N_29806);
or UO_2892 (O_2892,N_29987,N_29729);
or UO_2893 (O_2893,N_29737,N_29771);
and UO_2894 (O_2894,N_29964,N_29986);
nand UO_2895 (O_2895,N_29873,N_29952);
nor UO_2896 (O_2896,N_29763,N_29723);
xnor UO_2897 (O_2897,N_29909,N_29785);
and UO_2898 (O_2898,N_29891,N_29955);
nor UO_2899 (O_2899,N_29856,N_29712);
and UO_2900 (O_2900,N_29951,N_29801);
nand UO_2901 (O_2901,N_29757,N_29970);
nand UO_2902 (O_2902,N_29984,N_29862);
nor UO_2903 (O_2903,N_29911,N_29852);
or UO_2904 (O_2904,N_29789,N_29860);
nor UO_2905 (O_2905,N_29986,N_29906);
or UO_2906 (O_2906,N_29823,N_29775);
or UO_2907 (O_2907,N_29802,N_29923);
or UO_2908 (O_2908,N_29756,N_29716);
nand UO_2909 (O_2909,N_29750,N_29820);
and UO_2910 (O_2910,N_29706,N_29970);
or UO_2911 (O_2911,N_29805,N_29757);
xnor UO_2912 (O_2912,N_29968,N_29767);
nand UO_2913 (O_2913,N_29815,N_29846);
nand UO_2914 (O_2914,N_29965,N_29713);
xor UO_2915 (O_2915,N_29799,N_29822);
nor UO_2916 (O_2916,N_29754,N_29867);
nand UO_2917 (O_2917,N_29967,N_29813);
xor UO_2918 (O_2918,N_29920,N_29892);
or UO_2919 (O_2919,N_29971,N_29762);
xnor UO_2920 (O_2920,N_29896,N_29789);
nor UO_2921 (O_2921,N_29922,N_29979);
and UO_2922 (O_2922,N_29767,N_29858);
nand UO_2923 (O_2923,N_29700,N_29924);
xor UO_2924 (O_2924,N_29701,N_29824);
nand UO_2925 (O_2925,N_29979,N_29807);
or UO_2926 (O_2926,N_29967,N_29815);
or UO_2927 (O_2927,N_29831,N_29817);
xnor UO_2928 (O_2928,N_29743,N_29748);
and UO_2929 (O_2929,N_29945,N_29983);
nand UO_2930 (O_2930,N_29824,N_29759);
and UO_2931 (O_2931,N_29798,N_29817);
nand UO_2932 (O_2932,N_29995,N_29919);
or UO_2933 (O_2933,N_29779,N_29889);
and UO_2934 (O_2934,N_29933,N_29967);
and UO_2935 (O_2935,N_29832,N_29814);
xor UO_2936 (O_2936,N_29722,N_29848);
xor UO_2937 (O_2937,N_29962,N_29847);
or UO_2938 (O_2938,N_29967,N_29872);
xnor UO_2939 (O_2939,N_29884,N_29714);
and UO_2940 (O_2940,N_29768,N_29951);
and UO_2941 (O_2941,N_29787,N_29960);
or UO_2942 (O_2942,N_29936,N_29726);
and UO_2943 (O_2943,N_29761,N_29922);
nand UO_2944 (O_2944,N_29709,N_29787);
or UO_2945 (O_2945,N_29827,N_29954);
and UO_2946 (O_2946,N_29804,N_29996);
or UO_2947 (O_2947,N_29921,N_29806);
or UO_2948 (O_2948,N_29925,N_29944);
nand UO_2949 (O_2949,N_29978,N_29727);
xor UO_2950 (O_2950,N_29814,N_29876);
nor UO_2951 (O_2951,N_29813,N_29887);
nand UO_2952 (O_2952,N_29925,N_29942);
and UO_2953 (O_2953,N_29802,N_29787);
and UO_2954 (O_2954,N_29906,N_29761);
or UO_2955 (O_2955,N_29722,N_29977);
or UO_2956 (O_2956,N_29990,N_29810);
xnor UO_2957 (O_2957,N_29942,N_29963);
and UO_2958 (O_2958,N_29934,N_29931);
and UO_2959 (O_2959,N_29800,N_29822);
xor UO_2960 (O_2960,N_29864,N_29986);
nand UO_2961 (O_2961,N_29887,N_29941);
nand UO_2962 (O_2962,N_29918,N_29880);
xnor UO_2963 (O_2963,N_29972,N_29739);
xor UO_2964 (O_2964,N_29938,N_29765);
nand UO_2965 (O_2965,N_29837,N_29976);
or UO_2966 (O_2966,N_29800,N_29777);
nand UO_2967 (O_2967,N_29837,N_29736);
or UO_2968 (O_2968,N_29821,N_29736);
and UO_2969 (O_2969,N_29940,N_29929);
nor UO_2970 (O_2970,N_29945,N_29893);
and UO_2971 (O_2971,N_29940,N_29779);
or UO_2972 (O_2972,N_29815,N_29736);
nand UO_2973 (O_2973,N_29710,N_29850);
and UO_2974 (O_2974,N_29823,N_29750);
xnor UO_2975 (O_2975,N_29967,N_29805);
nand UO_2976 (O_2976,N_29918,N_29865);
xnor UO_2977 (O_2977,N_29885,N_29719);
and UO_2978 (O_2978,N_29928,N_29719);
or UO_2979 (O_2979,N_29924,N_29865);
or UO_2980 (O_2980,N_29904,N_29835);
xor UO_2981 (O_2981,N_29723,N_29831);
nor UO_2982 (O_2982,N_29761,N_29835);
xnor UO_2983 (O_2983,N_29715,N_29783);
nand UO_2984 (O_2984,N_29771,N_29715);
nor UO_2985 (O_2985,N_29942,N_29760);
nand UO_2986 (O_2986,N_29909,N_29888);
nor UO_2987 (O_2987,N_29968,N_29821);
nor UO_2988 (O_2988,N_29892,N_29836);
or UO_2989 (O_2989,N_29892,N_29801);
nor UO_2990 (O_2990,N_29808,N_29786);
xnor UO_2991 (O_2991,N_29907,N_29711);
xnor UO_2992 (O_2992,N_29886,N_29800);
and UO_2993 (O_2993,N_29795,N_29721);
nand UO_2994 (O_2994,N_29732,N_29847);
xor UO_2995 (O_2995,N_29813,N_29976);
nor UO_2996 (O_2996,N_29907,N_29718);
and UO_2997 (O_2997,N_29870,N_29821);
or UO_2998 (O_2998,N_29994,N_29977);
or UO_2999 (O_2999,N_29972,N_29859);
xor UO_3000 (O_3000,N_29932,N_29871);
nand UO_3001 (O_3001,N_29969,N_29981);
or UO_3002 (O_3002,N_29846,N_29869);
and UO_3003 (O_3003,N_29751,N_29771);
xor UO_3004 (O_3004,N_29890,N_29816);
xnor UO_3005 (O_3005,N_29992,N_29737);
nor UO_3006 (O_3006,N_29819,N_29754);
nand UO_3007 (O_3007,N_29903,N_29914);
xor UO_3008 (O_3008,N_29799,N_29815);
nand UO_3009 (O_3009,N_29792,N_29883);
or UO_3010 (O_3010,N_29805,N_29780);
xnor UO_3011 (O_3011,N_29821,N_29789);
nor UO_3012 (O_3012,N_29887,N_29718);
nand UO_3013 (O_3013,N_29978,N_29833);
and UO_3014 (O_3014,N_29736,N_29842);
xnor UO_3015 (O_3015,N_29725,N_29993);
nor UO_3016 (O_3016,N_29834,N_29739);
nor UO_3017 (O_3017,N_29825,N_29767);
or UO_3018 (O_3018,N_29762,N_29943);
nor UO_3019 (O_3019,N_29895,N_29822);
nand UO_3020 (O_3020,N_29766,N_29734);
and UO_3021 (O_3021,N_29774,N_29922);
nor UO_3022 (O_3022,N_29727,N_29703);
or UO_3023 (O_3023,N_29847,N_29772);
xnor UO_3024 (O_3024,N_29742,N_29884);
and UO_3025 (O_3025,N_29925,N_29737);
or UO_3026 (O_3026,N_29931,N_29981);
or UO_3027 (O_3027,N_29916,N_29884);
nor UO_3028 (O_3028,N_29798,N_29984);
nand UO_3029 (O_3029,N_29704,N_29715);
nand UO_3030 (O_3030,N_29785,N_29781);
nand UO_3031 (O_3031,N_29770,N_29711);
xor UO_3032 (O_3032,N_29926,N_29931);
or UO_3033 (O_3033,N_29857,N_29729);
or UO_3034 (O_3034,N_29813,N_29986);
nor UO_3035 (O_3035,N_29927,N_29833);
and UO_3036 (O_3036,N_29903,N_29857);
nand UO_3037 (O_3037,N_29889,N_29756);
or UO_3038 (O_3038,N_29939,N_29752);
xnor UO_3039 (O_3039,N_29974,N_29833);
or UO_3040 (O_3040,N_29996,N_29780);
or UO_3041 (O_3041,N_29932,N_29836);
nand UO_3042 (O_3042,N_29836,N_29997);
or UO_3043 (O_3043,N_29837,N_29908);
or UO_3044 (O_3044,N_29931,N_29954);
and UO_3045 (O_3045,N_29795,N_29941);
xnor UO_3046 (O_3046,N_29739,N_29899);
or UO_3047 (O_3047,N_29984,N_29801);
and UO_3048 (O_3048,N_29718,N_29744);
and UO_3049 (O_3049,N_29877,N_29902);
xor UO_3050 (O_3050,N_29888,N_29848);
or UO_3051 (O_3051,N_29813,N_29731);
or UO_3052 (O_3052,N_29739,N_29747);
xnor UO_3053 (O_3053,N_29702,N_29965);
nor UO_3054 (O_3054,N_29976,N_29719);
nor UO_3055 (O_3055,N_29996,N_29999);
nand UO_3056 (O_3056,N_29755,N_29941);
nor UO_3057 (O_3057,N_29990,N_29834);
or UO_3058 (O_3058,N_29844,N_29922);
and UO_3059 (O_3059,N_29705,N_29706);
xor UO_3060 (O_3060,N_29954,N_29784);
or UO_3061 (O_3061,N_29983,N_29894);
xnor UO_3062 (O_3062,N_29917,N_29851);
or UO_3063 (O_3063,N_29717,N_29913);
nand UO_3064 (O_3064,N_29826,N_29849);
nand UO_3065 (O_3065,N_29856,N_29961);
nand UO_3066 (O_3066,N_29761,N_29831);
and UO_3067 (O_3067,N_29705,N_29899);
nor UO_3068 (O_3068,N_29973,N_29836);
or UO_3069 (O_3069,N_29861,N_29788);
nand UO_3070 (O_3070,N_29960,N_29758);
and UO_3071 (O_3071,N_29828,N_29876);
and UO_3072 (O_3072,N_29911,N_29931);
xor UO_3073 (O_3073,N_29700,N_29758);
nor UO_3074 (O_3074,N_29705,N_29843);
xnor UO_3075 (O_3075,N_29801,N_29794);
xnor UO_3076 (O_3076,N_29941,N_29849);
or UO_3077 (O_3077,N_29877,N_29923);
or UO_3078 (O_3078,N_29778,N_29968);
and UO_3079 (O_3079,N_29811,N_29974);
nand UO_3080 (O_3080,N_29808,N_29880);
nand UO_3081 (O_3081,N_29952,N_29785);
or UO_3082 (O_3082,N_29885,N_29778);
xor UO_3083 (O_3083,N_29930,N_29902);
xnor UO_3084 (O_3084,N_29830,N_29700);
nor UO_3085 (O_3085,N_29879,N_29989);
or UO_3086 (O_3086,N_29982,N_29944);
or UO_3087 (O_3087,N_29941,N_29768);
and UO_3088 (O_3088,N_29868,N_29999);
and UO_3089 (O_3089,N_29983,N_29842);
nand UO_3090 (O_3090,N_29704,N_29840);
and UO_3091 (O_3091,N_29988,N_29989);
xor UO_3092 (O_3092,N_29817,N_29992);
nor UO_3093 (O_3093,N_29888,N_29973);
xor UO_3094 (O_3094,N_29844,N_29875);
nand UO_3095 (O_3095,N_29882,N_29966);
xor UO_3096 (O_3096,N_29858,N_29863);
or UO_3097 (O_3097,N_29771,N_29767);
nand UO_3098 (O_3098,N_29839,N_29797);
xnor UO_3099 (O_3099,N_29951,N_29749);
nor UO_3100 (O_3100,N_29803,N_29748);
and UO_3101 (O_3101,N_29885,N_29739);
nand UO_3102 (O_3102,N_29928,N_29986);
xnor UO_3103 (O_3103,N_29747,N_29917);
or UO_3104 (O_3104,N_29701,N_29707);
nor UO_3105 (O_3105,N_29707,N_29865);
xor UO_3106 (O_3106,N_29814,N_29768);
nand UO_3107 (O_3107,N_29962,N_29729);
or UO_3108 (O_3108,N_29866,N_29808);
nor UO_3109 (O_3109,N_29988,N_29991);
and UO_3110 (O_3110,N_29742,N_29869);
nor UO_3111 (O_3111,N_29952,N_29765);
nor UO_3112 (O_3112,N_29836,N_29702);
nand UO_3113 (O_3113,N_29881,N_29860);
nand UO_3114 (O_3114,N_29822,N_29823);
xor UO_3115 (O_3115,N_29736,N_29721);
xor UO_3116 (O_3116,N_29929,N_29861);
and UO_3117 (O_3117,N_29939,N_29747);
xor UO_3118 (O_3118,N_29805,N_29898);
nand UO_3119 (O_3119,N_29938,N_29738);
or UO_3120 (O_3120,N_29982,N_29865);
or UO_3121 (O_3121,N_29855,N_29847);
xnor UO_3122 (O_3122,N_29942,N_29905);
or UO_3123 (O_3123,N_29839,N_29829);
and UO_3124 (O_3124,N_29737,N_29750);
nor UO_3125 (O_3125,N_29886,N_29748);
nor UO_3126 (O_3126,N_29777,N_29738);
and UO_3127 (O_3127,N_29847,N_29924);
nand UO_3128 (O_3128,N_29705,N_29822);
xor UO_3129 (O_3129,N_29801,N_29753);
nor UO_3130 (O_3130,N_29937,N_29865);
and UO_3131 (O_3131,N_29922,N_29701);
nand UO_3132 (O_3132,N_29860,N_29757);
or UO_3133 (O_3133,N_29810,N_29752);
nand UO_3134 (O_3134,N_29913,N_29882);
and UO_3135 (O_3135,N_29709,N_29861);
xnor UO_3136 (O_3136,N_29992,N_29965);
nand UO_3137 (O_3137,N_29999,N_29828);
nand UO_3138 (O_3138,N_29989,N_29968);
or UO_3139 (O_3139,N_29727,N_29804);
xnor UO_3140 (O_3140,N_29820,N_29834);
or UO_3141 (O_3141,N_29997,N_29784);
nor UO_3142 (O_3142,N_29819,N_29931);
or UO_3143 (O_3143,N_29917,N_29785);
or UO_3144 (O_3144,N_29855,N_29814);
xnor UO_3145 (O_3145,N_29827,N_29801);
nor UO_3146 (O_3146,N_29797,N_29816);
xnor UO_3147 (O_3147,N_29878,N_29993);
or UO_3148 (O_3148,N_29996,N_29986);
and UO_3149 (O_3149,N_29740,N_29861);
and UO_3150 (O_3150,N_29782,N_29862);
nor UO_3151 (O_3151,N_29837,N_29711);
xnor UO_3152 (O_3152,N_29905,N_29951);
nor UO_3153 (O_3153,N_29930,N_29817);
nor UO_3154 (O_3154,N_29754,N_29854);
nor UO_3155 (O_3155,N_29911,N_29863);
nor UO_3156 (O_3156,N_29942,N_29954);
xor UO_3157 (O_3157,N_29844,N_29887);
xnor UO_3158 (O_3158,N_29959,N_29705);
and UO_3159 (O_3159,N_29901,N_29736);
xor UO_3160 (O_3160,N_29763,N_29769);
or UO_3161 (O_3161,N_29888,N_29806);
and UO_3162 (O_3162,N_29936,N_29737);
and UO_3163 (O_3163,N_29758,N_29729);
nor UO_3164 (O_3164,N_29890,N_29876);
and UO_3165 (O_3165,N_29898,N_29770);
and UO_3166 (O_3166,N_29795,N_29700);
or UO_3167 (O_3167,N_29816,N_29972);
xnor UO_3168 (O_3168,N_29875,N_29893);
nor UO_3169 (O_3169,N_29799,N_29985);
nand UO_3170 (O_3170,N_29970,N_29730);
nand UO_3171 (O_3171,N_29845,N_29770);
and UO_3172 (O_3172,N_29901,N_29802);
nor UO_3173 (O_3173,N_29820,N_29833);
xnor UO_3174 (O_3174,N_29863,N_29727);
xnor UO_3175 (O_3175,N_29877,N_29827);
and UO_3176 (O_3176,N_29963,N_29798);
nand UO_3177 (O_3177,N_29818,N_29742);
or UO_3178 (O_3178,N_29945,N_29733);
nand UO_3179 (O_3179,N_29972,N_29706);
nor UO_3180 (O_3180,N_29759,N_29813);
or UO_3181 (O_3181,N_29963,N_29987);
nand UO_3182 (O_3182,N_29707,N_29843);
or UO_3183 (O_3183,N_29788,N_29813);
and UO_3184 (O_3184,N_29859,N_29771);
nand UO_3185 (O_3185,N_29790,N_29854);
nand UO_3186 (O_3186,N_29835,N_29756);
and UO_3187 (O_3187,N_29986,N_29973);
or UO_3188 (O_3188,N_29740,N_29726);
nand UO_3189 (O_3189,N_29796,N_29822);
or UO_3190 (O_3190,N_29734,N_29812);
nor UO_3191 (O_3191,N_29720,N_29761);
or UO_3192 (O_3192,N_29868,N_29758);
and UO_3193 (O_3193,N_29829,N_29857);
nor UO_3194 (O_3194,N_29744,N_29730);
or UO_3195 (O_3195,N_29896,N_29883);
xnor UO_3196 (O_3196,N_29991,N_29849);
or UO_3197 (O_3197,N_29998,N_29840);
nand UO_3198 (O_3198,N_29986,N_29750);
nor UO_3199 (O_3199,N_29861,N_29894);
nor UO_3200 (O_3200,N_29913,N_29939);
nand UO_3201 (O_3201,N_29971,N_29828);
nor UO_3202 (O_3202,N_29987,N_29925);
and UO_3203 (O_3203,N_29806,N_29827);
nand UO_3204 (O_3204,N_29818,N_29768);
nand UO_3205 (O_3205,N_29920,N_29787);
xor UO_3206 (O_3206,N_29970,N_29926);
or UO_3207 (O_3207,N_29965,N_29949);
or UO_3208 (O_3208,N_29922,N_29851);
and UO_3209 (O_3209,N_29971,N_29906);
xnor UO_3210 (O_3210,N_29805,N_29901);
or UO_3211 (O_3211,N_29981,N_29759);
nand UO_3212 (O_3212,N_29942,N_29823);
or UO_3213 (O_3213,N_29703,N_29701);
xor UO_3214 (O_3214,N_29812,N_29769);
nor UO_3215 (O_3215,N_29732,N_29834);
or UO_3216 (O_3216,N_29790,N_29776);
nand UO_3217 (O_3217,N_29786,N_29968);
nand UO_3218 (O_3218,N_29822,N_29825);
and UO_3219 (O_3219,N_29847,N_29895);
nor UO_3220 (O_3220,N_29980,N_29818);
or UO_3221 (O_3221,N_29808,N_29921);
and UO_3222 (O_3222,N_29728,N_29998);
xnor UO_3223 (O_3223,N_29743,N_29988);
or UO_3224 (O_3224,N_29774,N_29847);
nand UO_3225 (O_3225,N_29801,N_29856);
nand UO_3226 (O_3226,N_29815,N_29784);
and UO_3227 (O_3227,N_29874,N_29936);
or UO_3228 (O_3228,N_29946,N_29791);
and UO_3229 (O_3229,N_29897,N_29733);
and UO_3230 (O_3230,N_29872,N_29959);
nor UO_3231 (O_3231,N_29852,N_29702);
nand UO_3232 (O_3232,N_29777,N_29723);
nor UO_3233 (O_3233,N_29899,N_29908);
xor UO_3234 (O_3234,N_29999,N_29800);
nand UO_3235 (O_3235,N_29858,N_29724);
and UO_3236 (O_3236,N_29795,N_29799);
nor UO_3237 (O_3237,N_29858,N_29827);
nand UO_3238 (O_3238,N_29884,N_29917);
nor UO_3239 (O_3239,N_29909,N_29908);
xnor UO_3240 (O_3240,N_29809,N_29821);
nor UO_3241 (O_3241,N_29884,N_29812);
nor UO_3242 (O_3242,N_29905,N_29884);
or UO_3243 (O_3243,N_29805,N_29716);
nor UO_3244 (O_3244,N_29953,N_29911);
and UO_3245 (O_3245,N_29872,N_29748);
or UO_3246 (O_3246,N_29807,N_29893);
nor UO_3247 (O_3247,N_29997,N_29742);
nand UO_3248 (O_3248,N_29892,N_29868);
nand UO_3249 (O_3249,N_29892,N_29911);
and UO_3250 (O_3250,N_29982,N_29726);
nand UO_3251 (O_3251,N_29924,N_29899);
and UO_3252 (O_3252,N_29958,N_29739);
and UO_3253 (O_3253,N_29897,N_29918);
or UO_3254 (O_3254,N_29775,N_29972);
and UO_3255 (O_3255,N_29893,N_29714);
xnor UO_3256 (O_3256,N_29778,N_29960);
nor UO_3257 (O_3257,N_29935,N_29963);
nand UO_3258 (O_3258,N_29791,N_29942);
or UO_3259 (O_3259,N_29881,N_29743);
and UO_3260 (O_3260,N_29898,N_29852);
nand UO_3261 (O_3261,N_29852,N_29859);
or UO_3262 (O_3262,N_29975,N_29781);
or UO_3263 (O_3263,N_29797,N_29997);
xnor UO_3264 (O_3264,N_29709,N_29729);
nor UO_3265 (O_3265,N_29953,N_29725);
nor UO_3266 (O_3266,N_29742,N_29754);
xor UO_3267 (O_3267,N_29748,N_29823);
and UO_3268 (O_3268,N_29746,N_29993);
nand UO_3269 (O_3269,N_29916,N_29994);
and UO_3270 (O_3270,N_29991,N_29746);
and UO_3271 (O_3271,N_29702,N_29775);
xnor UO_3272 (O_3272,N_29734,N_29910);
and UO_3273 (O_3273,N_29932,N_29929);
xor UO_3274 (O_3274,N_29891,N_29775);
xor UO_3275 (O_3275,N_29767,N_29853);
xnor UO_3276 (O_3276,N_29750,N_29864);
nand UO_3277 (O_3277,N_29903,N_29928);
xnor UO_3278 (O_3278,N_29729,N_29907);
xnor UO_3279 (O_3279,N_29811,N_29908);
and UO_3280 (O_3280,N_29719,N_29745);
and UO_3281 (O_3281,N_29846,N_29906);
or UO_3282 (O_3282,N_29832,N_29764);
and UO_3283 (O_3283,N_29958,N_29856);
and UO_3284 (O_3284,N_29919,N_29740);
nand UO_3285 (O_3285,N_29724,N_29995);
or UO_3286 (O_3286,N_29869,N_29898);
or UO_3287 (O_3287,N_29722,N_29836);
nand UO_3288 (O_3288,N_29993,N_29923);
xnor UO_3289 (O_3289,N_29914,N_29772);
or UO_3290 (O_3290,N_29713,N_29860);
xnor UO_3291 (O_3291,N_29910,N_29941);
and UO_3292 (O_3292,N_29910,N_29930);
nand UO_3293 (O_3293,N_29753,N_29976);
xor UO_3294 (O_3294,N_29704,N_29936);
xor UO_3295 (O_3295,N_29841,N_29714);
or UO_3296 (O_3296,N_29840,N_29928);
and UO_3297 (O_3297,N_29812,N_29862);
nor UO_3298 (O_3298,N_29855,N_29795);
xnor UO_3299 (O_3299,N_29722,N_29944);
nor UO_3300 (O_3300,N_29944,N_29713);
xor UO_3301 (O_3301,N_29835,N_29943);
nor UO_3302 (O_3302,N_29846,N_29750);
and UO_3303 (O_3303,N_29855,N_29762);
or UO_3304 (O_3304,N_29836,N_29714);
and UO_3305 (O_3305,N_29709,N_29791);
and UO_3306 (O_3306,N_29968,N_29811);
xnor UO_3307 (O_3307,N_29705,N_29793);
and UO_3308 (O_3308,N_29939,N_29862);
nor UO_3309 (O_3309,N_29953,N_29752);
nor UO_3310 (O_3310,N_29874,N_29716);
xor UO_3311 (O_3311,N_29824,N_29886);
or UO_3312 (O_3312,N_29734,N_29764);
and UO_3313 (O_3313,N_29897,N_29938);
nor UO_3314 (O_3314,N_29787,N_29923);
nor UO_3315 (O_3315,N_29871,N_29723);
nand UO_3316 (O_3316,N_29783,N_29795);
and UO_3317 (O_3317,N_29836,N_29989);
nor UO_3318 (O_3318,N_29850,N_29883);
and UO_3319 (O_3319,N_29830,N_29702);
and UO_3320 (O_3320,N_29823,N_29894);
and UO_3321 (O_3321,N_29824,N_29775);
or UO_3322 (O_3322,N_29889,N_29964);
or UO_3323 (O_3323,N_29892,N_29851);
and UO_3324 (O_3324,N_29771,N_29867);
and UO_3325 (O_3325,N_29997,N_29992);
and UO_3326 (O_3326,N_29988,N_29974);
xnor UO_3327 (O_3327,N_29773,N_29944);
or UO_3328 (O_3328,N_29788,N_29913);
nor UO_3329 (O_3329,N_29929,N_29783);
or UO_3330 (O_3330,N_29803,N_29985);
and UO_3331 (O_3331,N_29785,N_29890);
nor UO_3332 (O_3332,N_29724,N_29928);
or UO_3333 (O_3333,N_29883,N_29966);
xor UO_3334 (O_3334,N_29948,N_29916);
or UO_3335 (O_3335,N_29881,N_29980);
or UO_3336 (O_3336,N_29783,N_29744);
xor UO_3337 (O_3337,N_29978,N_29960);
nand UO_3338 (O_3338,N_29855,N_29937);
nand UO_3339 (O_3339,N_29945,N_29745);
nand UO_3340 (O_3340,N_29928,N_29981);
nand UO_3341 (O_3341,N_29980,N_29773);
nand UO_3342 (O_3342,N_29826,N_29926);
and UO_3343 (O_3343,N_29892,N_29854);
nor UO_3344 (O_3344,N_29865,N_29844);
nand UO_3345 (O_3345,N_29905,N_29844);
and UO_3346 (O_3346,N_29854,N_29702);
xnor UO_3347 (O_3347,N_29893,N_29886);
nand UO_3348 (O_3348,N_29844,N_29771);
xor UO_3349 (O_3349,N_29998,N_29941);
nor UO_3350 (O_3350,N_29814,N_29823);
nand UO_3351 (O_3351,N_29797,N_29895);
or UO_3352 (O_3352,N_29713,N_29871);
or UO_3353 (O_3353,N_29720,N_29882);
nand UO_3354 (O_3354,N_29741,N_29971);
or UO_3355 (O_3355,N_29802,N_29897);
nor UO_3356 (O_3356,N_29725,N_29718);
and UO_3357 (O_3357,N_29920,N_29936);
or UO_3358 (O_3358,N_29984,N_29961);
or UO_3359 (O_3359,N_29965,N_29739);
or UO_3360 (O_3360,N_29761,N_29887);
xnor UO_3361 (O_3361,N_29925,N_29969);
xor UO_3362 (O_3362,N_29893,N_29873);
nor UO_3363 (O_3363,N_29742,N_29795);
and UO_3364 (O_3364,N_29821,N_29706);
xnor UO_3365 (O_3365,N_29904,N_29911);
nor UO_3366 (O_3366,N_29982,N_29925);
and UO_3367 (O_3367,N_29956,N_29834);
xnor UO_3368 (O_3368,N_29768,N_29796);
nand UO_3369 (O_3369,N_29824,N_29991);
and UO_3370 (O_3370,N_29828,N_29765);
nand UO_3371 (O_3371,N_29920,N_29923);
nand UO_3372 (O_3372,N_29897,N_29765);
nor UO_3373 (O_3373,N_29725,N_29977);
nand UO_3374 (O_3374,N_29729,N_29790);
nor UO_3375 (O_3375,N_29843,N_29902);
or UO_3376 (O_3376,N_29802,N_29872);
and UO_3377 (O_3377,N_29732,N_29933);
or UO_3378 (O_3378,N_29841,N_29902);
or UO_3379 (O_3379,N_29816,N_29928);
or UO_3380 (O_3380,N_29901,N_29706);
or UO_3381 (O_3381,N_29718,N_29874);
nor UO_3382 (O_3382,N_29922,N_29827);
nor UO_3383 (O_3383,N_29795,N_29970);
and UO_3384 (O_3384,N_29770,N_29827);
or UO_3385 (O_3385,N_29930,N_29751);
nand UO_3386 (O_3386,N_29882,N_29826);
xor UO_3387 (O_3387,N_29702,N_29875);
xnor UO_3388 (O_3388,N_29791,N_29914);
xnor UO_3389 (O_3389,N_29825,N_29980);
nand UO_3390 (O_3390,N_29892,N_29834);
and UO_3391 (O_3391,N_29946,N_29867);
nor UO_3392 (O_3392,N_29793,N_29721);
and UO_3393 (O_3393,N_29890,N_29866);
or UO_3394 (O_3394,N_29842,N_29890);
nor UO_3395 (O_3395,N_29760,N_29881);
nand UO_3396 (O_3396,N_29719,N_29825);
xnor UO_3397 (O_3397,N_29930,N_29730);
or UO_3398 (O_3398,N_29744,N_29976);
and UO_3399 (O_3399,N_29975,N_29711);
nor UO_3400 (O_3400,N_29725,N_29807);
xnor UO_3401 (O_3401,N_29813,N_29783);
nand UO_3402 (O_3402,N_29754,N_29833);
or UO_3403 (O_3403,N_29852,N_29846);
nor UO_3404 (O_3404,N_29827,N_29854);
xor UO_3405 (O_3405,N_29701,N_29706);
nor UO_3406 (O_3406,N_29980,N_29863);
or UO_3407 (O_3407,N_29748,N_29810);
or UO_3408 (O_3408,N_29963,N_29777);
and UO_3409 (O_3409,N_29747,N_29738);
nand UO_3410 (O_3410,N_29764,N_29879);
nand UO_3411 (O_3411,N_29946,N_29729);
xnor UO_3412 (O_3412,N_29809,N_29964);
and UO_3413 (O_3413,N_29967,N_29948);
xnor UO_3414 (O_3414,N_29913,N_29793);
nor UO_3415 (O_3415,N_29742,N_29763);
nand UO_3416 (O_3416,N_29974,N_29930);
or UO_3417 (O_3417,N_29971,N_29876);
and UO_3418 (O_3418,N_29816,N_29986);
nand UO_3419 (O_3419,N_29981,N_29924);
or UO_3420 (O_3420,N_29993,N_29794);
nor UO_3421 (O_3421,N_29920,N_29971);
nand UO_3422 (O_3422,N_29994,N_29864);
xnor UO_3423 (O_3423,N_29977,N_29885);
xnor UO_3424 (O_3424,N_29863,N_29943);
xnor UO_3425 (O_3425,N_29993,N_29827);
xnor UO_3426 (O_3426,N_29742,N_29854);
nand UO_3427 (O_3427,N_29860,N_29970);
xnor UO_3428 (O_3428,N_29734,N_29846);
or UO_3429 (O_3429,N_29822,N_29923);
nand UO_3430 (O_3430,N_29861,N_29838);
xnor UO_3431 (O_3431,N_29964,N_29990);
nand UO_3432 (O_3432,N_29899,N_29883);
nand UO_3433 (O_3433,N_29752,N_29794);
nor UO_3434 (O_3434,N_29883,N_29926);
nand UO_3435 (O_3435,N_29819,N_29857);
nand UO_3436 (O_3436,N_29937,N_29778);
xnor UO_3437 (O_3437,N_29834,N_29825);
and UO_3438 (O_3438,N_29986,N_29823);
xnor UO_3439 (O_3439,N_29813,N_29989);
xor UO_3440 (O_3440,N_29720,N_29939);
or UO_3441 (O_3441,N_29810,N_29872);
xnor UO_3442 (O_3442,N_29993,N_29721);
xnor UO_3443 (O_3443,N_29715,N_29808);
nand UO_3444 (O_3444,N_29850,N_29815);
and UO_3445 (O_3445,N_29881,N_29775);
or UO_3446 (O_3446,N_29812,N_29793);
nand UO_3447 (O_3447,N_29961,N_29735);
xor UO_3448 (O_3448,N_29849,N_29831);
or UO_3449 (O_3449,N_29787,N_29765);
and UO_3450 (O_3450,N_29982,N_29857);
and UO_3451 (O_3451,N_29811,N_29929);
nor UO_3452 (O_3452,N_29953,N_29832);
nor UO_3453 (O_3453,N_29784,N_29723);
and UO_3454 (O_3454,N_29767,N_29963);
xnor UO_3455 (O_3455,N_29834,N_29873);
and UO_3456 (O_3456,N_29949,N_29814);
or UO_3457 (O_3457,N_29714,N_29737);
and UO_3458 (O_3458,N_29849,N_29841);
xnor UO_3459 (O_3459,N_29874,N_29722);
and UO_3460 (O_3460,N_29976,N_29856);
nor UO_3461 (O_3461,N_29742,N_29756);
nand UO_3462 (O_3462,N_29900,N_29708);
and UO_3463 (O_3463,N_29764,N_29884);
nand UO_3464 (O_3464,N_29811,N_29861);
nor UO_3465 (O_3465,N_29967,N_29787);
or UO_3466 (O_3466,N_29944,N_29943);
nand UO_3467 (O_3467,N_29933,N_29975);
nand UO_3468 (O_3468,N_29706,N_29707);
and UO_3469 (O_3469,N_29800,N_29941);
and UO_3470 (O_3470,N_29758,N_29794);
and UO_3471 (O_3471,N_29912,N_29780);
nand UO_3472 (O_3472,N_29890,N_29961);
or UO_3473 (O_3473,N_29952,N_29882);
or UO_3474 (O_3474,N_29896,N_29755);
or UO_3475 (O_3475,N_29798,N_29729);
nor UO_3476 (O_3476,N_29827,N_29901);
nor UO_3477 (O_3477,N_29721,N_29895);
or UO_3478 (O_3478,N_29944,N_29962);
xor UO_3479 (O_3479,N_29930,N_29735);
and UO_3480 (O_3480,N_29725,N_29787);
or UO_3481 (O_3481,N_29767,N_29758);
or UO_3482 (O_3482,N_29899,N_29733);
or UO_3483 (O_3483,N_29927,N_29760);
or UO_3484 (O_3484,N_29792,N_29717);
or UO_3485 (O_3485,N_29704,N_29939);
nor UO_3486 (O_3486,N_29824,N_29704);
or UO_3487 (O_3487,N_29779,N_29799);
and UO_3488 (O_3488,N_29818,N_29920);
or UO_3489 (O_3489,N_29729,N_29708);
nor UO_3490 (O_3490,N_29842,N_29953);
nor UO_3491 (O_3491,N_29835,N_29993);
xor UO_3492 (O_3492,N_29853,N_29967);
and UO_3493 (O_3493,N_29889,N_29741);
nand UO_3494 (O_3494,N_29889,N_29736);
xor UO_3495 (O_3495,N_29747,N_29710);
or UO_3496 (O_3496,N_29910,N_29832);
or UO_3497 (O_3497,N_29916,N_29944);
and UO_3498 (O_3498,N_29842,N_29831);
and UO_3499 (O_3499,N_29851,N_29925);
endmodule