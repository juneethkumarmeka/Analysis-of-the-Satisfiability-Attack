module basic_500_3000_500_6_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_462,In_242);
nor U1 (N_1,In_87,In_216);
nor U2 (N_2,In_178,In_266);
or U3 (N_3,In_147,In_268);
nor U4 (N_4,In_234,In_196);
xor U5 (N_5,In_374,In_494);
xor U6 (N_6,In_267,In_69);
nor U7 (N_7,In_390,In_326);
or U8 (N_8,In_394,In_411);
and U9 (N_9,In_354,In_324);
nor U10 (N_10,In_56,In_412);
and U11 (N_11,In_372,In_250);
or U12 (N_12,In_71,In_150);
or U13 (N_13,In_437,In_161);
and U14 (N_14,In_153,In_193);
nand U15 (N_15,In_103,In_88);
and U16 (N_16,In_190,In_291);
or U17 (N_17,In_49,In_122);
nand U18 (N_18,In_377,In_227);
or U19 (N_19,In_458,In_471);
nor U20 (N_20,In_422,In_481);
nand U21 (N_21,In_15,In_156);
xor U22 (N_22,In_138,In_479);
and U23 (N_23,In_383,In_259);
nand U24 (N_24,In_188,In_381);
and U25 (N_25,In_451,In_102);
xor U26 (N_26,In_167,In_106);
or U27 (N_27,In_172,In_319);
and U28 (N_28,In_455,In_357);
nor U29 (N_29,In_292,In_101);
nor U30 (N_30,In_174,In_154);
and U31 (N_31,In_456,In_264);
xnor U32 (N_32,In_429,In_197);
and U33 (N_33,In_212,In_339);
nand U34 (N_34,In_139,In_7);
or U35 (N_35,In_306,In_191);
xor U36 (N_36,In_130,In_123);
nand U37 (N_37,In_163,In_401);
and U38 (N_38,In_366,In_447);
nand U39 (N_39,In_485,In_72);
nand U40 (N_40,In_157,In_359);
nand U41 (N_41,In_367,In_175);
nor U42 (N_42,In_270,In_426);
or U43 (N_43,In_119,In_93);
nand U44 (N_44,In_322,In_10);
nand U45 (N_45,In_441,In_311);
and U46 (N_46,In_287,In_499);
and U47 (N_47,In_125,In_109);
nand U48 (N_48,In_21,In_98);
nor U49 (N_49,In_491,In_81);
nand U50 (N_50,In_201,In_151);
nor U51 (N_51,In_168,In_379);
nand U52 (N_52,In_364,In_164);
xnor U53 (N_53,In_137,In_331);
and U54 (N_54,In_111,In_64);
and U55 (N_55,In_496,In_179);
nand U56 (N_56,In_425,In_276);
nor U57 (N_57,In_31,In_129);
xor U58 (N_58,In_313,In_246);
nand U59 (N_59,In_240,In_484);
or U60 (N_60,In_296,In_382);
nor U61 (N_61,In_121,In_158);
or U62 (N_62,In_89,In_112);
or U63 (N_63,In_440,In_208);
and U64 (N_64,In_396,In_423);
nor U65 (N_65,In_171,In_32);
nand U66 (N_66,In_399,In_117);
xor U67 (N_67,In_0,In_41);
nand U68 (N_68,In_74,In_173);
nand U69 (N_69,In_134,In_397);
or U70 (N_70,In_323,In_464);
nand U71 (N_71,In_419,In_6);
or U72 (N_72,In_460,In_42);
nor U73 (N_73,In_220,In_206);
or U74 (N_74,In_439,In_207);
xor U75 (N_75,In_497,In_343);
or U76 (N_76,In_127,In_20);
nand U77 (N_77,In_90,In_335);
xor U78 (N_78,In_378,In_337);
and U79 (N_79,In_189,In_180);
xor U80 (N_80,In_493,In_318);
nand U81 (N_81,In_124,In_184);
nor U82 (N_82,In_146,In_169);
nand U83 (N_83,In_310,In_211);
nand U84 (N_84,In_376,In_434);
xnor U85 (N_85,In_239,In_24);
xor U86 (N_86,In_299,In_488);
xnor U87 (N_87,In_149,In_27);
or U88 (N_88,In_97,In_58);
nand U89 (N_89,In_294,In_274);
nor U90 (N_90,In_332,In_309);
or U91 (N_91,In_312,In_25);
xnor U92 (N_92,In_1,In_414);
xor U93 (N_93,In_51,In_62);
xnor U94 (N_94,In_77,In_83);
xor U95 (N_95,In_386,In_482);
and U96 (N_96,In_302,In_36);
and U97 (N_97,In_215,In_473);
nand U98 (N_98,In_255,In_445);
nand U99 (N_99,In_293,In_105);
or U100 (N_100,In_281,In_436);
or U101 (N_101,In_14,In_258);
nand U102 (N_102,In_286,In_280);
or U103 (N_103,In_263,In_476);
nor U104 (N_104,In_143,In_65);
and U105 (N_105,In_80,In_224);
and U106 (N_106,In_34,In_5);
and U107 (N_107,In_356,In_465);
or U108 (N_108,In_282,In_265);
xnor U109 (N_109,In_131,In_141);
nand U110 (N_110,In_373,In_30);
or U111 (N_111,In_39,In_432);
or U112 (N_112,In_495,In_384);
nor U113 (N_113,In_126,In_79);
and U114 (N_114,In_444,In_204);
or U115 (N_115,In_85,In_348);
nand U116 (N_116,In_375,In_229);
nand U117 (N_117,In_107,In_413);
nor U118 (N_118,In_132,In_448);
or U119 (N_119,In_285,In_162);
nand U120 (N_120,In_8,In_483);
nor U121 (N_121,In_75,In_334);
and U122 (N_122,In_490,In_78);
xnor U123 (N_123,In_408,In_283);
and U124 (N_124,In_279,In_290);
or U125 (N_125,In_463,In_450);
nor U126 (N_126,In_477,In_320);
nor U127 (N_127,In_289,In_330);
nand U128 (N_128,In_452,In_144);
and U129 (N_129,In_55,In_371);
xnor U130 (N_130,In_235,In_478);
xor U131 (N_131,In_469,In_388);
and U132 (N_132,In_489,In_213);
nor U133 (N_133,In_275,In_245);
xnor U134 (N_134,In_316,In_177);
xnor U135 (N_135,In_389,In_185);
xor U136 (N_136,In_438,In_116);
nor U137 (N_137,In_244,In_152);
and U138 (N_138,In_38,In_203);
xor U139 (N_139,In_353,In_314);
xnor U140 (N_140,In_182,In_108);
nand U141 (N_141,In_237,In_403);
nand U142 (N_142,In_99,In_352);
nor U143 (N_143,In_317,In_176);
or U144 (N_144,In_349,In_346);
xnor U145 (N_145,In_159,In_219);
and U146 (N_146,In_387,In_492);
and U147 (N_147,In_233,In_420);
or U148 (N_148,In_136,In_18);
and U149 (N_149,In_22,In_252);
or U150 (N_150,In_192,In_53);
and U151 (N_151,In_43,In_298);
or U152 (N_152,In_160,In_84);
and U153 (N_153,In_115,In_46);
nor U154 (N_154,In_170,In_454);
or U155 (N_155,In_57,In_37);
xnor U156 (N_156,In_230,In_363);
or U157 (N_157,In_241,In_23);
and U158 (N_158,In_68,In_35);
xnor U159 (N_159,In_305,In_205);
xnor U160 (N_160,In_166,In_328);
nand U161 (N_161,In_406,In_256);
and U162 (N_162,In_315,In_52);
nand U163 (N_163,In_91,In_214);
nor U164 (N_164,In_453,In_249);
nor U165 (N_165,In_13,In_321);
or U166 (N_166,In_409,In_195);
nand U167 (N_167,In_307,In_110);
xor U168 (N_168,In_466,In_95);
xor U169 (N_169,In_198,In_398);
and U170 (N_170,In_61,In_247);
nor U171 (N_171,In_135,In_449);
nor U172 (N_172,In_325,In_474);
or U173 (N_173,In_186,In_243);
or U174 (N_174,In_407,In_44);
xor U175 (N_175,In_418,In_142);
and U176 (N_176,In_100,In_16);
xnor U177 (N_177,In_350,In_114);
and U178 (N_178,In_4,In_427);
nand U179 (N_179,In_118,In_128);
and U180 (N_180,In_33,In_475);
xor U181 (N_181,In_200,In_48);
nand U182 (N_182,In_155,In_442);
or U183 (N_183,In_26,In_248);
xor U184 (N_184,In_40,In_217);
or U185 (N_185,In_301,In_54);
or U186 (N_186,In_12,In_113);
or U187 (N_187,In_210,In_470);
xor U188 (N_188,In_165,In_28);
xor U189 (N_189,In_254,In_410);
xnor U190 (N_190,In_29,In_368);
and U191 (N_191,In_86,In_459);
nand U192 (N_192,In_392,In_120);
xnor U193 (N_193,In_341,In_278);
nand U194 (N_194,In_370,In_424);
nand U195 (N_195,In_443,In_104);
and U196 (N_196,In_202,In_288);
nand U197 (N_197,In_96,In_238);
and U198 (N_198,In_277,In_486);
or U199 (N_199,In_9,In_405);
nand U200 (N_200,In_336,In_416);
xnor U201 (N_201,In_63,In_187);
nor U202 (N_202,In_428,In_480);
nor U203 (N_203,In_404,In_262);
and U204 (N_204,In_194,In_218);
and U205 (N_205,In_461,In_272);
nor U206 (N_206,In_430,In_271);
xnor U207 (N_207,In_385,In_226);
nor U208 (N_208,In_360,In_236);
or U209 (N_209,In_199,In_140);
xnor U210 (N_210,In_342,In_221);
or U211 (N_211,In_347,In_2);
xnor U212 (N_212,In_231,In_365);
nand U213 (N_213,In_433,In_468);
and U214 (N_214,In_369,In_82);
and U215 (N_215,In_225,In_183);
or U216 (N_216,In_329,In_209);
nor U217 (N_217,In_92,In_344);
and U218 (N_218,In_415,In_73);
nor U219 (N_219,In_50,In_395);
and U220 (N_220,In_59,In_284);
xnor U221 (N_221,In_261,In_421);
and U222 (N_222,In_380,In_60);
xnor U223 (N_223,In_223,In_17);
nor U224 (N_224,In_472,In_70);
nand U225 (N_225,In_327,In_145);
or U226 (N_226,In_232,In_457);
or U227 (N_227,In_11,In_393);
xnor U228 (N_228,In_47,In_345);
and U229 (N_229,In_351,In_487);
or U230 (N_230,In_45,In_308);
xnor U231 (N_231,In_417,In_400);
nor U232 (N_232,In_431,In_133);
or U233 (N_233,In_222,In_297);
or U234 (N_234,In_251,In_257);
nand U235 (N_235,In_253,In_19);
xor U236 (N_236,In_338,In_402);
nand U237 (N_237,In_361,In_148);
and U238 (N_238,In_66,In_467);
nor U239 (N_239,In_273,In_181);
nand U240 (N_240,In_498,In_304);
nor U241 (N_241,In_446,In_303);
or U242 (N_242,In_228,In_300);
and U243 (N_243,In_355,In_362);
and U244 (N_244,In_295,In_67);
or U245 (N_245,In_391,In_340);
nor U246 (N_246,In_358,In_94);
and U247 (N_247,In_3,In_260);
nand U248 (N_248,In_333,In_435);
xor U249 (N_249,In_269,In_76);
nor U250 (N_250,In_462,In_54);
nor U251 (N_251,In_424,In_233);
or U252 (N_252,In_411,In_383);
nand U253 (N_253,In_242,In_299);
xnor U254 (N_254,In_52,In_403);
or U255 (N_255,In_319,In_264);
nor U256 (N_256,In_445,In_383);
xor U257 (N_257,In_83,In_484);
xnor U258 (N_258,In_365,In_404);
nor U259 (N_259,In_299,In_121);
nor U260 (N_260,In_345,In_152);
nor U261 (N_261,In_299,In_108);
and U262 (N_262,In_451,In_307);
and U263 (N_263,In_407,In_150);
nor U264 (N_264,In_213,In_295);
and U265 (N_265,In_342,In_278);
nor U266 (N_266,In_494,In_146);
xnor U267 (N_267,In_259,In_484);
xor U268 (N_268,In_345,In_431);
and U269 (N_269,In_323,In_200);
nand U270 (N_270,In_430,In_2);
xor U271 (N_271,In_218,In_340);
nand U272 (N_272,In_404,In_340);
and U273 (N_273,In_294,In_394);
and U274 (N_274,In_306,In_246);
nor U275 (N_275,In_493,In_411);
or U276 (N_276,In_324,In_264);
xor U277 (N_277,In_126,In_393);
xor U278 (N_278,In_182,In_373);
nor U279 (N_279,In_40,In_393);
or U280 (N_280,In_75,In_247);
xor U281 (N_281,In_248,In_244);
nand U282 (N_282,In_292,In_180);
and U283 (N_283,In_90,In_349);
nor U284 (N_284,In_13,In_357);
xnor U285 (N_285,In_45,In_35);
nand U286 (N_286,In_41,In_274);
xor U287 (N_287,In_459,In_238);
nand U288 (N_288,In_66,In_7);
xor U289 (N_289,In_439,In_383);
xor U290 (N_290,In_171,In_206);
nor U291 (N_291,In_406,In_496);
and U292 (N_292,In_152,In_293);
xnor U293 (N_293,In_119,In_229);
or U294 (N_294,In_49,In_342);
xor U295 (N_295,In_351,In_5);
nor U296 (N_296,In_466,In_18);
nor U297 (N_297,In_132,In_302);
nand U298 (N_298,In_355,In_250);
nor U299 (N_299,In_274,In_273);
xnor U300 (N_300,In_223,In_177);
or U301 (N_301,In_447,In_260);
and U302 (N_302,In_495,In_361);
nor U303 (N_303,In_255,In_201);
nor U304 (N_304,In_64,In_446);
nand U305 (N_305,In_442,In_283);
or U306 (N_306,In_317,In_360);
xnor U307 (N_307,In_453,In_189);
or U308 (N_308,In_192,In_193);
or U309 (N_309,In_126,In_136);
xor U310 (N_310,In_90,In_144);
nor U311 (N_311,In_393,In_438);
nand U312 (N_312,In_412,In_260);
and U313 (N_313,In_441,In_91);
or U314 (N_314,In_280,In_144);
or U315 (N_315,In_405,In_27);
nand U316 (N_316,In_222,In_7);
nor U317 (N_317,In_488,In_420);
or U318 (N_318,In_341,In_422);
nor U319 (N_319,In_99,In_283);
or U320 (N_320,In_130,In_120);
xor U321 (N_321,In_477,In_198);
nor U322 (N_322,In_178,In_146);
or U323 (N_323,In_113,In_171);
and U324 (N_324,In_66,In_135);
xor U325 (N_325,In_93,In_101);
xnor U326 (N_326,In_262,In_276);
or U327 (N_327,In_432,In_255);
or U328 (N_328,In_124,In_349);
nand U329 (N_329,In_66,In_88);
and U330 (N_330,In_41,In_284);
nand U331 (N_331,In_66,In_108);
nand U332 (N_332,In_126,In_4);
or U333 (N_333,In_111,In_328);
nor U334 (N_334,In_212,In_278);
nor U335 (N_335,In_395,In_182);
nor U336 (N_336,In_466,In_277);
or U337 (N_337,In_297,In_431);
nor U338 (N_338,In_140,In_88);
and U339 (N_339,In_218,In_498);
or U340 (N_340,In_17,In_423);
nand U341 (N_341,In_150,In_277);
nor U342 (N_342,In_334,In_109);
nor U343 (N_343,In_36,In_382);
nor U344 (N_344,In_8,In_341);
or U345 (N_345,In_343,In_323);
nand U346 (N_346,In_177,In_12);
or U347 (N_347,In_221,In_109);
nor U348 (N_348,In_197,In_472);
nor U349 (N_349,In_149,In_48);
nand U350 (N_350,In_349,In_323);
xor U351 (N_351,In_448,In_499);
or U352 (N_352,In_188,In_228);
nor U353 (N_353,In_140,In_139);
nand U354 (N_354,In_297,In_225);
nand U355 (N_355,In_300,In_99);
or U356 (N_356,In_297,In_44);
xor U357 (N_357,In_414,In_15);
and U358 (N_358,In_200,In_106);
nand U359 (N_359,In_201,In_138);
and U360 (N_360,In_240,In_245);
or U361 (N_361,In_212,In_14);
nand U362 (N_362,In_191,In_314);
xnor U363 (N_363,In_452,In_261);
nor U364 (N_364,In_108,In_499);
nor U365 (N_365,In_355,In_24);
nand U366 (N_366,In_256,In_436);
or U367 (N_367,In_72,In_235);
xnor U368 (N_368,In_232,In_163);
or U369 (N_369,In_24,In_233);
xor U370 (N_370,In_266,In_244);
or U371 (N_371,In_379,In_182);
nand U372 (N_372,In_132,In_304);
nor U373 (N_373,In_260,In_113);
nand U374 (N_374,In_89,In_256);
nor U375 (N_375,In_316,In_0);
or U376 (N_376,In_282,In_351);
nand U377 (N_377,In_325,In_278);
and U378 (N_378,In_441,In_106);
or U379 (N_379,In_95,In_491);
nor U380 (N_380,In_235,In_52);
and U381 (N_381,In_265,In_151);
xor U382 (N_382,In_486,In_419);
and U383 (N_383,In_447,In_83);
and U384 (N_384,In_142,In_436);
nor U385 (N_385,In_110,In_14);
and U386 (N_386,In_65,In_218);
or U387 (N_387,In_302,In_408);
nor U388 (N_388,In_189,In_213);
and U389 (N_389,In_179,In_112);
nor U390 (N_390,In_224,In_373);
nor U391 (N_391,In_332,In_415);
nor U392 (N_392,In_265,In_115);
and U393 (N_393,In_343,In_187);
xor U394 (N_394,In_392,In_138);
xor U395 (N_395,In_213,In_60);
and U396 (N_396,In_407,In_212);
and U397 (N_397,In_192,In_381);
or U398 (N_398,In_125,In_128);
xnor U399 (N_399,In_346,In_417);
and U400 (N_400,In_72,In_143);
nand U401 (N_401,In_306,In_403);
nand U402 (N_402,In_400,In_277);
xnor U403 (N_403,In_232,In_330);
nand U404 (N_404,In_273,In_39);
or U405 (N_405,In_112,In_37);
or U406 (N_406,In_400,In_249);
or U407 (N_407,In_75,In_255);
nor U408 (N_408,In_472,In_19);
xor U409 (N_409,In_103,In_424);
or U410 (N_410,In_106,In_60);
nand U411 (N_411,In_96,In_218);
and U412 (N_412,In_65,In_231);
nor U413 (N_413,In_75,In_204);
and U414 (N_414,In_283,In_320);
and U415 (N_415,In_45,In_366);
nor U416 (N_416,In_396,In_103);
and U417 (N_417,In_66,In_210);
or U418 (N_418,In_104,In_457);
or U419 (N_419,In_477,In_46);
xnor U420 (N_420,In_404,In_9);
xor U421 (N_421,In_62,In_319);
xnor U422 (N_422,In_90,In_318);
nor U423 (N_423,In_343,In_136);
and U424 (N_424,In_46,In_1);
and U425 (N_425,In_256,In_329);
nand U426 (N_426,In_299,In_124);
or U427 (N_427,In_266,In_241);
and U428 (N_428,In_259,In_426);
and U429 (N_429,In_35,In_266);
xor U430 (N_430,In_265,In_66);
nor U431 (N_431,In_306,In_313);
nand U432 (N_432,In_468,In_318);
nor U433 (N_433,In_477,In_89);
xor U434 (N_434,In_156,In_98);
nor U435 (N_435,In_370,In_224);
and U436 (N_436,In_131,In_203);
nor U437 (N_437,In_236,In_490);
and U438 (N_438,In_91,In_310);
and U439 (N_439,In_351,In_456);
or U440 (N_440,In_100,In_352);
xor U441 (N_441,In_74,In_351);
or U442 (N_442,In_317,In_129);
nand U443 (N_443,In_122,In_143);
or U444 (N_444,In_159,In_372);
or U445 (N_445,In_267,In_143);
or U446 (N_446,In_410,In_173);
or U447 (N_447,In_110,In_130);
nand U448 (N_448,In_362,In_470);
nand U449 (N_449,In_402,In_81);
or U450 (N_450,In_81,In_263);
or U451 (N_451,In_266,In_58);
nor U452 (N_452,In_393,In_76);
nor U453 (N_453,In_248,In_342);
and U454 (N_454,In_391,In_425);
and U455 (N_455,In_94,In_467);
xor U456 (N_456,In_386,In_200);
and U457 (N_457,In_61,In_326);
and U458 (N_458,In_95,In_472);
xnor U459 (N_459,In_326,In_386);
nor U460 (N_460,In_357,In_167);
xor U461 (N_461,In_16,In_464);
and U462 (N_462,In_440,In_104);
or U463 (N_463,In_122,In_428);
and U464 (N_464,In_400,In_337);
or U465 (N_465,In_80,In_296);
or U466 (N_466,In_184,In_22);
nor U467 (N_467,In_68,In_345);
nor U468 (N_468,In_24,In_255);
nand U469 (N_469,In_484,In_302);
nand U470 (N_470,In_244,In_211);
or U471 (N_471,In_480,In_230);
or U472 (N_472,In_494,In_410);
xnor U473 (N_473,In_121,In_311);
and U474 (N_474,In_483,In_82);
or U475 (N_475,In_193,In_207);
or U476 (N_476,In_307,In_341);
xor U477 (N_477,In_59,In_445);
xor U478 (N_478,In_287,In_442);
xnor U479 (N_479,In_154,In_369);
nor U480 (N_480,In_344,In_211);
xor U481 (N_481,In_468,In_483);
or U482 (N_482,In_398,In_20);
or U483 (N_483,In_199,In_151);
or U484 (N_484,In_187,In_100);
xnor U485 (N_485,In_362,In_60);
nand U486 (N_486,In_162,In_400);
nor U487 (N_487,In_226,In_242);
and U488 (N_488,In_114,In_444);
or U489 (N_489,In_119,In_194);
and U490 (N_490,In_383,In_117);
or U491 (N_491,In_119,In_12);
or U492 (N_492,In_40,In_321);
or U493 (N_493,In_362,In_73);
or U494 (N_494,In_268,In_255);
xnor U495 (N_495,In_368,In_166);
xnor U496 (N_496,In_488,In_314);
nor U497 (N_497,In_6,In_224);
nor U498 (N_498,In_83,In_493);
nor U499 (N_499,In_474,In_348);
xor U500 (N_500,N_401,N_44);
nor U501 (N_501,N_300,N_232);
or U502 (N_502,N_445,N_324);
and U503 (N_503,N_180,N_349);
and U504 (N_504,N_385,N_475);
or U505 (N_505,N_163,N_468);
nand U506 (N_506,N_463,N_425);
and U507 (N_507,N_260,N_117);
nand U508 (N_508,N_166,N_162);
and U509 (N_509,N_296,N_101);
nor U510 (N_510,N_388,N_494);
and U511 (N_511,N_198,N_49);
and U512 (N_512,N_103,N_375);
or U513 (N_513,N_179,N_244);
nand U514 (N_514,N_4,N_146);
nor U515 (N_515,N_271,N_341);
xor U516 (N_516,N_334,N_18);
nand U517 (N_517,N_110,N_36);
nor U518 (N_518,N_245,N_471);
xnor U519 (N_519,N_48,N_92);
nand U520 (N_520,N_160,N_132);
nand U521 (N_521,N_256,N_342);
nor U522 (N_522,N_59,N_178);
nand U523 (N_523,N_99,N_81);
nand U524 (N_524,N_236,N_255);
nand U525 (N_525,N_0,N_104);
xor U526 (N_526,N_403,N_25);
nand U527 (N_527,N_220,N_69);
nor U528 (N_528,N_108,N_135);
and U529 (N_529,N_203,N_136);
and U530 (N_530,N_215,N_249);
or U531 (N_531,N_268,N_386);
and U532 (N_532,N_477,N_306);
and U533 (N_533,N_344,N_408);
or U534 (N_534,N_455,N_481);
xnor U535 (N_535,N_235,N_343);
xor U536 (N_536,N_60,N_152);
or U537 (N_537,N_347,N_176);
nor U538 (N_538,N_2,N_482);
and U539 (N_539,N_71,N_302);
or U540 (N_540,N_439,N_157);
nand U541 (N_541,N_274,N_363);
xnor U542 (N_542,N_116,N_214);
nand U543 (N_543,N_238,N_270);
and U544 (N_544,N_358,N_243);
xnor U545 (N_545,N_242,N_47);
xor U546 (N_546,N_45,N_451);
and U547 (N_547,N_326,N_170);
nor U548 (N_548,N_400,N_219);
and U549 (N_549,N_57,N_464);
xnor U550 (N_550,N_356,N_141);
and U551 (N_551,N_66,N_395);
and U552 (N_552,N_191,N_453);
nor U553 (N_553,N_221,N_419);
xor U554 (N_554,N_457,N_377);
nor U555 (N_555,N_320,N_113);
and U556 (N_556,N_458,N_133);
nand U557 (N_557,N_337,N_95);
xor U558 (N_558,N_246,N_360);
or U559 (N_559,N_391,N_74);
and U560 (N_560,N_366,N_493);
and U561 (N_561,N_79,N_291);
and U562 (N_562,N_316,N_308);
or U563 (N_563,N_143,N_28);
nand U564 (N_564,N_369,N_240);
nor U565 (N_565,N_350,N_126);
and U566 (N_566,N_259,N_367);
nor U567 (N_567,N_177,N_404);
nand U568 (N_568,N_124,N_204);
nand U569 (N_569,N_41,N_387);
and U570 (N_570,N_94,N_476);
and U571 (N_571,N_98,N_449);
nor U572 (N_572,N_254,N_286);
or U573 (N_573,N_210,N_325);
nand U574 (N_574,N_412,N_399);
xor U575 (N_575,N_150,N_431);
nand U576 (N_576,N_164,N_381);
or U577 (N_577,N_310,N_107);
xnor U578 (N_578,N_321,N_279);
or U579 (N_579,N_55,N_154);
nor U580 (N_580,N_9,N_466);
and U581 (N_581,N_346,N_423);
xnor U582 (N_582,N_277,N_26);
xnor U583 (N_583,N_196,N_261);
nor U584 (N_584,N_340,N_201);
and U585 (N_585,N_168,N_125);
xnor U586 (N_586,N_263,N_253);
xor U587 (N_587,N_495,N_488);
xor U588 (N_588,N_329,N_446);
xor U589 (N_589,N_32,N_409);
and U590 (N_590,N_156,N_183);
nor U591 (N_591,N_68,N_186);
and U592 (N_592,N_35,N_80);
or U593 (N_593,N_287,N_93);
xor U594 (N_594,N_289,N_461);
nor U595 (N_595,N_155,N_222);
or U596 (N_596,N_13,N_58);
and U597 (N_597,N_195,N_485);
or U598 (N_598,N_486,N_184);
or U599 (N_599,N_378,N_443);
or U600 (N_600,N_34,N_23);
nand U601 (N_601,N_478,N_102);
or U602 (N_602,N_389,N_20);
nor U603 (N_603,N_402,N_406);
and U604 (N_604,N_309,N_172);
nand U605 (N_605,N_288,N_84);
nor U606 (N_606,N_252,N_63);
nor U607 (N_607,N_371,N_118);
or U608 (N_608,N_67,N_305);
and U609 (N_609,N_293,N_149);
nand U610 (N_610,N_73,N_379);
xor U611 (N_611,N_330,N_284);
and U612 (N_612,N_262,N_364);
and U613 (N_613,N_322,N_472);
nand U614 (N_614,N_460,N_78);
and U615 (N_615,N_165,N_484);
and U616 (N_616,N_127,N_211);
nand U617 (N_617,N_161,N_123);
and U618 (N_618,N_173,N_7);
xnor U619 (N_619,N_447,N_352);
and U620 (N_620,N_437,N_440);
or U621 (N_621,N_335,N_248);
or U622 (N_622,N_10,N_185);
nand U623 (N_623,N_223,N_105);
nand U624 (N_624,N_442,N_392);
nor U625 (N_625,N_114,N_87);
and U626 (N_626,N_415,N_327);
nand U627 (N_627,N_297,N_16);
xor U628 (N_628,N_56,N_295);
or U629 (N_629,N_332,N_193);
nand U630 (N_630,N_54,N_17);
xor U631 (N_631,N_405,N_479);
xor U632 (N_632,N_22,N_111);
xnor U633 (N_633,N_280,N_454);
or U634 (N_634,N_72,N_197);
xor U635 (N_635,N_380,N_192);
nand U636 (N_636,N_231,N_351);
or U637 (N_637,N_413,N_75);
nor U638 (N_638,N_131,N_213);
or U639 (N_639,N_498,N_383);
nand U640 (N_640,N_122,N_151);
or U641 (N_641,N_91,N_64);
or U642 (N_642,N_134,N_489);
nor U643 (N_643,N_417,N_450);
nand U644 (N_644,N_353,N_421);
xor U645 (N_645,N_3,N_283);
or U646 (N_646,N_336,N_312);
nand U647 (N_647,N_467,N_224);
xor U648 (N_648,N_314,N_304);
nor U649 (N_649,N_130,N_33);
nand U650 (N_650,N_112,N_333);
and U651 (N_651,N_359,N_490);
nand U652 (N_652,N_6,N_171);
xnor U653 (N_653,N_24,N_227);
or U654 (N_654,N_411,N_434);
or U655 (N_655,N_348,N_376);
nor U656 (N_656,N_89,N_265);
and U657 (N_657,N_438,N_422);
nand U658 (N_658,N_394,N_175);
nand U659 (N_659,N_338,N_65);
nor U660 (N_660,N_237,N_96);
xor U661 (N_661,N_269,N_37);
nor U662 (N_662,N_382,N_31);
xnor U663 (N_663,N_448,N_361);
or U664 (N_664,N_469,N_470);
nor U665 (N_665,N_21,N_355);
and U666 (N_666,N_153,N_12);
and U667 (N_667,N_303,N_187);
or U668 (N_668,N_285,N_229);
xnor U669 (N_669,N_167,N_77);
and U670 (N_670,N_174,N_499);
nand U671 (N_671,N_319,N_15);
or U672 (N_672,N_483,N_444);
or U673 (N_673,N_272,N_426);
nor U674 (N_674,N_138,N_189);
and U675 (N_675,N_29,N_39);
xor U676 (N_676,N_129,N_148);
nor U677 (N_677,N_147,N_492);
or U678 (N_678,N_281,N_292);
and U679 (N_679,N_317,N_339);
or U680 (N_680,N_38,N_416);
and U681 (N_681,N_42,N_459);
nor U682 (N_682,N_424,N_207);
nand U683 (N_683,N_208,N_1);
nand U684 (N_684,N_487,N_40);
or U685 (N_685,N_428,N_61);
or U686 (N_686,N_436,N_331);
nand U687 (N_687,N_206,N_328);
nor U688 (N_688,N_241,N_11);
or U689 (N_689,N_465,N_414);
nor U690 (N_690,N_158,N_247);
and U691 (N_691,N_200,N_230);
and U692 (N_692,N_119,N_205);
and U693 (N_693,N_88,N_273);
or U694 (N_694,N_278,N_251);
xnor U695 (N_695,N_142,N_258);
or U696 (N_696,N_139,N_393);
xor U697 (N_697,N_496,N_396);
or U698 (N_698,N_8,N_323);
or U699 (N_699,N_307,N_365);
and U700 (N_700,N_27,N_264);
xnor U701 (N_701,N_372,N_427);
xnor U702 (N_702,N_410,N_290);
nor U703 (N_703,N_14,N_86);
nor U704 (N_704,N_234,N_311);
xnor U705 (N_705,N_239,N_169);
nand U706 (N_706,N_30,N_474);
and U707 (N_707,N_19,N_362);
and U708 (N_708,N_52,N_267);
nor U709 (N_709,N_145,N_212);
and U710 (N_710,N_51,N_121);
and U711 (N_711,N_140,N_384);
or U712 (N_712,N_120,N_199);
or U713 (N_713,N_76,N_433);
nand U714 (N_714,N_301,N_83);
xor U715 (N_715,N_354,N_217);
xnor U716 (N_716,N_315,N_473);
nor U717 (N_717,N_480,N_70);
xor U718 (N_718,N_345,N_370);
or U719 (N_719,N_46,N_441);
or U720 (N_720,N_497,N_194);
or U721 (N_721,N_407,N_115);
and U722 (N_722,N_188,N_5);
xor U723 (N_723,N_318,N_452);
nand U724 (N_724,N_225,N_275);
or U725 (N_725,N_373,N_435);
nor U726 (N_726,N_398,N_226);
nor U727 (N_727,N_250,N_456);
xor U728 (N_728,N_257,N_228);
nand U729 (N_729,N_429,N_159);
nor U730 (N_730,N_90,N_233);
or U731 (N_731,N_420,N_397);
nor U732 (N_732,N_97,N_432);
and U733 (N_733,N_216,N_299);
xor U734 (N_734,N_294,N_106);
xnor U735 (N_735,N_43,N_144);
xnor U736 (N_736,N_368,N_276);
and U737 (N_737,N_181,N_53);
nor U738 (N_738,N_100,N_218);
nor U739 (N_739,N_109,N_82);
xor U740 (N_740,N_418,N_190);
or U741 (N_741,N_62,N_137);
nand U742 (N_742,N_202,N_298);
and U743 (N_743,N_50,N_390);
or U744 (N_744,N_266,N_491);
xnor U745 (N_745,N_182,N_430);
xnor U746 (N_746,N_85,N_209);
nand U747 (N_747,N_313,N_357);
nand U748 (N_748,N_282,N_462);
xnor U749 (N_749,N_374,N_128);
nor U750 (N_750,N_330,N_355);
or U751 (N_751,N_421,N_215);
nor U752 (N_752,N_362,N_285);
and U753 (N_753,N_414,N_45);
nand U754 (N_754,N_330,N_421);
or U755 (N_755,N_461,N_207);
or U756 (N_756,N_173,N_405);
or U757 (N_757,N_124,N_337);
xnor U758 (N_758,N_127,N_117);
and U759 (N_759,N_338,N_31);
nand U760 (N_760,N_140,N_110);
xnor U761 (N_761,N_346,N_384);
xnor U762 (N_762,N_364,N_99);
nor U763 (N_763,N_57,N_331);
or U764 (N_764,N_466,N_298);
and U765 (N_765,N_379,N_324);
xor U766 (N_766,N_93,N_234);
nand U767 (N_767,N_60,N_116);
xor U768 (N_768,N_497,N_5);
or U769 (N_769,N_58,N_467);
or U770 (N_770,N_205,N_212);
nor U771 (N_771,N_84,N_453);
xor U772 (N_772,N_176,N_172);
xor U773 (N_773,N_291,N_216);
or U774 (N_774,N_19,N_417);
xor U775 (N_775,N_491,N_123);
nand U776 (N_776,N_496,N_285);
nand U777 (N_777,N_73,N_136);
nand U778 (N_778,N_5,N_291);
nor U779 (N_779,N_131,N_238);
or U780 (N_780,N_316,N_420);
xor U781 (N_781,N_241,N_238);
nand U782 (N_782,N_148,N_276);
or U783 (N_783,N_397,N_427);
xor U784 (N_784,N_349,N_23);
or U785 (N_785,N_361,N_9);
or U786 (N_786,N_39,N_290);
nor U787 (N_787,N_260,N_219);
xor U788 (N_788,N_434,N_437);
and U789 (N_789,N_364,N_148);
nor U790 (N_790,N_307,N_438);
xor U791 (N_791,N_486,N_249);
or U792 (N_792,N_274,N_142);
xor U793 (N_793,N_432,N_44);
xor U794 (N_794,N_496,N_365);
and U795 (N_795,N_275,N_487);
or U796 (N_796,N_460,N_445);
or U797 (N_797,N_168,N_231);
nor U798 (N_798,N_14,N_78);
xnor U799 (N_799,N_263,N_206);
nand U800 (N_800,N_417,N_233);
xnor U801 (N_801,N_355,N_120);
nand U802 (N_802,N_290,N_158);
nand U803 (N_803,N_243,N_50);
or U804 (N_804,N_459,N_26);
or U805 (N_805,N_375,N_109);
xor U806 (N_806,N_17,N_42);
or U807 (N_807,N_266,N_102);
nand U808 (N_808,N_374,N_444);
nor U809 (N_809,N_299,N_354);
nand U810 (N_810,N_211,N_130);
or U811 (N_811,N_307,N_136);
or U812 (N_812,N_274,N_71);
nand U813 (N_813,N_443,N_58);
nor U814 (N_814,N_473,N_104);
or U815 (N_815,N_337,N_403);
nand U816 (N_816,N_261,N_186);
nand U817 (N_817,N_368,N_421);
and U818 (N_818,N_242,N_192);
and U819 (N_819,N_233,N_207);
nand U820 (N_820,N_123,N_53);
xor U821 (N_821,N_351,N_387);
or U822 (N_822,N_31,N_367);
nand U823 (N_823,N_267,N_113);
xnor U824 (N_824,N_347,N_98);
xor U825 (N_825,N_261,N_471);
or U826 (N_826,N_449,N_409);
nor U827 (N_827,N_168,N_321);
or U828 (N_828,N_213,N_415);
xor U829 (N_829,N_98,N_71);
xnor U830 (N_830,N_21,N_286);
and U831 (N_831,N_175,N_390);
nand U832 (N_832,N_469,N_147);
nand U833 (N_833,N_37,N_366);
xnor U834 (N_834,N_194,N_140);
or U835 (N_835,N_254,N_455);
and U836 (N_836,N_33,N_434);
or U837 (N_837,N_319,N_205);
nand U838 (N_838,N_14,N_113);
nand U839 (N_839,N_280,N_180);
or U840 (N_840,N_286,N_131);
and U841 (N_841,N_253,N_271);
or U842 (N_842,N_445,N_348);
nor U843 (N_843,N_297,N_191);
nor U844 (N_844,N_132,N_241);
and U845 (N_845,N_383,N_402);
nor U846 (N_846,N_85,N_233);
or U847 (N_847,N_360,N_55);
or U848 (N_848,N_278,N_317);
and U849 (N_849,N_302,N_347);
and U850 (N_850,N_130,N_290);
nor U851 (N_851,N_119,N_437);
or U852 (N_852,N_30,N_253);
xor U853 (N_853,N_39,N_407);
nor U854 (N_854,N_308,N_400);
nor U855 (N_855,N_65,N_220);
nand U856 (N_856,N_339,N_33);
xnor U857 (N_857,N_442,N_283);
xnor U858 (N_858,N_257,N_308);
xnor U859 (N_859,N_393,N_452);
nor U860 (N_860,N_263,N_422);
and U861 (N_861,N_281,N_270);
nor U862 (N_862,N_377,N_481);
and U863 (N_863,N_224,N_352);
xor U864 (N_864,N_90,N_182);
or U865 (N_865,N_314,N_76);
nor U866 (N_866,N_150,N_183);
nor U867 (N_867,N_27,N_108);
or U868 (N_868,N_362,N_286);
xnor U869 (N_869,N_24,N_191);
xnor U870 (N_870,N_412,N_308);
and U871 (N_871,N_261,N_361);
and U872 (N_872,N_460,N_17);
nor U873 (N_873,N_122,N_464);
xnor U874 (N_874,N_176,N_489);
nor U875 (N_875,N_35,N_99);
nor U876 (N_876,N_5,N_62);
or U877 (N_877,N_3,N_223);
nand U878 (N_878,N_326,N_229);
xnor U879 (N_879,N_479,N_163);
nand U880 (N_880,N_450,N_463);
and U881 (N_881,N_100,N_389);
or U882 (N_882,N_140,N_58);
or U883 (N_883,N_467,N_107);
or U884 (N_884,N_105,N_470);
xnor U885 (N_885,N_175,N_391);
or U886 (N_886,N_87,N_470);
nor U887 (N_887,N_388,N_489);
or U888 (N_888,N_418,N_133);
or U889 (N_889,N_363,N_49);
xor U890 (N_890,N_130,N_297);
xnor U891 (N_891,N_148,N_78);
or U892 (N_892,N_347,N_116);
nor U893 (N_893,N_366,N_483);
nor U894 (N_894,N_282,N_213);
xor U895 (N_895,N_276,N_223);
and U896 (N_896,N_84,N_348);
nand U897 (N_897,N_117,N_341);
nand U898 (N_898,N_451,N_294);
and U899 (N_899,N_371,N_398);
xnor U900 (N_900,N_488,N_497);
and U901 (N_901,N_202,N_328);
nor U902 (N_902,N_155,N_495);
and U903 (N_903,N_56,N_319);
nor U904 (N_904,N_0,N_231);
nand U905 (N_905,N_389,N_290);
xnor U906 (N_906,N_310,N_177);
xnor U907 (N_907,N_452,N_29);
and U908 (N_908,N_404,N_91);
or U909 (N_909,N_330,N_5);
xor U910 (N_910,N_48,N_269);
nand U911 (N_911,N_16,N_90);
nand U912 (N_912,N_223,N_482);
xnor U913 (N_913,N_498,N_402);
xor U914 (N_914,N_293,N_101);
nand U915 (N_915,N_348,N_14);
and U916 (N_916,N_498,N_434);
and U917 (N_917,N_339,N_10);
nor U918 (N_918,N_454,N_417);
nor U919 (N_919,N_179,N_117);
nand U920 (N_920,N_111,N_452);
xor U921 (N_921,N_110,N_377);
or U922 (N_922,N_323,N_209);
or U923 (N_923,N_419,N_322);
nor U924 (N_924,N_83,N_249);
and U925 (N_925,N_374,N_427);
nor U926 (N_926,N_385,N_477);
and U927 (N_927,N_87,N_490);
nand U928 (N_928,N_377,N_155);
xor U929 (N_929,N_420,N_359);
nand U930 (N_930,N_185,N_69);
and U931 (N_931,N_350,N_106);
or U932 (N_932,N_286,N_339);
nand U933 (N_933,N_255,N_325);
and U934 (N_934,N_389,N_297);
nor U935 (N_935,N_364,N_494);
nand U936 (N_936,N_308,N_170);
nor U937 (N_937,N_315,N_431);
and U938 (N_938,N_187,N_10);
nor U939 (N_939,N_130,N_240);
nor U940 (N_940,N_300,N_185);
and U941 (N_941,N_383,N_477);
nand U942 (N_942,N_450,N_435);
or U943 (N_943,N_473,N_368);
or U944 (N_944,N_499,N_415);
or U945 (N_945,N_479,N_309);
nand U946 (N_946,N_102,N_169);
nand U947 (N_947,N_297,N_152);
nor U948 (N_948,N_186,N_104);
nand U949 (N_949,N_214,N_42);
nand U950 (N_950,N_26,N_137);
nand U951 (N_951,N_116,N_307);
xor U952 (N_952,N_327,N_471);
nor U953 (N_953,N_454,N_392);
and U954 (N_954,N_468,N_132);
or U955 (N_955,N_74,N_352);
nand U956 (N_956,N_306,N_484);
nor U957 (N_957,N_293,N_160);
nor U958 (N_958,N_7,N_273);
or U959 (N_959,N_165,N_335);
and U960 (N_960,N_353,N_40);
and U961 (N_961,N_393,N_6);
nand U962 (N_962,N_129,N_141);
nor U963 (N_963,N_67,N_109);
or U964 (N_964,N_47,N_57);
or U965 (N_965,N_483,N_72);
and U966 (N_966,N_428,N_456);
and U967 (N_967,N_420,N_33);
xor U968 (N_968,N_281,N_342);
xor U969 (N_969,N_138,N_334);
nor U970 (N_970,N_155,N_11);
or U971 (N_971,N_165,N_65);
nand U972 (N_972,N_289,N_193);
nor U973 (N_973,N_335,N_163);
xnor U974 (N_974,N_357,N_242);
or U975 (N_975,N_264,N_218);
and U976 (N_976,N_288,N_360);
and U977 (N_977,N_334,N_291);
nor U978 (N_978,N_287,N_31);
or U979 (N_979,N_335,N_44);
nor U980 (N_980,N_203,N_172);
nand U981 (N_981,N_119,N_171);
xnor U982 (N_982,N_381,N_202);
nor U983 (N_983,N_254,N_495);
xnor U984 (N_984,N_76,N_336);
xor U985 (N_985,N_176,N_226);
or U986 (N_986,N_97,N_446);
xnor U987 (N_987,N_204,N_316);
and U988 (N_988,N_410,N_352);
and U989 (N_989,N_161,N_480);
or U990 (N_990,N_393,N_441);
nor U991 (N_991,N_423,N_164);
and U992 (N_992,N_299,N_427);
nand U993 (N_993,N_436,N_157);
xor U994 (N_994,N_85,N_119);
and U995 (N_995,N_26,N_128);
or U996 (N_996,N_470,N_70);
or U997 (N_997,N_254,N_80);
nor U998 (N_998,N_307,N_178);
nor U999 (N_999,N_396,N_329);
nand U1000 (N_1000,N_805,N_891);
or U1001 (N_1001,N_621,N_853);
nand U1002 (N_1002,N_749,N_708);
xnor U1003 (N_1003,N_548,N_847);
xnor U1004 (N_1004,N_961,N_850);
nand U1005 (N_1005,N_661,N_768);
nand U1006 (N_1006,N_818,N_945);
nand U1007 (N_1007,N_523,N_792);
or U1008 (N_1008,N_518,N_529);
and U1009 (N_1009,N_758,N_726);
nand U1010 (N_1010,N_806,N_832);
xor U1011 (N_1011,N_907,N_838);
nor U1012 (N_1012,N_900,N_807);
and U1013 (N_1013,N_931,N_755);
xnor U1014 (N_1014,N_656,N_982);
nand U1015 (N_1015,N_941,N_845);
and U1016 (N_1016,N_546,N_933);
and U1017 (N_1017,N_700,N_864);
and U1018 (N_1018,N_667,N_738);
xnor U1019 (N_1019,N_851,N_544);
or U1020 (N_1020,N_728,N_837);
xor U1021 (N_1021,N_731,N_831);
or U1022 (N_1022,N_815,N_684);
or U1023 (N_1023,N_527,N_710);
xor U1024 (N_1024,N_742,N_631);
nand U1025 (N_1025,N_522,N_826);
nor U1026 (N_1026,N_926,N_670);
and U1027 (N_1027,N_735,N_510);
and U1028 (N_1028,N_689,N_607);
nor U1029 (N_1029,N_543,N_812);
xnor U1030 (N_1030,N_617,N_743);
or U1031 (N_1031,N_757,N_965);
nand U1032 (N_1032,N_869,N_545);
xor U1033 (N_1033,N_683,N_587);
and U1034 (N_1034,N_777,N_620);
or U1035 (N_1035,N_686,N_939);
xnor U1036 (N_1036,N_551,N_693);
xnor U1037 (N_1037,N_886,N_990);
or U1038 (N_1038,N_882,N_761);
nand U1039 (N_1039,N_764,N_935);
and U1040 (N_1040,N_920,N_930);
and U1041 (N_1041,N_912,N_740);
and U1042 (N_1042,N_873,N_919);
xor U1043 (N_1043,N_553,N_950);
and U1044 (N_1044,N_730,N_594);
and U1045 (N_1045,N_592,N_820);
xor U1046 (N_1046,N_707,N_947);
nor U1047 (N_1047,N_713,N_836);
and U1048 (N_1048,N_765,N_937);
nor U1049 (N_1049,N_517,N_896);
and U1050 (N_1050,N_802,N_974);
and U1051 (N_1051,N_558,N_932);
or U1052 (N_1052,N_664,N_663);
nand U1053 (N_1053,N_817,N_923);
and U1054 (N_1054,N_719,N_879);
and U1055 (N_1055,N_784,N_632);
xor U1056 (N_1056,N_789,N_659);
nor U1057 (N_1057,N_692,N_840);
xor U1058 (N_1058,N_960,N_952);
or U1059 (N_1059,N_734,N_622);
nor U1060 (N_1060,N_903,N_775);
or U1061 (N_1061,N_550,N_998);
nand U1062 (N_1062,N_598,N_662);
and U1063 (N_1063,N_911,N_858);
xor U1064 (N_1064,N_701,N_729);
or U1065 (N_1065,N_898,N_916);
nand U1066 (N_1066,N_557,N_613);
nor U1067 (N_1067,N_855,N_660);
nand U1068 (N_1068,N_590,N_841);
xnor U1069 (N_1069,N_893,N_991);
nor U1070 (N_1070,N_653,N_530);
xnor U1071 (N_1071,N_681,N_872);
and U1072 (N_1072,N_630,N_509);
nor U1073 (N_1073,N_819,N_574);
and U1074 (N_1074,N_672,N_500);
and U1075 (N_1075,N_508,N_650);
and U1076 (N_1076,N_781,N_671);
or U1077 (N_1077,N_636,N_536);
or U1078 (N_1078,N_801,N_868);
nand U1079 (N_1079,N_969,N_793);
and U1080 (N_1080,N_834,N_605);
nand U1081 (N_1081,N_588,N_843);
xnor U1082 (N_1082,N_526,N_910);
and U1083 (N_1083,N_624,N_967);
or U1084 (N_1084,N_721,N_582);
xnor U1085 (N_1085,N_501,N_874);
xnor U1086 (N_1086,N_634,N_609);
nor U1087 (N_1087,N_674,N_778);
nand U1088 (N_1088,N_814,N_637);
or U1089 (N_1089,N_809,N_563);
nand U1090 (N_1090,N_779,N_810);
nand U1091 (N_1091,N_943,N_769);
or U1092 (N_1092,N_828,N_720);
or U1093 (N_1093,N_862,N_601);
nand U1094 (N_1094,N_676,N_573);
or U1095 (N_1095,N_655,N_995);
nor U1096 (N_1096,N_766,N_575);
nand U1097 (N_1097,N_669,N_954);
and U1098 (N_1098,N_914,N_964);
nand U1099 (N_1099,N_959,N_860);
xor U1100 (N_1100,N_983,N_762);
nand U1101 (N_1101,N_569,N_830);
nor U1102 (N_1102,N_880,N_559);
or U1103 (N_1103,N_870,N_725);
and U1104 (N_1104,N_854,N_895);
and U1105 (N_1105,N_875,N_540);
nand U1106 (N_1106,N_606,N_507);
or U1107 (N_1107,N_816,N_827);
xnor U1108 (N_1108,N_984,N_652);
nor U1109 (N_1109,N_852,N_541);
nor U1110 (N_1110,N_780,N_736);
nand U1111 (N_1111,N_866,N_716);
nand U1112 (N_1112,N_562,N_856);
nor U1113 (N_1113,N_963,N_748);
and U1114 (N_1114,N_744,N_901);
xnor U1115 (N_1115,N_584,N_904);
or U1116 (N_1116,N_773,N_822);
nand U1117 (N_1117,N_833,N_798);
xor U1118 (N_1118,N_786,N_994);
nor U1119 (N_1119,N_796,N_657);
or U1120 (N_1120,N_846,N_724);
nand U1121 (N_1121,N_682,N_648);
xnor U1122 (N_1122,N_934,N_608);
and U1123 (N_1123,N_532,N_953);
nand U1124 (N_1124,N_596,N_927);
and U1125 (N_1125,N_889,N_804);
nor U1126 (N_1126,N_987,N_694);
nor U1127 (N_1127,N_884,N_679);
nand U1128 (N_1128,N_715,N_811);
or U1129 (N_1129,N_938,N_723);
xor U1130 (N_1130,N_703,N_752);
or U1131 (N_1131,N_610,N_695);
nor U1132 (N_1132,N_973,N_772);
and U1133 (N_1133,N_942,N_929);
nor U1134 (N_1134,N_746,N_909);
xor U1135 (N_1135,N_503,N_842);
or U1136 (N_1136,N_917,N_638);
nor U1137 (N_1137,N_745,N_625);
nor U1138 (N_1138,N_774,N_839);
and U1139 (N_1139,N_794,N_698);
and U1140 (N_1140,N_712,N_576);
and U1141 (N_1141,N_589,N_504);
nand U1142 (N_1142,N_999,N_554);
nor U1143 (N_1143,N_642,N_883);
xor U1144 (N_1144,N_711,N_565);
and U1145 (N_1145,N_640,N_612);
or U1146 (N_1146,N_788,N_673);
and U1147 (N_1147,N_922,N_787);
nor U1148 (N_1148,N_603,N_611);
xnor U1149 (N_1149,N_646,N_865);
nand U1150 (N_1150,N_892,N_966);
and U1151 (N_1151,N_813,N_680);
nor U1152 (N_1152,N_525,N_581);
xor U1153 (N_1153,N_844,N_519);
nand U1154 (N_1154,N_675,N_633);
nand U1155 (N_1155,N_600,N_685);
and U1156 (N_1156,N_580,N_829);
or U1157 (N_1157,N_702,N_595);
nor U1158 (N_1158,N_754,N_705);
nor U1159 (N_1159,N_717,N_785);
nand U1160 (N_1160,N_876,N_531);
xor U1161 (N_1161,N_528,N_668);
or U1162 (N_1162,N_968,N_678);
or U1163 (N_1163,N_714,N_513);
nand U1164 (N_1164,N_997,N_956);
nand U1165 (N_1165,N_645,N_951);
or U1166 (N_1166,N_666,N_552);
nand U1167 (N_1167,N_549,N_859);
and U1168 (N_1168,N_972,N_928);
nor U1169 (N_1169,N_626,N_616);
xnor U1170 (N_1170,N_718,N_516);
nand U1171 (N_1171,N_515,N_514);
xor U1172 (N_1172,N_770,N_771);
and U1173 (N_1173,N_512,N_753);
or U1174 (N_1174,N_696,N_913);
xnor U1175 (N_1175,N_795,N_560);
xor U1176 (N_1176,N_857,N_722);
nor U1177 (N_1177,N_849,N_727);
xor U1178 (N_1178,N_647,N_741);
xor U1179 (N_1179,N_591,N_732);
nand U1180 (N_1180,N_782,N_848);
or U1181 (N_1181,N_586,N_691);
and U1182 (N_1182,N_690,N_665);
or U1183 (N_1183,N_906,N_975);
nand U1184 (N_1184,N_538,N_767);
nor U1185 (N_1185,N_555,N_988);
and U1186 (N_1186,N_957,N_733);
or U1187 (N_1187,N_924,N_567);
nand U1188 (N_1188,N_750,N_791);
nor U1189 (N_1189,N_888,N_905);
or U1190 (N_1190,N_980,N_948);
xnor U1191 (N_1191,N_627,N_800);
and U1192 (N_1192,N_566,N_955);
nor U1193 (N_1193,N_658,N_604);
and U1194 (N_1194,N_643,N_881);
or U1195 (N_1195,N_824,N_783);
and U1196 (N_1196,N_654,N_902);
nand U1197 (N_1197,N_688,N_564);
nand U1198 (N_1198,N_602,N_887);
and U1199 (N_1199,N_949,N_547);
nand U1200 (N_1200,N_709,N_585);
or U1201 (N_1201,N_537,N_577);
and U1202 (N_1202,N_885,N_521);
xnor U1203 (N_1203,N_985,N_760);
or U1204 (N_1204,N_572,N_897);
and U1205 (N_1205,N_561,N_986);
nand U1206 (N_1206,N_506,N_799);
or U1207 (N_1207,N_803,N_597);
nand U1208 (N_1208,N_992,N_520);
nor U1209 (N_1209,N_556,N_977);
nor U1210 (N_1210,N_918,N_583);
or U1211 (N_1211,N_511,N_534);
xor U1212 (N_1212,N_699,N_970);
nor U1213 (N_1213,N_524,N_790);
nor U1214 (N_1214,N_635,N_776);
and U1215 (N_1215,N_505,N_867);
or U1216 (N_1216,N_808,N_871);
nand U1217 (N_1217,N_542,N_940);
and U1218 (N_1218,N_877,N_677);
nand U1219 (N_1219,N_976,N_944);
xnor U1220 (N_1220,N_539,N_946);
nand U1221 (N_1221,N_502,N_861);
xor U1222 (N_1222,N_568,N_639);
nand U1223 (N_1223,N_925,N_644);
nand U1224 (N_1224,N_649,N_962);
nor U1225 (N_1225,N_825,N_981);
nand U1226 (N_1226,N_570,N_618);
and U1227 (N_1227,N_958,N_593);
xor U1228 (N_1228,N_993,N_894);
or U1229 (N_1229,N_614,N_651);
nand U1230 (N_1230,N_890,N_706);
or U1231 (N_1231,N_687,N_747);
or U1232 (N_1232,N_979,N_629);
or U1233 (N_1233,N_641,N_823);
nor U1234 (N_1234,N_978,N_915);
nor U1235 (N_1235,N_533,N_737);
nor U1236 (N_1236,N_835,N_623);
nand U1237 (N_1237,N_821,N_615);
xor U1238 (N_1238,N_863,N_899);
and U1239 (N_1239,N_878,N_751);
or U1240 (N_1240,N_619,N_756);
nor U1241 (N_1241,N_599,N_989);
nor U1242 (N_1242,N_628,N_739);
or U1243 (N_1243,N_535,N_759);
nand U1244 (N_1244,N_936,N_971);
xor U1245 (N_1245,N_763,N_697);
xnor U1246 (N_1246,N_797,N_704);
nand U1247 (N_1247,N_921,N_578);
and U1248 (N_1248,N_908,N_571);
and U1249 (N_1249,N_996,N_579);
nand U1250 (N_1250,N_643,N_835);
nand U1251 (N_1251,N_579,N_503);
xnor U1252 (N_1252,N_635,N_563);
and U1253 (N_1253,N_661,N_526);
nand U1254 (N_1254,N_718,N_624);
xnor U1255 (N_1255,N_589,N_832);
xnor U1256 (N_1256,N_696,N_952);
nand U1257 (N_1257,N_787,N_853);
xor U1258 (N_1258,N_730,N_690);
nand U1259 (N_1259,N_586,N_595);
and U1260 (N_1260,N_795,N_926);
nor U1261 (N_1261,N_892,N_517);
or U1262 (N_1262,N_679,N_572);
nor U1263 (N_1263,N_786,N_662);
nor U1264 (N_1264,N_761,N_886);
and U1265 (N_1265,N_501,N_694);
and U1266 (N_1266,N_662,N_560);
or U1267 (N_1267,N_611,N_676);
nor U1268 (N_1268,N_524,N_715);
and U1269 (N_1269,N_665,N_621);
nand U1270 (N_1270,N_824,N_853);
or U1271 (N_1271,N_590,N_974);
nand U1272 (N_1272,N_516,N_907);
or U1273 (N_1273,N_926,N_721);
or U1274 (N_1274,N_836,N_732);
or U1275 (N_1275,N_736,N_583);
xor U1276 (N_1276,N_686,N_891);
nand U1277 (N_1277,N_797,N_535);
and U1278 (N_1278,N_551,N_902);
or U1279 (N_1279,N_934,N_984);
nand U1280 (N_1280,N_825,N_884);
xor U1281 (N_1281,N_637,N_729);
nor U1282 (N_1282,N_825,N_639);
xor U1283 (N_1283,N_916,N_773);
xor U1284 (N_1284,N_835,N_708);
nor U1285 (N_1285,N_616,N_588);
or U1286 (N_1286,N_513,N_813);
xor U1287 (N_1287,N_795,N_937);
nor U1288 (N_1288,N_503,N_820);
xor U1289 (N_1289,N_761,N_939);
nor U1290 (N_1290,N_750,N_557);
xor U1291 (N_1291,N_552,N_886);
nand U1292 (N_1292,N_792,N_682);
nor U1293 (N_1293,N_501,N_808);
nand U1294 (N_1294,N_786,N_501);
xor U1295 (N_1295,N_959,N_783);
xor U1296 (N_1296,N_703,N_827);
xnor U1297 (N_1297,N_965,N_619);
nor U1298 (N_1298,N_605,N_744);
or U1299 (N_1299,N_715,N_858);
nor U1300 (N_1300,N_872,N_568);
and U1301 (N_1301,N_559,N_813);
xnor U1302 (N_1302,N_843,N_700);
nor U1303 (N_1303,N_883,N_898);
nor U1304 (N_1304,N_861,N_552);
nand U1305 (N_1305,N_767,N_826);
xor U1306 (N_1306,N_653,N_825);
or U1307 (N_1307,N_608,N_631);
and U1308 (N_1308,N_677,N_538);
nor U1309 (N_1309,N_767,N_520);
or U1310 (N_1310,N_566,N_788);
and U1311 (N_1311,N_809,N_863);
and U1312 (N_1312,N_515,N_903);
nand U1313 (N_1313,N_520,N_581);
xnor U1314 (N_1314,N_521,N_721);
xor U1315 (N_1315,N_777,N_692);
nand U1316 (N_1316,N_849,N_716);
xor U1317 (N_1317,N_811,N_798);
nor U1318 (N_1318,N_564,N_717);
nor U1319 (N_1319,N_595,N_521);
nand U1320 (N_1320,N_578,N_837);
nand U1321 (N_1321,N_623,N_942);
and U1322 (N_1322,N_583,N_672);
nand U1323 (N_1323,N_817,N_674);
or U1324 (N_1324,N_701,N_570);
xor U1325 (N_1325,N_716,N_795);
xnor U1326 (N_1326,N_578,N_544);
nor U1327 (N_1327,N_793,N_802);
nand U1328 (N_1328,N_589,N_572);
nand U1329 (N_1329,N_534,N_576);
nand U1330 (N_1330,N_910,N_685);
nor U1331 (N_1331,N_929,N_620);
xor U1332 (N_1332,N_569,N_867);
and U1333 (N_1333,N_871,N_548);
and U1334 (N_1334,N_929,N_506);
nor U1335 (N_1335,N_966,N_924);
xor U1336 (N_1336,N_924,N_962);
nor U1337 (N_1337,N_607,N_559);
nor U1338 (N_1338,N_815,N_642);
nor U1339 (N_1339,N_922,N_572);
or U1340 (N_1340,N_737,N_877);
nand U1341 (N_1341,N_749,N_958);
xnor U1342 (N_1342,N_558,N_642);
nand U1343 (N_1343,N_593,N_979);
or U1344 (N_1344,N_643,N_539);
or U1345 (N_1345,N_853,N_989);
and U1346 (N_1346,N_646,N_631);
xor U1347 (N_1347,N_790,N_800);
and U1348 (N_1348,N_559,N_973);
or U1349 (N_1349,N_949,N_574);
and U1350 (N_1350,N_904,N_927);
or U1351 (N_1351,N_587,N_758);
xnor U1352 (N_1352,N_887,N_895);
and U1353 (N_1353,N_698,N_526);
or U1354 (N_1354,N_961,N_794);
xnor U1355 (N_1355,N_881,N_630);
or U1356 (N_1356,N_948,N_957);
nor U1357 (N_1357,N_838,N_686);
or U1358 (N_1358,N_520,N_843);
nand U1359 (N_1359,N_551,N_575);
or U1360 (N_1360,N_548,N_587);
nand U1361 (N_1361,N_679,N_787);
xnor U1362 (N_1362,N_990,N_511);
or U1363 (N_1363,N_631,N_670);
and U1364 (N_1364,N_644,N_629);
and U1365 (N_1365,N_773,N_771);
or U1366 (N_1366,N_882,N_923);
xor U1367 (N_1367,N_665,N_568);
or U1368 (N_1368,N_961,N_863);
nor U1369 (N_1369,N_886,N_714);
or U1370 (N_1370,N_580,N_659);
and U1371 (N_1371,N_864,N_693);
or U1372 (N_1372,N_984,N_996);
nand U1373 (N_1373,N_536,N_638);
and U1374 (N_1374,N_789,N_623);
xor U1375 (N_1375,N_665,N_777);
nor U1376 (N_1376,N_539,N_932);
or U1377 (N_1377,N_971,N_912);
xnor U1378 (N_1378,N_537,N_680);
or U1379 (N_1379,N_880,N_738);
nor U1380 (N_1380,N_661,N_739);
and U1381 (N_1381,N_621,N_672);
or U1382 (N_1382,N_546,N_892);
nand U1383 (N_1383,N_914,N_687);
and U1384 (N_1384,N_783,N_994);
nor U1385 (N_1385,N_838,N_812);
and U1386 (N_1386,N_686,N_834);
xor U1387 (N_1387,N_628,N_695);
and U1388 (N_1388,N_862,N_619);
or U1389 (N_1389,N_942,N_673);
nor U1390 (N_1390,N_532,N_688);
nand U1391 (N_1391,N_557,N_914);
nand U1392 (N_1392,N_611,N_873);
or U1393 (N_1393,N_590,N_605);
xnor U1394 (N_1394,N_723,N_631);
nor U1395 (N_1395,N_517,N_613);
and U1396 (N_1396,N_975,N_670);
nor U1397 (N_1397,N_753,N_628);
nand U1398 (N_1398,N_563,N_550);
nand U1399 (N_1399,N_588,N_548);
and U1400 (N_1400,N_635,N_679);
xnor U1401 (N_1401,N_632,N_862);
and U1402 (N_1402,N_969,N_708);
and U1403 (N_1403,N_888,N_724);
nand U1404 (N_1404,N_792,N_651);
or U1405 (N_1405,N_513,N_869);
or U1406 (N_1406,N_544,N_864);
nor U1407 (N_1407,N_921,N_766);
or U1408 (N_1408,N_974,N_636);
nor U1409 (N_1409,N_985,N_742);
nand U1410 (N_1410,N_870,N_592);
nand U1411 (N_1411,N_791,N_578);
xnor U1412 (N_1412,N_865,N_806);
and U1413 (N_1413,N_564,N_758);
xnor U1414 (N_1414,N_636,N_659);
xor U1415 (N_1415,N_783,N_738);
nand U1416 (N_1416,N_874,N_949);
nand U1417 (N_1417,N_813,N_924);
xor U1418 (N_1418,N_717,N_824);
nor U1419 (N_1419,N_524,N_862);
xor U1420 (N_1420,N_862,N_600);
nand U1421 (N_1421,N_619,N_849);
xnor U1422 (N_1422,N_572,N_880);
nor U1423 (N_1423,N_728,N_641);
nor U1424 (N_1424,N_913,N_862);
or U1425 (N_1425,N_928,N_694);
xnor U1426 (N_1426,N_879,N_673);
and U1427 (N_1427,N_859,N_683);
and U1428 (N_1428,N_603,N_526);
and U1429 (N_1429,N_544,N_792);
or U1430 (N_1430,N_700,N_930);
or U1431 (N_1431,N_786,N_754);
and U1432 (N_1432,N_760,N_881);
or U1433 (N_1433,N_610,N_869);
xor U1434 (N_1434,N_628,N_625);
nand U1435 (N_1435,N_682,N_921);
and U1436 (N_1436,N_540,N_764);
or U1437 (N_1437,N_783,N_511);
nand U1438 (N_1438,N_961,N_706);
nand U1439 (N_1439,N_568,N_683);
nor U1440 (N_1440,N_637,N_577);
and U1441 (N_1441,N_777,N_977);
and U1442 (N_1442,N_721,N_834);
or U1443 (N_1443,N_795,N_884);
nand U1444 (N_1444,N_545,N_851);
nand U1445 (N_1445,N_529,N_854);
nand U1446 (N_1446,N_614,N_598);
xnor U1447 (N_1447,N_544,N_681);
and U1448 (N_1448,N_710,N_740);
nand U1449 (N_1449,N_735,N_870);
or U1450 (N_1450,N_679,N_757);
xnor U1451 (N_1451,N_639,N_793);
xnor U1452 (N_1452,N_973,N_924);
or U1453 (N_1453,N_997,N_766);
or U1454 (N_1454,N_633,N_765);
nand U1455 (N_1455,N_763,N_602);
and U1456 (N_1456,N_886,N_706);
and U1457 (N_1457,N_565,N_780);
and U1458 (N_1458,N_797,N_996);
xnor U1459 (N_1459,N_752,N_503);
nor U1460 (N_1460,N_874,N_646);
xor U1461 (N_1461,N_875,N_909);
nor U1462 (N_1462,N_953,N_580);
or U1463 (N_1463,N_543,N_839);
nor U1464 (N_1464,N_595,N_775);
nand U1465 (N_1465,N_882,N_773);
nor U1466 (N_1466,N_910,N_909);
or U1467 (N_1467,N_921,N_510);
xor U1468 (N_1468,N_834,N_829);
nor U1469 (N_1469,N_972,N_784);
nand U1470 (N_1470,N_561,N_999);
nand U1471 (N_1471,N_698,N_613);
xnor U1472 (N_1472,N_907,N_760);
or U1473 (N_1473,N_733,N_597);
nand U1474 (N_1474,N_681,N_925);
nand U1475 (N_1475,N_843,N_771);
nor U1476 (N_1476,N_657,N_707);
or U1477 (N_1477,N_703,N_927);
and U1478 (N_1478,N_709,N_572);
or U1479 (N_1479,N_634,N_957);
nor U1480 (N_1480,N_787,N_646);
or U1481 (N_1481,N_859,N_782);
nor U1482 (N_1482,N_908,N_766);
or U1483 (N_1483,N_891,N_739);
xnor U1484 (N_1484,N_525,N_669);
or U1485 (N_1485,N_546,N_841);
nand U1486 (N_1486,N_939,N_715);
and U1487 (N_1487,N_981,N_882);
nor U1488 (N_1488,N_675,N_944);
or U1489 (N_1489,N_518,N_606);
and U1490 (N_1490,N_978,N_852);
nor U1491 (N_1491,N_741,N_554);
nor U1492 (N_1492,N_767,N_768);
nor U1493 (N_1493,N_572,N_566);
nand U1494 (N_1494,N_596,N_925);
xnor U1495 (N_1495,N_925,N_856);
nor U1496 (N_1496,N_995,N_725);
xor U1497 (N_1497,N_534,N_951);
nor U1498 (N_1498,N_848,N_619);
and U1499 (N_1499,N_776,N_605);
or U1500 (N_1500,N_1309,N_1256);
xnor U1501 (N_1501,N_1450,N_1091);
xor U1502 (N_1502,N_1164,N_1492);
nor U1503 (N_1503,N_1083,N_1000);
nor U1504 (N_1504,N_1004,N_1114);
nand U1505 (N_1505,N_1463,N_1145);
or U1506 (N_1506,N_1305,N_1404);
or U1507 (N_1507,N_1456,N_1345);
and U1508 (N_1508,N_1433,N_1316);
or U1509 (N_1509,N_1128,N_1082);
xnor U1510 (N_1510,N_1424,N_1179);
and U1511 (N_1511,N_1297,N_1076);
nand U1512 (N_1512,N_1488,N_1344);
or U1513 (N_1513,N_1471,N_1219);
xor U1514 (N_1514,N_1451,N_1234);
nand U1515 (N_1515,N_1363,N_1105);
and U1516 (N_1516,N_1079,N_1267);
or U1517 (N_1517,N_1360,N_1005);
and U1518 (N_1518,N_1125,N_1214);
nand U1519 (N_1519,N_1059,N_1428);
xor U1520 (N_1520,N_1330,N_1074);
nand U1521 (N_1521,N_1268,N_1474);
xor U1522 (N_1522,N_1314,N_1054);
and U1523 (N_1523,N_1047,N_1013);
nor U1524 (N_1524,N_1255,N_1092);
and U1525 (N_1525,N_1303,N_1045);
nand U1526 (N_1526,N_1044,N_1495);
xnor U1527 (N_1527,N_1352,N_1132);
xor U1528 (N_1528,N_1347,N_1065);
and U1529 (N_1529,N_1393,N_1354);
and U1530 (N_1530,N_1294,N_1279);
and U1531 (N_1531,N_1479,N_1181);
and U1532 (N_1532,N_1208,N_1236);
and U1533 (N_1533,N_1251,N_1289);
nand U1534 (N_1534,N_1009,N_1455);
or U1535 (N_1535,N_1253,N_1020);
or U1536 (N_1536,N_1356,N_1361);
nor U1537 (N_1537,N_1295,N_1468);
and U1538 (N_1538,N_1315,N_1384);
and U1539 (N_1539,N_1312,N_1235);
and U1540 (N_1540,N_1197,N_1319);
xor U1541 (N_1541,N_1185,N_1221);
or U1542 (N_1542,N_1438,N_1244);
nand U1543 (N_1543,N_1414,N_1489);
xnor U1544 (N_1544,N_1041,N_1337);
and U1545 (N_1545,N_1032,N_1407);
xnor U1546 (N_1546,N_1043,N_1058);
xor U1547 (N_1547,N_1093,N_1411);
or U1548 (N_1548,N_1001,N_1148);
xor U1549 (N_1549,N_1037,N_1496);
nand U1550 (N_1550,N_1080,N_1340);
or U1551 (N_1551,N_1423,N_1118);
and U1552 (N_1552,N_1188,N_1122);
and U1553 (N_1553,N_1406,N_1176);
nor U1554 (N_1554,N_1353,N_1408);
nand U1555 (N_1555,N_1369,N_1473);
xnor U1556 (N_1556,N_1292,N_1184);
nand U1557 (N_1557,N_1341,N_1410);
nand U1558 (N_1558,N_1426,N_1087);
nor U1559 (N_1559,N_1095,N_1444);
and U1560 (N_1560,N_1225,N_1030);
xor U1561 (N_1561,N_1383,N_1212);
or U1562 (N_1562,N_1374,N_1209);
xor U1563 (N_1563,N_1480,N_1282);
nor U1564 (N_1564,N_1026,N_1343);
nor U1565 (N_1565,N_1313,N_1447);
and U1566 (N_1566,N_1391,N_1089);
nand U1567 (N_1567,N_1137,N_1230);
nand U1568 (N_1568,N_1216,N_1227);
nor U1569 (N_1569,N_1346,N_1431);
nor U1570 (N_1570,N_1382,N_1263);
nor U1571 (N_1571,N_1469,N_1231);
or U1572 (N_1572,N_1483,N_1250);
or U1573 (N_1573,N_1323,N_1386);
or U1574 (N_1574,N_1098,N_1016);
nor U1575 (N_1575,N_1335,N_1155);
xor U1576 (N_1576,N_1121,N_1202);
and U1577 (N_1577,N_1034,N_1023);
and U1578 (N_1578,N_1085,N_1284);
nor U1579 (N_1579,N_1126,N_1245);
nor U1580 (N_1580,N_1127,N_1362);
or U1581 (N_1581,N_1207,N_1106);
xor U1582 (N_1582,N_1086,N_1099);
or U1583 (N_1583,N_1206,N_1421);
or U1584 (N_1584,N_1146,N_1075);
or U1585 (N_1585,N_1420,N_1425);
nand U1586 (N_1586,N_1301,N_1376);
nor U1587 (N_1587,N_1116,N_1049);
or U1588 (N_1588,N_1258,N_1320);
and U1589 (N_1589,N_1381,N_1419);
xnor U1590 (N_1590,N_1432,N_1152);
nand U1591 (N_1591,N_1033,N_1435);
xor U1592 (N_1592,N_1183,N_1130);
nand U1593 (N_1593,N_1403,N_1464);
nor U1594 (N_1594,N_1102,N_1220);
nand U1595 (N_1595,N_1266,N_1154);
nor U1596 (N_1596,N_1460,N_1186);
nand U1597 (N_1597,N_1304,N_1171);
or U1598 (N_1598,N_1167,N_1409);
or U1599 (N_1599,N_1133,N_1014);
xnor U1600 (N_1600,N_1194,N_1229);
and U1601 (N_1601,N_1311,N_1057);
xor U1602 (N_1602,N_1276,N_1103);
and U1603 (N_1603,N_1417,N_1046);
nor U1604 (N_1604,N_1124,N_1056);
nand U1605 (N_1605,N_1416,N_1373);
or U1606 (N_1606,N_1178,N_1213);
or U1607 (N_1607,N_1296,N_1144);
or U1608 (N_1608,N_1170,N_1071);
or U1609 (N_1609,N_1405,N_1441);
nand U1610 (N_1610,N_1070,N_1430);
xor U1611 (N_1611,N_1191,N_1240);
xor U1612 (N_1612,N_1298,N_1090);
nand U1613 (N_1613,N_1210,N_1010);
xor U1614 (N_1614,N_1198,N_1201);
and U1615 (N_1615,N_1217,N_1375);
or U1616 (N_1616,N_1072,N_1387);
and U1617 (N_1617,N_1241,N_1142);
and U1618 (N_1618,N_1285,N_1084);
or U1619 (N_1619,N_1108,N_1100);
nand U1620 (N_1620,N_1112,N_1274);
nor U1621 (N_1621,N_1002,N_1454);
xnor U1622 (N_1622,N_1446,N_1331);
xor U1623 (N_1623,N_1465,N_1060);
xor U1624 (N_1624,N_1445,N_1307);
or U1625 (N_1625,N_1200,N_1119);
nand U1626 (N_1626,N_1169,N_1302);
or U1627 (N_1627,N_1392,N_1064);
nor U1628 (N_1628,N_1135,N_1415);
xor U1629 (N_1629,N_1461,N_1088);
and U1630 (N_1630,N_1358,N_1139);
xor U1631 (N_1631,N_1242,N_1475);
or U1632 (N_1632,N_1272,N_1104);
nand U1633 (N_1633,N_1336,N_1401);
nor U1634 (N_1634,N_1243,N_1097);
nand U1635 (N_1635,N_1394,N_1436);
xnor U1636 (N_1636,N_1310,N_1173);
nand U1637 (N_1637,N_1481,N_1482);
xor U1638 (N_1638,N_1291,N_1003);
xor U1639 (N_1639,N_1031,N_1019);
nor U1640 (N_1640,N_1174,N_1264);
or U1641 (N_1641,N_1028,N_1136);
or U1642 (N_1642,N_1324,N_1478);
nor U1643 (N_1643,N_1380,N_1081);
nor U1644 (N_1644,N_1215,N_1390);
and U1645 (N_1645,N_1467,N_1288);
xor U1646 (N_1646,N_1252,N_1151);
xnor U1647 (N_1647,N_1271,N_1163);
or U1648 (N_1648,N_1308,N_1277);
and U1649 (N_1649,N_1027,N_1487);
or U1650 (N_1650,N_1063,N_1224);
and U1651 (N_1651,N_1110,N_1379);
or U1652 (N_1652,N_1300,N_1138);
xor U1653 (N_1653,N_1254,N_1349);
xnor U1654 (N_1654,N_1040,N_1328);
or U1655 (N_1655,N_1395,N_1494);
or U1656 (N_1656,N_1156,N_1491);
and U1657 (N_1657,N_1348,N_1018);
nand U1658 (N_1658,N_1364,N_1134);
nor U1659 (N_1659,N_1117,N_1143);
or U1660 (N_1660,N_1094,N_1287);
or U1661 (N_1661,N_1233,N_1205);
or U1662 (N_1662,N_1462,N_1477);
nand U1663 (N_1663,N_1377,N_1398);
nand U1664 (N_1664,N_1029,N_1223);
nand U1665 (N_1665,N_1286,N_1195);
and U1666 (N_1666,N_1490,N_1499);
nor U1667 (N_1667,N_1422,N_1062);
xor U1668 (N_1668,N_1015,N_1237);
or U1669 (N_1669,N_1055,N_1452);
nand U1670 (N_1670,N_1333,N_1260);
and U1671 (N_1671,N_1193,N_1321);
nand U1672 (N_1672,N_1283,N_1189);
or U1673 (N_1673,N_1351,N_1342);
nor U1674 (N_1674,N_1325,N_1168);
xor U1675 (N_1675,N_1273,N_1318);
nand U1676 (N_1676,N_1306,N_1449);
or U1677 (N_1677,N_1149,N_1367);
and U1678 (N_1678,N_1073,N_1024);
nand U1679 (N_1679,N_1153,N_1442);
nand U1680 (N_1680,N_1101,N_1008);
and U1681 (N_1681,N_1036,N_1109);
and U1682 (N_1682,N_1190,N_1261);
or U1683 (N_1683,N_1131,N_1397);
xor U1684 (N_1684,N_1115,N_1498);
nor U1685 (N_1685,N_1035,N_1365);
nand U1686 (N_1686,N_1443,N_1484);
nor U1687 (N_1687,N_1402,N_1187);
nor U1688 (N_1688,N_1021,N_1355);
xnor U1689 (N_1689,N_1158,N_1412);
xor U1690 (N_1690,N_1476,N_1453);
nand U1691 (N_1691,N_1068,N_1222);
nor U1692 (N_1692,N_1011,N_1140);
xor U1693 (N_1693,N_1275,N_1427);
or U1694 (N_1694,N_1161,N_1147);
and U1695 (N_1695,N_1434,N_1270);
and U1696 (N_1696,N_1472,N_1339);
nand U1697 (N_1697,N_1048,N_1199);
and U1698 (N_1698,N_1378,N_1322);
nor U1699 (N_1699,N_1162,N_1357);
nand U1700 (N_1700,N_1350,N_1107);
nand U1701 (N_1701,N_1067,N_1053);
nor U1702 (N_1702,N_1388,N_1025);
nor U1703 (N_1703,N_1334,N_1177);
nand U1704 (N_1704,N_1159,N_1281);
xor U1705 (N_1705,N_1069,N_1257);
nor U1706 (N_1706,N_1448,N_1440);
xnor U1707 (N_1707,N_1457,N_1165);
xor U1708 (N_1708,N_1247,N_1012);
nor U1709 (N_1709,N_1238,N_1228);
xor U1710 (N_1710,N_1203,N_1180);
or U1711 (N_1711,N_1196,N_1317);
and U1712 (N_1712,N_1413,N_1262);
nor U1713 (N_1713,N_1326,N_1051);
nand U1714 (N_1714,N_1486,N_1400);
or U1715 (N_1715,N_1141,N_1470);
and U1716 (N_1716,N_1497,N_1182);
or U1717 (N_1717,N_1017,N_1007);
and U1718 (N_1718,N_1061,N_1204);
or U1719 (N_1719,N_1459,N_1050);
nor U1720 (N_1720,N_1172,N_1248);
xnor U1721 (N_1721,N_1466,N_1371);
xnor U1722 (N_1722,N_1429,N_1327);
and U1723 (N_1723,N_1160,N_1366);
or U1724 (N_1724,N_1096,N_1111);
and U1725 (N_1725,N_1370,N_1006);
and U1726 (N_1726,N_1150,N_1218);
and U1727 (N_1727,N_1439,N_1458);
nor U1728 (N_1728,N_1052,N_1293);
xor U1729 (N_1729,N_1157,N_1129);
or U1730 (N_1730,N_1332,N_1039);
or U1731 (N_1731,N_1259,N_1290);
nand U1732 (N_1732,N_1249,N_1226);
and U1733 (N_1733,N_1396,N_1485);
nor U1734 (N_1734,N_1022,N_1192);
and U1735 (N_1735,N_1166,N_1437);
xor U1736 (N_1736,N_1329,N_1299);
nand U1737 (N_1737,N_1278,N_1113);
nor U1738 (N_1738,N_1372,N_1368);
nor U1739 (N_1739,N_1280,N_1246);
or U1740 (N_1740,N_1175,N_1211);
xnor U1741 (N_1741,N_1123,N_1066);
nand U1742 (N_1742,N_1359,N_1418);
nand U1743 (N_1743,N_1389,N_1399);
nor U1744 (N_1744,N_1269,N_1385);
and U1745 (N_1745,N_1239,N_1338);
xor U1746 (N_1746,N_1078,N_1038);
xor U1747 (N_1747,N_1042,N_1265);
nand U1748 (N_1748,N_1232,N_1493);
or U1749 (N_1749,N_1120,N_1077);
or U1750 (N_1750,N_1267,N_1434);
or U1751 (N_1751,N_1224,N_1015);
xor U1752 (N_1752,N_1138,N_1317);
and U1753 (N_1753,N_1386,N_1393);
and U1754 (N_1754,N_1038,N_1234);
nand U1755 (N_1755,N_1388,N_1425);
nand U1756 (N_1756,N_1452,N_1490);
or U1757 (N_1757,N_1493,N_1233);
xor U1758 (N_1758,N_1176,N_1205);
and U1759 (N_1759,N_1378,N_1014);
nand U1760 (N_1760,N_1191,N_1476);
and U1761 (N_1761,N_1053,N_1476);
nand U1762 (N_1762,N_1411,N_1226);
and U1763 (N_1763,N_1172,N_1302);
nand U1764 (N_1764,N_1028,N_1031);
or U1765 (N_1765,N_1286,N_1345);
nor U1766 (N_1766,N_1466,N_1218);
xor U1767 (N_1767,N_1135,N_1037);
or U1768 (N_1768,N_1274,N_1379);
or U1769 (N_1769,N_1324,N_1318);
xor U1770 (N_1770,N_1444,N_1013);
and U1771 (N_1771,N_1235,N_1097);
or U1772 (N_1772,N_1181,N_1151);
nor U1773 (N_1773,N_1296,N_1099);
or U1774 (N_1774,N_1186,N_1271);
nor U1775 (N_1775,N_1076,N_1328);
and U1776 (N_1776,N_1117,N_1472);
or U1777 (N_1777,N_1355,N_1454);
and U1778 (N_1778,N_1239,N_1371);
nor U1779 (N_1779,N_1012,N_1403);
or U1780 (N_1780,N_1363,N_1396);
xor U1781 (N_1781,N_1412,N_1313);
nor U1782 (N_1782,N_1054,N_1432);
or U1783 (N_1783,N_1386,N_1396);
or U1784 (N_1784,N_1440,N_1262);
xor U1785 (N_1785,N_1005,N_1230);
and U1786 (N_1786,N_1209,N_1367);
or U1787 (N_1787,N_1413,N_1043);
nor U1788 (N_1788,N_1080,N_1028);
or U1789 (N_1789,N_1029,N_1269);
nor U1790 (N_1790,N_1464,N_1215);
or U1791 (N_1791,N_1384,N_1034);
xor U1792 (N_1792,N_1498,N_1478);
xnor U1793 (N_1793,N_1333,N_1374);
nand U1794 (N_1794,N_1203,N_1194);
and U1795 (N_1795,N_1306,N_1346);
nand U1796 (N_1796,N_1486,N_1020);
and U1797 (N_1797,N_1371,N_1403);
xor U1798 (N_1798,N_1054,N_1310);
nand U1799 (N_1799,N_1306,N_1136);
and U1800 (N_1800,N_1029,N_1421);
nand U1801 (N_1801,N_1038,N_1016);
xor U1802 (N_1802,N_1393,N_1054);
nand U1803 (N_1803,N_1276,N_1346);
nand U1804 (N_1804,N_1310,N_1385);
xor U1805 (N_1805,N_1228,N_1065);
nand U1806 (N_1806,N_1107,N_1085);
or U1807 (N_1807,N_1265,N_1466);
and U1808 (N_1808,N_1280,N_1034);
and U1809 (N_1809,N_1024,N_1142);
and U1810 (N_1810,N_1434,N_1125);
nand U1811 (N_1811,N_1137,N_1390);
nand U1812 (N_1812,N_1323,N_1236);
and U1813 (N_1813,N_1434,N_1088);
xnor U1814 (N_1814,N_1113,N_1424);
nor U1815 (N_1815,N_1338,N_1291);
nand U1816 (N_1816,N_1045,N_1007);
and U1817 (N_1817,N_1122,N_1242);
xor U1818 (N_1818,N_1319,N_1083);
xnor U1819 (N_1819,N_1469,N_1052);
nor U1820 (N_1820,N_1436,N_1488);
or U1821 (N_1821,N_1374,N_1181);
nor U1822 (N_1822,N_1156,N_1465);
xor U1823 (N_1823,N_1193,N_1095);
nand U1824 (N_1824,N_1193,N_1145);
xor U1825 (N_1825,N_1006,N_1269);
nor U1826 (N_1826,N_1388,N_1010);
nand U1827 (N_1827,N_1359,N_1457);
and U1828 (N_1828,N_1462,N_1356);
or U1829 (N_1829,N_1123,N_1181);
xnor U1830 (N_1830,N_1168,N_1169);
or U1831 (N_1831,N_1482,N_1027);
or U1832 (N_1832,N_1442,N_1433);
or U1833 (N_1833,N_1189,N_1237);
nand U1834 (N_1834,N_1104,N_1178);
xor U1835 (N_1835,N_1191,N_1343);
and U1836 (N_1836,N_1257,N_1336);
xnor U1837 (N_1837,N_1308,N_1063);
nor U1838 (N_1838,N_1110,N_1093);
nor U1839 (N_1839,N_1185,N_1032);
and U1840 (N_1840,N_1311,N_1395);
xnor U1841 (N_1841,N_1205,N_1009);
nand U1842 (N_1842,N_1376,N_1449);
xor U1843 (N_1843,N_1409,N_1281);
nand U1844 (N_1844,N_1478,N_1408);
and U1845 (N_1845,N_1098,N_1022);
nor U1846 (N_1846,N_1167,N_1494);
and U1847 (N_1847,N_1405,N_1400);
or U1848 (N_1848,N_1492,N_1093);
xnor U1849 (N_1849,N_1438,N_1039);
nor U1850 (N_1850,N_1353,N_1210);
and U1851 (N_1851,N_1429,N_1095);
or U1852 (N_1852,N_1474,N_1168);
or U1853 (N_1853,N_1105,N_1122);
nor U1854 (N_1854,N_1073,N_1010);
and U1855 (N_1855,N_1011,N_1166);
xnor U1856 (N_1856,N_1081,N_1037);
or U1857 (N_1857,N_1448,N_1114);
xnor U1858 (N_1858,N_1409,N_1158);
and U1859 (N_1859,N_1361,N_1308);
nand U1860 (N_1860,N_1175,N_1300);
nor U1861 (N_1861,N_1223,N_1349);
nor U1862 (N_1862,N_1049,N_1122);
nand U1863 (N_1863,N_1427,N_1127);
and U1864 (N_1864,N_1076,N_1168);
nor U1865 (N_1865,N_1428,N_1075);
xnor U1866 (N_1866,N_1499,N_1273);
xnor U1867 (N_1867,N_1279,N_1004);
or U1868 (N_1868,N_1424,N_1131);
or U1869 (N_1869,N_1060,N_1439);
nand U1870 (N_1870,N_1395,N_1286);
nor U1871 (N_1871,N_1436,N_1216);
or U1872 (N_1872,N_1139,N_1122);
xnor U1873 (N_1873,N_1159,N_1042);
and U1874 (N_1874,N_1174,N_1324);
nand U1875 (N_1875,N_1190,N_1070);
xor U1876 (N_1876,N_1394,N_1466);
xor U1877 (N_1877,N_1011,N_1119);
xor U1878 (N_1878,N_1155,N_1212);
xor U1879 (N_1879,N_1137,N_1476);
xnor U1880 (N_1880,N_1176,N_1381);
nand U1881 (N_1881,N_1119,N_1378);
nand U1882 (N_1882,N_1184,N_1130);
or U1883 (N_1883,N_1117,N_1486);
and U1884 (N_1884,N_1325,N_1057);
nor U1885 (N_1885,N_1456,N_1243);
or U1886 (N_1886,N_1336,N_1435);
and U1887 (N_1887,N_1043,N_1322);
nand U1888 (N_1888,N_1109,N_1309);
xnor U1889 (N_1889,N_1406,N_1097);
nand U1890 (N_1890,N_1015,N_1218);
and U1891 (N_1891,N_1410,N_1106);
and U1892 (N_1892,N_1363,N_1310);
or U1893 (N_1893,N_1347,N_1098);
nor U1894 (N_1894,N_1443,N_1082);
nand U1895 (N_1895,N_1020,N_1003);
nand U1896 (N_1896,N_1406,N_1193);
or U1897 (N_1897,N_1458,N_1153);
nand U1898 (N_1898,N_1050,N_1231);
nand U1899 (N_1899,N_1307,N_1258);
nor U1900 (N_1900,N_1452,N_1006);
or U1901 (N_1901,N_1490,N_1193);
or U1902 (N_1902,N_1187,N_1275);
xor U1903 (N_1903,N_1467,N_1338);
and U1904 (N_1904,N_1366,N_1384);
and U1905 (N_1905,N_1488,N_1273);
nor U1906 (N_1906,N_1022,N_1319);
or U1907 (N_1907,N_1397,N_1386);
xor U1908 (N_1908,N_1232,N_1291);
nand U1909 (N_1909,N_1481,N_1040);
and U1910 (N_1910,N_1450,N_1123);
and U1911 (N_1911,N_1364,N_1023);
nor U1912 (N_1912,N_1451,N_1325);
or U1913 (N_1913,N_1425,N_1145);
or U1914 (N_1914,N_1234,N_1283);
nor U1915 (N_1915,N_1020,N_1403);
xor U1916 (N_1916,N_1477,N_1226);
nand U1917 (N_1917,N_1281,N_1400);
nor U1918 (N_1918,N_1423,N_1181);
and U1919 (N_1919,N_1123,N_1258);
nand U1920 (N_1920,N_1235,N_1172);
nor U1921 (N_1921,N_1016,N_1458);
nor U1922 (N_1922,N_1221,N_1321);
nand U1923 (N_1923,N_1418,N_1051);
xor U1924 (N_1924,N_1100,N_1359);
nand U1925 (N_1925,N_1161,N_1431);
and U1926 (N_1926,N_1266,N_1041);
nand U1927 (N_1927,N_1114,N_1224);
nand U1928 (N_1928,N_1148,N_1276);
xnor U1929 (N_1929,N_1053,N_1304);
nor U1930 (N_1930,N_1453,N_1007);
xor U1931 (N_1931,N_1174,N_1110);
nor U1932 (N_1932,N_1389,N_1404);
and U1933 (N_1933,N_1053,N_1062);
nand U1934 (N_1934,N_1114,N_1149);
nand U1935 (N_1935,N_1290,N_1449);
xor U1936 (N_1936,N_1172,N_1282);
nor U1937 (N_1937,N_1267,N_1096);
nor U1938 (N_1938,N_1212,N_1419);
nand U1939 (N_1939,N_1310,N_1190);
xnor U1940 (N_1940,N_1389,N_1075);
or U1941 (N_1941,N_1106,N_1000);
and U1942 (N_1942,N_1061,N_1340);
xor U1943 (N_1943,N_1306,N_1356);
and U1944 (N_1944,N_1183,N_1499);
xor U1945 (N_1945,N_1498,N_1143);
nor U1946 (N_1946,N_1445,N_1302);
nor U1947 (N_1947,N_1428,N_1247);
nor U1948 (N_1948,N_1290,N_1344);
or U1949 (N_1949,N_1367,N_1053);
xor U1950 (N_1950,N_1100,N_1279);
or U1951 (N_1951,N_1391,N_1034);
or U1952 (N_1952,N_1349,N_1377);
and U1953 (N_1953,N_1260,N_1330);
xor U1954 (N_1954,N_1347,N_1484);
nor U1955 (N_1955,N_1300,N_1133);
or U1956 (N_1956,N_1435,N_1050);
nand U1957 (N_1957,N_1235,N_1282);
xnor U1958 (N_1958,N_1499,N_1110);
or U1959 (N_1959,N_1319,N_1130);
nor U1960 (N_1960,N_1448,N_1198);
and U1961 (N_1961,N_1072,N_1197);
xnor U1962 (N_1962,N_1342,N_1461);
nand U1963 (N_1963,N_1249,N_1281);
or U1964 (N_1964,N_1189,N_1363);
nor U1965 (N_1965,N_1379,N_1485);
and U1966 (N_1966,N_1272,N_1461);
and U1967 (N_1967,N_1179,N_1398);
nor U1968 (N_1968,N_1338,N_1044);
nor U1969 (N_1969,N_1172,N_1347);
xor U1970 (N_1970,N_1160,N_1449);
and U1971 (N_1971,N_1112,N_1433);
and U1972 (N_1972,N_1321,N_1173);
xor U1973 (N_1973,N_1035,N_1243);
xor U1974 (N_1974,N_1221,N_1054);
and U1975 (N_1975,N_1029,N_1142);
nor U1976 (N_1976,N_1348,N_1176);
nand U1977 (N_1977,N_1186,N_1304);
xor U1978 (N_1978,N_1459,N_1000);
and U1979 (N_1979,N_1361,N_1425);
xor U1980 (N_1980,N_1079,N_1306);
nor U1981 (N_1981,N_1283,N_1421);
nand U1982 (N_1982,N_1120,N_1097);
nor U1983 (N_1983,N_1036,N_1151);
or U1984 (N_1984,N_1499,N_1407);
nand U1985 (N_1985,N_1024,N_1425);
xor U1986 (N_1986,N_1403,N_1184);
nand U1987 (N_1987,N_1063,N_1276);
nor U1988 (N_1988,N_1030,N_1145);
nand U1989 (N_1989,N_1065,N_1395);
or U1990 (N_1990,N_1417,N_1081);
nor U1991 (N_1991,N_1366,N_1483);
or U1992 (N_1992,N_1243,N_1352);
and U1993 (N_1993,N_1313,N_1125);
nand U1994 (N_1994,N_1113,N_1355);
nor U1995 (N_1995,N_1466,N_1458);
or U1996 (N_1996,N_1327,N_1370);
xnor U1997 (N_1997,N_1272,N_1076);
nand U1998 (N_1998,N_1178,N_1301);
nor U1999 (N_1999,N_1405,N_1157);
nand U2000 (N_2000,N_1899,N_1503);
nand U2001 (N_2001,N_1998,N_1594);
nor U2002 (N_2002,N_1919,N_1871);
or U2003 (N_2003,N_1885,N_1581);
nand U2004 (N_2004,N_1556,N_1873);
or U2005 (N_2005,N_1506,N_1927);
nand U2006 (N_2006,N_1531,N_1595);
nor U2007 (N_2007,N_1913,N_1995);
and U2008 (N_2008,N_1533,N_1662);
and U2009 (N_2009,N_1790,N_1601);
and U2010 (N_2010,N_1675,N_1818);
or U2011 (N_2011,N_1887,N_1981);
and U2012 (N_2012,N_1648,N_1750);
or U2013 (N_2013,N_1747,N_1759);
nand U2014 (N_2014,N_1572,N_1532);
and U2015 (N_2015,N_1612,N_1916);
nor U2016 (N_2016,N_1692,N_1744);
and U2017 (N_2017,N_1856,N_1574);
and U2018 (N_2018,N_1943,N_1700);
nand U2019 (N_2019,N_1688,N_1898);
or U2020 (N_2020,N_1569,N_1632);
xor U2021 (N_2021,N_1973,N_1693);
nand U2022 (N_2022,N_1705,N_1638);
or U2023 (N_2023,N_1925,N_1965);
or U2024 (N_2024,N_1729,N_1691);
and U2025 (N_2025,N_1970,N_1893);
xor U2026 (N_2026,N_1554,N_1855);
nor U2027 (N_2027,N_1507,N_1950);
and U2028 (N_2028,N_1961,N_1683);
or U2029 (N_2029,N_1817,N_1733);
or U2030 (N_2030,N_1980,N_1912);
and U2031 (N_2031,N_1639,N_1593);
xnor U2032 (N_2032,N_1796,N_1557);
nor U2033 (N_2033,N_1754,N_1960);
nor U2034 (N_2034,N_1968,N_1504);
or U2035 (N_2035,N_1578,N_1780);
nor U2036 (N_2036,N_1876,N_1978);
and U2037 (N_2037,N_1822,N_1728);
nor U2038 (N_2038,N_1529,N_1623);
xnor U2039 (N_2039,N_1618,N_1988);
nor U2040 (N_2040,N_1722,N_1999);
nand U2041 (N_2041,N_1828,N_1910);
xnor U2042 (N_2042,N_1591,N_1918);
or U2043 (N_2043,N_1837,N_1651);
or U2044 (N_2044,N_1841,N_1677);
nor U2045 (N_2045,N_1826,N_1636);
or U2046 (N_2046,N_1582,N_1795);
nand U2047 (N_2047,N_1809,N_1509);
and U2048 (N_2048,N_1838,N_1707);
or U2049 (N_2049,N_1971,N_1672);
nor U2050 (N_2050,N_1550,N_1902);
and U2051 (N_2051,N_1984,N_1619);
or U2052 (N_2052,N_1694,N_1966);
or U2053 (N_2053,N_1549,N_1717);
nor U2054 (N_2054,N_1541,N_1629);
nand U2055 (N_2055,N_1610,N_1931);
xnor U2056 (N_2056,N_1643,N_1954);
and U2057 (N_2057,N_1654,N_1952);
xor U2058 (N_2058,N_1777,N_1989);
nand U2059 (N_2059,N_1656,N_1868);
or U2060 (N_2060,N_1706,N_1637);
or U2061 (N_2061,N_1860,N_1908);
or U2062 (N_2062,N_1634,N_1975);
and U2063 (N_2063,N_1686,N_1781);
nand U2064 (N_2064,N_1830,N_1928);
xor U2065 (N_2065,N_1977,N_1606);
nand U2066 (N_2066,N_1527,N_1834);
nand U2067 (N_2067,N_1511,N_1586);
xor U2068 (N_2068,N_1821,N_1732);
nor U2069 (N_2069,N_1811,N_1864);
nor U2070 (N_2070,N_1682,N_1888);
xor U2071 (N_2071,N_1911,N_1583);
xor U2072 (N_2072,N_1624,N_1650);
xor U2073 (N_2073,N_1563,N_1842);
nor U2074 (N_2074,N_1752,N_1616);
nand U2075 (N_2075,N_1832,N_1720);
xnor U2076 (N_2076,N_1579,N_1799);
nand U2077 (N_2077,N_1521,N_1807);
xnor U2078 (N_2078,N_1690,N_1661);
or U2079 (N_2079,N_1857,N_1939);
xor U2080 (N_2080,N_1784,N_1835);
or U2081 (N_2081,N_1801,N_1515);
xnor U2082 (N_2082,N_1644,N_1671);
nor U2083 (N_2083,N_1696,N_1813);
xnor U2084 (N_2084,N_1520,N_1814);
xnor U2085 (N_2085,N_1502,N_1559);
xor U2086 (N_2086,N_1877,N_1763);
or U2087 (N_2087,N_1798,N_1646);
nand U2088 (N_2088,N_1501,N_1831);
nor U2089 (N_2089,N_1879,N_1680);
and U2090 (N_2090,N_1674,N_1957);
and U2091 (N_2091,N_1820,N_1847);
nor U2092 (N_2092,N_1839,N_1940);
nand U2093 (N_2093,N_1766,N_1884);
and U2094 (N_2094,N_1553,N_1551);
nand U2095 (N_2095,N_1866,N_1577);
nor U2096 (N_2096,N_1737,N_1769);
and U2097 (N_2097,N_1566,N_1915);
xnor U2098 (N_2098,N_1562,N_1921);
and U2099 (N_2099,N_1914,N_1567);
xnor U2100 (N_2100,N_1738,N_1851);
xnor U2101 (N_2101,N_1512,N_1552);
xor U2102 (N_2102,N_1513,N_1805);
nor U2103 (N_2103,N_1575,N_1542);
nor U2104 (N_2104,N_1904,N_1723);
or U2105 (N_2105,N_1518,N_1959);
nor U2106 (N_2106,N_1663,N_1901);
and U2107 (N_2107,N_1770,N_1976);
nand U2108 (N_2108,N_1776,N_1649);
and U2109 (N_2109,N_1749,N_1714);
or U2110 (N_2110,N_1843,N_1709);
and U2111 (N_2111,N_1526,N_1742);
and U2112 (N_2112,N_1875,N_1819);
or U2113 (N_2113,N_1882,N_1953);
nor U2114 (N_2114,N_1628,N_1755);
and U2115 (N_2115,N_1955,N_1734);
or U2116 (N_2116,N_1547,N_1545);
xor U2117 (N_2117,N_1779,N_1558);
xor U2118 (N_2118,N_1548,N_1889);
xnor U2119 (N_2119,N_1708,N_1844);
and U2120 (N_2120,N_1872,N_1712);
nor U2121 (N_2121,N_1703,N_1715);
xor U2122 (N_2122,N_1865,N_1560);
nand U2123 (N_2123,N_1956,N_1555);
nand U2124 (N_2124,N_1909,N_1540);
nand U2125 (N_2125,N_1568,N_1588);
nor U2126 (N_2126,N_1768,N_1640);
and U2127 (N_2127,N_1785,N_1510);
nand U2128 (N_2128,N_1571,N_1840);
nor U2129 (N_2129,N_1972,N_1938);
nor U2130 (N_2130,N_1967,N_1580);
nor U2131 (N_2131,N_1958,N_1861);
xor U2132 (N_2132,N_1815,N_1711);
nor U2133 (N_2133,N_1676,N_1621);
nor U2134 (N_2134,N_1516,N_1525);
nand U2135 (N_2135,N_1534,N_1762);
nand U2136 (N_2136,N_1543,N_1791);
nand U2137 (N_2137,N_1725,N_1930);
nor U2138 (N_2138,N_1753,N_1765);
nand U2139 (N_2139,N_1764,N_1922);
and U2140 (N_2140,N_1994,N_1642);
nor U2141 (N_2141,N_1743,N_1808);
and U2142 (N_2142,N_1736,N_1679);
nor U2143 (N_2143,N_1681,N_1891);
or U2144 (N_2144,N_1824,N_1685);
xor U2145 (N_2145,N_1848,N_1539);
xor U2146 (N_2146,N_1936,N_1829);
nor U2147 (N_2147,N_1782,N_1617);
or U2148 (N_2148,N_1528,N_1993);
nor U2149 (N_2149,N_1787,N_1933);
nand U2150 (N_2150,N_1945,N_1983);
and U2151 (N_2151,N_1850,N_1935);
nor U2152 (N_2152,N_1987,N_1695);
and U2153 (N_2153,N_1608,N_1620);
and U2154 (N_2154,N_1645,N_1853);
nor U2155 (N_2155,N_1730,N_1992);
nor U2156 (N_2156,N_1812,N_1990);
or U2157 (N_2157,N_1599,N_1716);
nand U2158 (N_2158,N_1757,N_1963);
nor U2159 (N_2159,N_1756,N_1721);
nor U2160 (N_2160,N_1854,N_1788);
or U2161 (N_2161,N_1783,N_1614);
nor U2162 (N_2162,N_1886,N_1974);
nand U2163 (N_2163,N_1699,N_1804);
or U2164 (N_2164,N_1923,N_1613);
nor U2165 (N_2165,N_1767,N_1584);
nand U2166 (N_2166,N_1985,N_1573);
nand U2167 (N_2167,N_1576,N_1626);
and U2168 (N_2168,N_1827,N_1803);
or U2169 (N_2169,N_1964,N_1689);
nand U2170 (N_2170,N_1878,N_1687);
nand U2171 (N_2171,N_1745,N_1704);
and U2172 (N_2172,N_1603,N_1622);
or U2173 (N_2173,N_1932,N_1863);
or U2174 (N_2174,N_1774,N_1845);
and U2175 (N_2175,N_1741,N_1655);
and U2176 (N_2176,N_1590,N_1997);
and U2177 (N_2177,N_1962,N_1657);
nor U2178 (N_2178,N_1806,N_1561);
and U2179 (N_2179,N_1773,N_1800);
nor U2180 (N_2180,N_1810,N_1701);
nor U2181 (N_2181,N_1710,N_1894);
nand U2182 (N_2182,N_1727,N_1949);
or U2183 (N_2183,N_1934,N_1607);
nor U2184 (N_2184,N_1598,N_1678);
nor U2185 (N_2185,N_1890,N_1836);
nor U2186 (N_2186,N_1937,N_1786);
xnor U2187 (N_2187,N_1740,N_1862);
or U2188 (N_2188,N_1917,N_1641);
xnor U2189 (N_2189,N_1615,N_1713);
nor U2190 (N_2190,N_1895,N_1630);
nand U2191 (N_2191,N_1587,N_1986);
nand U2192 (N_2192,N_1726,N_1697);
nor U2193 (N_2193,N_1524,N_1647);
nand U2194 (N_2194,N_1538,N_1523);
and U2195 (N_2195,N_1635,N_1668);
xnor U2196 (N_2196,N_1514,N_1565);
xnor U2197 (N_2197,N_1665,N_1905);
xor U2198 (N_2198,N_1920,N_1982);
xor U2199 (N_2199,N_1673,N_1944);
or U2200 (N_2200,N_1536,N_1991);
and U2201 (N_2201,N_1670,N_1941);
or U2202 (N_2202,N_1761,N_1631);
xor U2203 (N_2203,N_1772,N_1969);
xnor U2204 (N_2204,N_1698,N_1658);
or U2205 (N_2205,N_1896,N_1924);
or U2206 (N_2206,N_1846,N_1719);
nor U2207 (N_2207,N_1669,N_1883);
or U2208 (N_2208,N_1906,N_1942);
or U2209 (N_2209,N_1816,N_1602);
and U2210 (N_2210,N_1519,N_1794);
or U2211 (N_2211,N_1667,N_1739);
nand U2212 (N_2212,N_1625,N_1731);
or U2213 (N_2213,N_1535,N_1659);
nor U2214 (N_2214,N_1627,N_1979);
or U2215 (N_2215,N_1600,N_1793);
and U2216 (N_2216,N_1867,N_1858);
and U2217 (N_2217,N_1530,N_1564);
and U2218 (N_2218,N_1948,N_1609);
nor U2219 (N_2219,N_1881,N_1597);
nand U2220 (N_2220,N_1500,N_1505);
xor U2221 (N_2221,N_1748,N_1897);
and U2222 (N_2222,N_1570,N_1746);
xor U2223 (N_2223,N_1684,N_1522);
xnor U2224 (N_2224,N_1849,N_1605);
or U2225 (N_2225,N_1604,N_1508);
or U2226 (N_2226,N_1596,N_1892);
and U2227 (N_2227,N_1546,N_1585);
and U2228 (N_2228,N_1778,N_1859);
xnor U2229 (N_2229,N_1775,N_1633);
or U2230 (N_2230,N_1903,N_1537);
or U2231 (N_2231,N_1758,N_1825);
nor U2232 (N_2232,N_1900,N_1870);
or U2233 (N_2233,N_1592,N_1724);
nor U2234 (N_2234,N_1751,N_1660);
nand U2235 (N_2235,N_1517,N_1802);
or U2236 (N_2236,N_1926,N_1869);
or U2237 (N_2237,N_1544,N_1664);
nand U2238 (N_2238,N_1823,N_1880);
and U2239 (N_2239,N_1929,N_1702);
and U2240 (N_2240,N_1996,N_1946);
or U2241 (N_2241,N_1666,N_1833);
and U2242 (N_2242,N_1907,N_1874);
or U2243 (N_2243,N_1771,N_1611);
or U2244 (N_2244,N_1792,N_1653);
and U2245 (N_2245,N_1718,N_1797);
nor U2246 (N_2246,N_1852,N_1589);
and U2247 (N_2247,N_1789,N_1951);
xnor U2248 (N_2248,N_1947,N_1760);
nand U2249 (N_2249,N_1735,N_1652);
nor U2250 (N_2250,N_1938,N_1658);
and U2251 (N_2251,N_1707,N_1644);
and U2252 (N_2252,N_1836,N_1666);
nor U2253 (N_2253,N_1808,N_1637);
nand U2254 (N_2254,N_1697,N_1758);
or U2255 (N_2255,N_1990,N_1610);
nor U2256 (N_2256,N_1878,N_1949);
nor U2257 (N_2257,N_1919,N_1828);
nand U2258 (N_2258,N_1571,N_1594);
or U2259 (N_2259,N_1691,N_1736);
nor U2260 (N_2260,N_1508,N_1756);
nand U2261 (N_2261,N_1754,N_1595);
nor U2262 (N_2262,N_1857,N_1752);
xor U2263 (N_2263,N_1627,N_1637);
and U2264 (N_2264,N_1998,N_1893);
xnor U2265 (N_2265,N_1934,N_1564);
or U2266 (N_2266,N_1842,N_1649);
and U2267 (N_2267,N_1521,N_1685);
nor U2268 (N_2268,N_1549,N_1574);
xor U2269 (N_2269,N_1748,N_1715);
xnor U2270 (N_2270,N_1784,N_1810);
nand U2271 (N_2271,N_1754,N_1512);
nand U2272 (N_2272,N_1956,N_1668);
xnor U2273 (N_2273,N_1767,N_1615);
or U2274 (N_2274,N_1747,N_1695);
nand U2275 (N_2275,N_1508,N_1686);
nor U2276 (N_2276,N_1514,N_1987);
xnor U2277 (N_2277,N_1677,N_1768);
nand U2278 (N_2278,N_1707,N_1871);
xnor U2279 (N_2279,N_1914,N_1643);
xnor U2280 (N_2280,N_1776,N_1596);
nand U2281 (N_2281,N_1604,N_1673);
or U2282 (N_2282,N_1947,N_1607);
nor U2283 (N_2283,N_1559,N_1600);
nand U2284 (N_2284,N_1547,N_1881);
or U2285 (N_2285,N_1725,N_1632);
nand U2286 (N_2286,N_1930,N_1592);
nor U2287 (N_2287,N_1746,N_1924);
or U2288 (N_2288,N_1699,N_1637);
nand U2289 (N_2289,N_1695,N_1589);
nor U2290 (N_2290,N_1711,N_1579);
xor U2291 (N_2291,N_1779,N_1946);
nand U2292 (N_2292,N_1816,N_1860);
or U2293 (N_2293,N_1890,N_1818);
and U2294 (N_2294,N_1673,N_1981);
nand U2295 (N_2295,N_1778,N_1966);
nand U2296 (N_2296,N_1762,N_1690);
or U2297 (N_2297,N_1529,N_1539);
nand U2298 (N_2298,N_1991,N_1711);
nand U2299 (N_2299,N_1714,N_1876);
and U2300 (N_2300,N_1529,N_1584);
nand U2301 (N_2301,N_1634,N_1945);
nor U2302 (N_2302,N_1793,N_1544);
nor U2303 (N_2303,N_1995,N_1827);
nand U2304 (N_2304,N_1825,N_1570);
or U2305 (N_2305,N_1820,N_1692);
nand U2306 (N_2306,N_1849,N_1859);
nor U2307 (N_2307,N_1723,N_1611);
or U2308 (N_2308,N_1542,N_1615);
nand U2309 (N_2309,N_1968,N_1774);
xnor U2310 (N_2310,N_1921,N_1942);
xor U2311 (N_2311,N_1963,N_1720);
and U2312 (N_2312,N_1649,N_1550);
xnor U2313 (N_2313,N_1573,N_1797);
nand U2314 (N_2314,N_1896,N_1925);
or U2315 (N_2315,N_1939,N_1733);
or U2316 (N_2316,N_1720,N_1757);
nand U2317 (N_2317,N_1975,N_1779);
nand U2318 (N_2318,N_1617,N_1561);
xor U2319 (N_2319,N_1650,N_1710);
and U2320 (N_2320,N_1763,N_1696);
nor U2321 (N_2321,N_1929,N_1545);
and U2322 (N_2322,N_1727,N_1758);
nand U2323 (N_2323,N_1906,N_1712);
or U2324 (N_2324,N_1914,N_1512);
nor U2325 (N_2325,N_1738,N_1928);
nand U2326 (N_2326,N_1679,N_1830);
or U2327 (N_2327,N_1630,N_1644);
nor U2328 (N_2328,N_1724,N_1591);
and U2329 (N_2329,N_1760,N_1976);
nor U2330 (N_2330,N_1978,N_1816);
or U2331 (N_2331,N_1666,N_1882);
nor U2332 (N_2332,N_1618,N_1593);
nor U2333 (N_2333,N_1543,N_1666);
and U2334 (N_2334,N_1706,N_1578);
and U2335 (N_2335,N_1726,N_1585);
nor U2336 (N_2336,N_1861,N_1779);
and U2337 (N_2337,N_1851,N_1771);
nor U2338 (N_2338,N_1753,N_1839);
nand U2339 (N_2339,N_1962,N_1929);
and U2340 (N_2340,N_1546,N_1655);
and U2341 (N_2341,N_1753,N_1676);
nor U2342 (N_2342,N_1837,N_1988);
xor U2343 (N_2343,N_1664,N_1923);
and U2344 (N_2344,N_1638,N_1654);
and U2345 (N_2345,N_1875,N_1886);
and U2346 (N_2346,N_1707,N_1849);
nand U2347 (N_2347,N_1576,N_1967);
nand U2348 (N_2348,N_1771,N_1539);
nand U2349 (N_2349,N_1797,N_1598);
or U2350 (N_2350,N_1893,N_1811);
or U2351 (N_2351,N_1854,N_1745);
nand U2352 (N_2352,N_1869,N_1521);
and U2353 (N_2353,N_1653,N_1559);
or U2354 (N_2354,N_1917,N_1680);
or U2355 (N_2355,N_1694,N_1577);
nor U2356 (N_2356,N_1645,N_1818);
nor U2357 (N_2357,N_1872,N_1900);
or U2358 (N_2358,N_1774,N_1590);
and U2359 (N_2359,N_1770,N_1591);
xnor U2360 (N_2360,N_1880,N_1957);
or U2361 (N_2361,N_1536,N_1911);
or U2362 (N_2362,N_1574,N_1605);
or U2363 (N_2363,N_1831,N_1802);
nor U2364 (N_2364,N_1757,N_1671);
and U2365 (N_2365,N_1621,N_1875);
and U2366 (N_2366,N_1821,N_1659);
nand U2367 (N_2367,N_1692,N_1518);
and U2368 (N_2368,N_1854,N_1698);
nand U2369 (N_2369,N_1642,N_1803);
and U2370 (N_2370,N_1709,N_1589);
xor U2371 (N_2371,N_1905,N_1564);
nand U2372 (N_2372,N_1678,N_1661);
or U2373 (N_2373,N_1804,N_1999);
nand U2374 (N_2374,N_1516,N_1702);
nand U2375 (N_2375,N_1949,N_1954);
nand U2376 (N_2376,N_1744,N_1579);
nor U2377 (N_2377,N_1567,N_1660);
nand U2378 (N_2378,N_1782,N_1884);
nor U2379 (N_2379,N_1898,N_1781);
nand U2380 (N_2380,N_1888,N_1556);
or U2381 (N_2381,N_1727,N_1759);
xor U2382 (N_2382,N_1852,N_1979);
or U2383 (N_2383,N_1909,N_1617);
xnor U2384 (N_2384,N_1920,N_1899);
nand U2385 (N_2385,N_1607,N_1877);
nand U2386 (N_2386,N_1966,N_1796);
nand U2387 (N_2387,N_1779,N_1767);
xor U2388 (N_2388,N_1735,N_1942);
and U2389 (N_2389,N_1896,N_1947);
xor U2390 (N_2390,N_1751,N_1691);
and U2391 (N_2391,N_1897,N_1911);
nor U2392 (N_2392,N_1723,N_1733);
nor U2393 (N_2393,N_1690,N_1737);
nand U2394 (N_2394,N_1536,N_1531);
xor U2395 (N_2395,N_1909,N_1698);
and U2396 (N_2396,N_1685,N_1916);
or U2397 (N_2397,N_1740,N_1839);
xor U2398 (N_2398,N_1630,N_1914);
and U2399 (N_2399,N_1894,N_1718);
or U2400 (N_2400,N_1634,N_1749);
or U2401 (N_2401,N_1520,N_1799);
nand U2402 (N_2402,N_1826,N_1737);
or U2403 (N_2403,N_1974,N_1834);
and U2404 (N_2404,N_1774,N_1637);
nand U2405 (N_2405,N_1853,N_1784);
or U2406 (N_2406,N_1863,N_1803);
or U2407 (N_2407,N_1691,N_1715);
nand U2408 (N_2408,N_1866,N_1776);
and U2409 (N_2409,N_1783,N_1786);
xor U2410 (N_2410,N_1662,N_1973);
and U2411 (N_2411,N_1781,N_1561);
or U2412 (N_2412,N_1996,N_1966);
or U2413 (N_2413,N_1873,N_1870);
nand U2414 (N_2414,N_1816,N_1583);
nor U2415 (N_2415,N_1882,N_1888);
xor U2416 (N_2416,N_1820,N_1727);
xnor U2417 (N_2417,N_1674,N_1902);
xnor U2418 (N_2418,N_1641,N_1926);
or U2419 (N_2419,N_1501,N_1944);
and U2420 (N_2420,N_1882,N_1821);
nor U2421 (N_2421,N_1979,N_1570);
nand U2422 (N_2422,N_1901,N_1844);
or U2423 (N_2423,N_1736,N_1733);
nor U2424 (N_2424,N_1769,N_1603);
or U2425 (N_2425,N_1894,N_1748);
or U2426 (N_2426,N_1980,N_1901);
and U2427 (N_2427,N_1798,N_1952);
nand U2428 (N_2428,N_1685,N_1939);
and U2429 (N_2429,N_1729,N_1815);
nor U2430 (N_2430,N_1986,N_1755);
nor U2431 (N_2431,N_1876,N_1626);
nand U2432 (N_2432,N_1572,N_1746);
nor U2433 (N_2433,N_1614,N_1800);
or U2434 (N_2434,N_1588,N_1748);
xor U2435 (N_2435,N_1808,N_1759);
nand U2436 (N_2436,N_1816,N_1565);
or U2437 (N_2437,N_1807,N_1551);
or U2438 (N_2438,N_1577,N_1996);
nor U2439 (N_2439,N_1892,N_1812);
and U2440 (N_2440,N_1997,N_1521);
and U2441 (N_2441,N_1758,N_1925);
or U2442 (N_2442,N_1737,N_1816);
nand U2443 (N_2443,N_1730,N_1579);
and U2444 (N_2444,N_1945,N_1812);
nor U2445 (N_2445,N_1954,N_1907);
nand U2446 (N_2446,N_1721,N_1916);
nand U2447 (N_2447,N_1710,N_1601);
or U2448 (N_2448,N_1865,N_1606);
and U2449 (N_2449,N_1768,N_1732);
nor U2450 (N_2450,N_1598,N_1706);
xor U2451 (N_2451,N_1957,N_1923);
xnor U2452 (N_2452,N_1663,N_1838);
and U2453 (N_2453,N_1716,N_1913);
nand U2454 (N_2454,N_1670,N_1726);
nor U2455 (N_2455,N_1806,N_1580);
and U2456 (N_2456,N_1606,N_1971);
xor U2457 (N_2457,N_1994,N_1862);
nor U2458 (N_2458,N_1809,N_1900);
nor U2459 (N_2459,N_1604,N_1851);
nand U2460 (N_2460,N_1771,N_1888);
xnor U2461 (N_2461,N_1661,N_1891);
and U2462 (N_2462,N_1679,N_1952);
or U2463 (N_2463,N_1613,N_1872);
nor U2464 (N_2464,N_1861,N_1836);
and U2465 (N_2465,N_1920,N_1705);
xor U2466 (N_2466,N_1890,N_1865);
or U2467 (N_2467,N_1646,N_1593);
nand U2468 (N_2468,N_1766,N_1576);
or U2469 (N_2469,N_1932,N_1777);
nor U2470 (N_2470,N_1876,N_1861);
and U2471 (N_2471,N_1960,N_1861);
or U2472 (N_2472,N_1738,N_1660);
or U2473 (N_2473,N_1622,N_1521);
xnor U2474 (N_2474,N_1721,N_1762);
nor U2475 (N_2475,N_1978,N_1524);
nand U2476 (N_2476,N_1545,N_1636);
nor U2477 (N_2477,N_1673,N_1974);
nor U2478 (N_2478,N_1547,N_1768);
xnor U2479 (N_2479,N_1999,N_1896);
and U2480 (N_2480,N_1698,N_1534);
nor U2481 (N_2481,N_1944,N_1863);
nor U2482 (N_2482,N_1932,N_1517);
xor U2483 (N_2483,N_1778,N_1712);
xnor U2484 (N_2484,N_1513,N_1607);
or U2485 (N_2485,N_1791,N_1517);
xor U2486 (N_2486,N_1880,N_1679);
xnor U2487 (N_2487,N_1657,N_1501);
xnor U2488 (N_2488,N_1687,N_1809);
or U2489 (N_2489,N_1718,N_1838);
nor U2490 (N_2490,N_1772,N_1684);
nor U2491 (N_2491,N_1926,N_1814);
or U2492 (N_2492,N_1516,N_1594);
xnor U2493 (N_2493,N_1512,N_1747);
nor U2494 (N_2494,N_1586,N_1835);
xnor U2495 (N_2495,N_1933,N_1778);
nor U2496 (N_2496,N_1756,N_1917);
and U2497 (N_2497,N_1692,N_1695);
nor U2498 (N_2498,N_1757,N_1825);
and U2499 (N_2499,N_1845,N_1603);
or U2500 (N_2500,N_2403,N_2026);
or U2501 (N_2501,N_2289,N_2390);
and U2502 (N_2502,N_2030,N_2050);
or U2503 (N_2503,N_2330,N_2135);
nand U2504 (N_2504,N_2016,N_2239);
xnor U2505 (N_2505,N_2283,N_2182);
nand U2506 (N_2506,N_2272,N_2144);
xnor U2507 (N_2507,N_2373,N_2037);
or U2508 (N_2508,N_2290,N_2313);
and U2509 (N_2509,N_2394,N_2271);
nor U2510 (N_2510,N_2268,N_2348);
nor U2511 (N_2511,N_2459,N_2183);
nor U2512 (N_2512,N_2365,N_2265);
and U2513 (N_2513,N_2380,N_2109);
or U2514 (N_2514,N_2375,N_2022);
xor U2515 (N_2515,N_2275,N_2127);
or U2516 (N_2516,N_2303,N_2049);
nor U2517 (N_2517,N_2349,N_2370);
nand U2518 (N_2518,N_2464,N_2364);
nand U2519 (N_2519,N_2029,N_2273);
nor U2520 (N_2520,N_2320,N_2072);
nor U2521 (N_2521,N_2294,N_2287);
or U2522 (N_2522,N_2211,N_2034);
or U2523 (N_2523,N_2124,N_2422);
or U2524 (N_2524,N_2443,N_2085);
nor U2525 (N_2525,N_2151,N_2008);
xor U2526 (N_2526,N_2028,N_2453);
or U2527 (N_2527,N_2233,N_2446);
or U2528 (N_2528,N_2070,N_2323);
or U2529 (N_2529,N_2048,N_2417);
nand U2530 (N_2530,N_2346,N_2131);
or U2531 (N_2531,N_2335,N_2165);
or U2532 (N_2532,N_2156,N_2209);
nor U2533 (N_2533,N_2033,N_2445);
or U2534 (N_2534,N_2126,N_2471);
and U2535 (N_2535,N_2399,N_2001);
nor U2536 (N_2536,N_2059,N_2351);
and U2537 (N_2537,N_2477,N_2478);
nor U2538 (N_2538,N_2042,N_2189);
and U2539 (N_2539,N_2243,N_2087);
xor U2540 (N_2540,N_2485,N_2014);
nand U2541 (N_2541,N_2021,N_2123);
or U2542 (N_2542,N_2047,N_2291);
nand U2543 (N_2543,N_2460,N_2089);
or U2544 (N_2544,N_2244,N_2054);
nand U2545 (N_2545,N_2095,N_2164);
and U2546 (N_2546,N_2121,N_2322);
and U2547 (N_2547,N_2492,N_2230);
or U2548 (N_2548,N_2263,N_2497);
and U2549 (N_2549,N_2377,N_2279);
nor U2550 (N_2550,N_2111,N_2331);
xor U2551 (N_2551,N_2483,N_2077);
nand U2552 (N_2552,N_2411,N_2012);
and U2553 (N_2553,N_2005,N_2473);
nand U2554 (N_2554,N_2101,N_2440);
nor U2555 (N_2555,N_2385,N_2193);
nor U2556 (N_2556,N_2476,N_2451);
xnor U2557 (N_2557,N_2134,N_2307);
nand U2558 (N_2558,N_2137,N_2342);
or U2559 (N_2559,N_2425,N_2309);
or U2560 (N_2560,N_2073,N_2337);
and U2561 (N_2561,N_2391,N_2115);
or U2562 (N_2562,N_2332,N_2196);
nor U2563 (N_2563,N_2241,N_2299);
nand U2564 (N_2564,N_2490,N_2097);
nand U2565 (N_2565,N_2400,N_2000);
and U2566 (N_2566,N_2174,N_2438);
nor U2567 (N_2567,N_2247,N_2019);
xor U2568 (N_2568,N_2347,N_2061);
or U2569 (N_2569,N_2458,N_2282);
and U2570 (N_2570,N_2249,N_2103);
or U2571 (N_2571,N_2105,N_2318);
and U2572 (N_2572,N_2338,N_2494);
nor U2573 (N_2573,N_2013,N_2444);
and U2574 (N_2574,N_2392,N_2217);
nor U2575 (N_2575,N_2402,N_2065);
nand U2576 (N_2576,N_2213,N_2172);
xor U2577 (N_2577,N_2128,N_2468);
nand U2578 (N_2578,N_2122,N_2024);
nand U2579 (N_2579,N_2187,N_2130);
and U2580 (N_2580,N_2314,N_2071);
and U2581 (N_2581,N_2043,N_2110);
xor U2582 (N_2582,N_2099,N_2107);
nor U2583 (N_2583,N_2441,N_2310);
nor U2584 (N_2584,N_2256,N_2401);
or U2585 (N_2585,N_2051,N_2415);
xor U2586 (N_2586,N_2469,N_2218);
or U2587 (N_2587,N_2360,N_2255);
nand U2588 (N_2588,N_2363,N_2448);
nand U2589 (N_2589,N_2129,N_2094);
xnor U2590 (N_2590,N_2152,N_2383);
and U2591 (N_2591,N_2496,N_2421);
nand U2592 (N_2592,N_2173,N_2226);
nand U2593 (N_2593,N_2006,N_2430);
and U2594 (N_2594,N_2112,N_2202);
and U2595 (N_2595,N_2205,N_2133);
nand U2596 (N_2596,N_2092,N_2482);
or U2597 (N_2597,N_2428,N_2449);
or U2598 (N_2598,N_2486,N_2457);
nand U2599 (N_2599,N_2393,N_2186);
nor U2600 (N_2600,N_2082,N_2161);
nand U2601 (N_2601,N_2274,N_2308);
nor U2602 (N_2602,N_2336,N_2058);
and U2603 (N_2603,N_2035,N_2248);
and U2604 (N_2604,N_2168,N_2145);
and U2605 (N_2605,N_2491,N_2067);
nand U2606 (N_2606,N_2465,N_2228);
or U2607 (N_2607,N_2484,N_2276);
nor U2608 (N_2608,N_2177,N_2237);
nor U2609 (N_2609,N_2254,N_2378);
nand U2610 (N_2610,N_2044,N_2104);
nand U2611 (N_2611,N_2431,N_2192);
nand U2612 (N_2612,N_2084,N_2064);
nand U2613 (N_2613,N_2260,N_2052);
and U2614 (N_2614,N_2020,N_2297);
xor U2615 (N_2615,N_2231,N_2147);
nor U2616 (N_2616,N_2352,N_2113);
and U2617 (N_2617,N_2015,N_2433);
nor U2618 (N_2618,N_2120,N_2406);
nand U2619 (N_2619,N_2435,N_2143);
or U2620 (N_2620,N_2132,N_2463);
nor U2621 (N_2621,N_2389,N_2295);
or U2622 (N_2622,N_2055,N_2262);
nand U2623 (N_2623,N_2139,N_2079);
or U2624 (N_2624,N_2138,N_2327);
and U2625 (N_2625,N_2442,N_2093);
and U2626 (N_2626,N_2454,N_2286);
and U2627 (N_2627,N_2190,N_2447);
or U2628 (N_2628,N_2304,N_2366);
nor U2629 (N_2629,N_2040,N_2432);
xor U2630 (N_2630,N_2136,N_2158);
xnor U2631 (N_2631,N_2036,N_2096);
and U2632 (N_2632,N_2345,N_2329);
or U2633 (N_2633,N_2056,N_2009);
nor U2634 (N_2634,N_2155,N_2114);
nor U2635 (N_2635,N_2208,N_2199);
xor U2636 (N_2636,N_2369,N_2046);
nor U2637 (N_2637,N_2188,N_2269);
and U2638 (N_2638,N_2371,N_2429);
or U2639 (N_2639,N_2160,N_2277);
and U2640 (N_2640,N_2357,N_2367);
nor U2641 (N_2641,N_2225,N_2078);
xor U2642 (N_2642,N_2398,N_2060);
or U2643 (N_2643,N_2066,N_2281);
nor U2644 (N_2644,N_2359,N_2206);
and U2645 (N_2645,N_2409,N_2343);
nand U2646 (N_2646,N_2362,N_2220);
or U2647 (N_2647,N_2075,N_2414);
or U2648 (N_2648,N_2166,N_2475);
nand U2649 (N_2649,N_2372,N_2242);
and U2650 (N_2650,N_2162,N_2334);
nor U2651 (N_2651,N_2057,N_2002);
or U2652 (N_2652,N_2288,N_2227);
or U2653 (N_2653,N_2305,N_2424);
nor U2654 (N_2654,N_2253,N_2240);
xor U2655 (N_2655,N_2434,N_2023);
and U2656 (N_2656,N_2210,N_2266);
and U2657 (N_2657,N_2236,N_2149);
nand U2658 (N_2658,N_2474,N_2354);
and U2659 (N_2659,N_2419,N_2219);
or U2660 (N_2660,N_2148,N_2038);
nand U2661 (N_2661,N_2499,N_2039);
or U2662 (N_2662,N_2495,N_2204);
and U2663 (N_2663,N_2141,N_2410);
nor U2664 (N_2664,N_2376,N_2068);
or U2665 (N_2665,N_2339,N_2361);
or U2666 (N_2666,N_2452,N_2293);
xnor U2667 (N_2667,N_2498,N_2238);
and U2668 (N_2668,N_2150,N_2081);
nand U2669 (N_2669,N_2436,N_2063);
nand U2670 (N_2670,N_2181,N_2080);
nor U2671 (N_2671,N_2207,N_2197);
and U2672 (N_2672,N_2259,N_2176);
and U2673 (N_2673,N_2258,N_2203);
nor U2674 (N_2674,N_2179,N_2326);
and U2675 (N_2675,N_2032,N_2062);
nor U2676 (N_2676,N_2379,N_2387);
and U2677 (N_2677,N_2250,N_2386);
nor U2678 (N_2678,N_2450,N_2027);
nor U2679 (N_2679,N_2041,N_2280);
nand U2680 (N_2680,N_2312,N_2153);
nand U2681 (N_2681,N_2427,N_2224);
nand U2682 (N_2682,N_2221,N_2157);
xnor U2683 (N_2683,N_2201,N_2185);
xnor U2684 (N_2684,N_2355,N_2396);
nor U2685 (N_2685,N_2340,N_2108);
nand U2686 (N_2686,N_2083,N_2397);
xor U2687 (N_2687,N_2098,N_2480);
nor U2688 (N_2688,N_2461,N_2316);
xnor U2689 (N_2689,N_2317,N_2010);
and U2690 (N_2690,N_2292,N_2298);
nand U2691 (N_2691,N_2493,N_2353);
nand U2692 (N_2692,N_2423,N_2328);
or U2693 (N_2693,N_2102,N_2200);
and U2694 (N_2694,N_2116,N_2426);
nand U2695 (N_2695,N_2088,N_2350);
nor U2696 (N_2696,N_2489,N_2302);
or U2697 (N_2697,N_2358,N_2455);
nand U2698 (N_2698,N_2408,N_2344);
or U2699 (N_2699,N_2214,N_2167);
nor U2700 (N_2700,N_2488,N_2466);
nand U2701 (N_2701,N_2234,N_2481);
and U2702 (N_2702,N_2053,N_2017);
xnor U2703 (N_2703,N_2223,N_2222);
nand U2704 (N_2704,N_2229,N_2170);
or U2705 (N_2705,N_2456,N_2384);
xnor U2706 (N_2706,N_2086,N_2025);
or U2707 (N_2707,N_2119,N_2154);
and U2708 (N_2708,N_2175,N_2315);
xnor U2709 (N_2709,N_2163,N_2003);
xnor U2710 (N_2710,N_2074,N_2416);
nand U2711 (N_2711,N_2420,N_2178);
or U2712 (N_2712,N_2341,N_2246);
and U2713 (N_2713,N_2198,N_2270);
nor U2714 (N_2714,N_2252,N_2285);
xor U2715 (N_2715,N_2333,N_2300);
or U2716 (N_2716,N_2031,N_2467);
and U2717 (N_2717,N_2479,N_2382);
nand U2718 (N_2718,N_2267,N_2215);
and U2719 (N_2719,N_2251,N_2118);
or U2720 (N_2720,N_2090,N_2159);
and U2721 (N_2721,N_2325,N_2169);
and U2722 (N_2722,N_2437,N_2356);
and U2723 (N_2723,N_2418,N_2125);
xnor U2724 (N_2724,N_2045,N_2407);
xnor U2725 (N_2725,N_2412,N_2171);
xor U2726 (N_2726,N_2306,N_2368);
xnor U2727 (N_2727,N_2462,N_2194);
xor U2728 (N_2728,N_2076,N_2284);
nand U2729 (N_2729,N_2413,N_2232);
nor U2730 (N_2730,N_2069,N_2007);
or U2731 (N_2731,N_2235,N_2404);
nand U2732 (N_2732,N_2106,N_2487);
nand U2733 (N_2733,N_2278,N_2319);
xnor U2734 (N_2734,N_2004,N_2395);
and U2735 (N_2735,N_2142,N_2191);
xor U2736 (N_2736,N_2100,N_2180);
or U2737 (N_2737,N_2261,N_2195);
nand U2738 (N_2738,N_2324,N_2018);
nor U2739 (N_2739,N_2212,N_2301);
xnor U2740 (N_2740,N_2011,N_2470);
nand U2741 (N_2741,N_2321,N_2091);
nor U2742 (N_2742,N_2374,N_2216);
xor U2743 (N_2743,N_2146,N_2117);
xnor U2744 (N_2744,N_2184,N_2439);
nand U2745 (N_2745,N_2140,N_2311);
and U2746 (N_2746,N_2264,N_2257);
nand U2747 (N_2747,N_2472,N_2388);
and U2748 (N_2748,N_2296,N_2381);
and U2749 (N_2749,N_2405,N_2245);
xor U2750 (N_2750,N_2449,N_2397);
and U2751 (N_2751,N_2017,N_2187);
nand U2752 (N_2752,N_2147,N_2377);
or U2753 (N_2753,N_2348,N_2045);
nor U2754 (N_2754,N_2396,N_2227);
and U2755 (N_2755,N_2345,N_2225);
nor U2756 (N_2756,N_2376,N_2475);
nor U2757 (N_2757,N_2167,N_2463);
nand U2758 (N_2758,N_2009,N_2405);
or U2759 (N_2759,N_2360,N_2376);
and U2760 (N_2760,N_2037,N_2486);
and U2761 (N_2761,N_2117,N_2289);
and U2762 (N_2762,N_2297,N_2268);
nor U2763 (N_2763,N_2188,N_2205);
nor U2764 (N_2764,N_2340,N_2229);
xnor U2765 (N_2765,N_2439,N_2037);
or U2766 (N_2766,N_2051,N_2248);
nor U2767 (N_2767,N_2448,N_2460);
nand U2768 (N_2768,N_2164,N_2254);
nand U2769 (N_2769,N_2332,N_2494);
nor U2770 (N_2770,N_2312,N_2479);
nor U2771 (N_2771,N_2384,N_2268);
and U2772 (N_2772,N_2311,N_2223);
or U2773 (N_2773,N_2112,N_2176);
nand U2774 (N_2774,N_2325,N_2490);
or U2775 (N_2775,N_2481,N_2361);
and U2776 (N_2776,N_2077,N_2257);
xnor U2777 (N_2777,N_2135,N_2476);
or U2778 (N_2778,N_2342,N_2129);
or U2779 (N_2779,N_2120,N_2165);
nand U2780 (N_2780,N_2232,N_2336);
and U2781 (N_2781,N_2027,N_2307);
xor U2782 (N_2782,N_2446,N_2141);
and U2783 (N_2783,N_2205,N_2408);
nand U2784 (N_2784,N_2431,N_2156);
or U2785 (N_2785,N_2338,N_2359);
nand U2786 (N_2786,N_2413,N_2272);
or U2787 (N_2787,N_2360,N_2344);
xor U2788 (N_2788,N_2238,N_2435);
or U2789 (N_2789,N_2106,N_2459);
nand U2790 (N_2790,N_2029,N_2307);
or U2791 (N_2791,N_2231,N_2232);
xnor U2792 (N_2792,N_2153,N_2009);
nand U2793 (N_2793,N_2317,N_2002);
nor U2794 (N_2794,N_2374,N_2119);
xor U2795 (N_2795,N_2449,N_2184);
and U2796 (N_2796,N_2270,N_2265);
or U2797 (N_2797,N_2217,N_2131);
or U2798 (N_2798,N_2069,N_2209);
nand U2799 (N_2799,N_2133,N_2427);
and U2800 (N_2800,N_2226,N_2043);
xor U2801 (N_2801,N_2279,N_2162);
xnor U2802 (N_2802,N_2059,N_2148);
xor U2803 (N_2803,N_2085,N_2230);
or U2804 (N_2804,N_2370,N_2130);
nor U2805 (N_2805,N_2494,N_2149);
nand U2806 (N_2806,N_2270,N_2394);
and U2807 (N_2807,N_2310,N_2294);
or U2808 (N_2808,N_2206,N_2226);
nand U2809 (N_2809,N_2221,N_2019);
and U2810 (N_2810,N_2058,N_2420);
xor U2811 (N_2811,N_2131,N_2294);
nor U2812 (N_2812,N_2381,N_2230);
nor U2813 (N_2813,N_2229,N_2215);
xor U2814 (N_2814,N_2470,N_2111);
nand U2815 (N_2815,N_2072,N_2075);
and U2816 (N_2816,N_2138,N_2452);
or U2817 (N_2817,N_2104,N_2458);
and U2818 (N_2818,N_2048,N_2308);
xor U2819 (N_2819,N_2439,N_2328);
xnor U2820 (N_2820,N_2105,N_2275);
nand U2821 (N_2821,N_2466,N_2291);
nor U2822 (N_2822,N_2023,N_2456);
and U2823 (N_2823,N_2235,N_2169);
xor U2824 (N_2824,N_2092,N_2057);
and U2825 (N_2825,N_2471,N_2239);
or U2826 (N_2826,N_2194,N_2401);
or U2827 (N_2827,N_2294,N_2055);
xnor U2828 (N_2828,N_2258,N_2102);
or U2829 (N_2829,N_2485,N_2410);
xnor U2830 (N_2830,N_2118,N_2294);
xnor U2831 (N_2831,N_2067,N_2247);
nand U2832 (N_2832,N_2441,N_2115);
nor U2833 (N_2833,N_2125,N_2248);
xor U2834 (N_2834,N_2022,N_2497);
nand U2835 (N_2835,N_2268,N_2219);
nand U2836 (N_2836,N_2362,N_2131);
or U2837 (N_2837,N_2217,N_2118);
or U2838 (N_2838,N_2067,N_2007);
nor U2839 (N_2839,N_2114,N_2169);
or U2840 (N_2840,N_2313,N_2402);
nor U2841 (N_2841,N_2010,N_2083);
nor U2842 (N_2842,N_2454,N_2380);
xor U2843 (N_2843,N_2380,N_2062);
and U2844 (N_2844,N_2300,N_2329);
and U2845 (N_2845,N_2272,N_2376);
or U2846 (N_2846,N_2167,N_2145);
or U2847 (N_2847,N_2490,N_2464);
xor U2848 (N_2848,N_2041,N_2207);
xnor U2849 (N_2849,N_2353,N_2260);
nor U2850 (N_2850,N_2046,N_2428);
nor U2851 (N_2851,N_2089,N_2350);
or U2852 (N_2852,N_2417,N_2319);
nand U2853 (N_2853,N_2272,N_2421);
nand U2854 (N_2854,N_2068,N_2192);
or U2855 (N_2855,N_2374,N_2212);
or U2856 (N_2856,N_2478,N_2125);
xor U2857 (N_2857,N_2053,N_2125);
or U2858 (N_2858,N_2214,N_2244);
and U2859 (N_2859,N_2211,N_2329);
xnor U2860 (N_2860,N_2083,N_2246);
nand U2861 (N_2861,N_2097,N_2246);
xnor U2862 (N_2862,N_2394,N_2116);
nor U2863 (N_2863,N_2203,N_2349);
and U2864 (N_2864,N_2288,N_2205);
nor U2865 (N_2865,N_2316,N_2399);
or U2866 (N_2866,N_2455,N_2219);
and U2867 (N_2867,N_2115,N_2251);
or U2868 (N_2868,N_2304,N_2106);
and U2869 (N_2869,N_2019,N_2078);
nor U2870 (N_2870,N_2446,N_2084);
nor U2871 (N_2871,N_2455,N_2142);
nand U2872 (N_2872,N_2082,N_2022);
nor U2873 (N_2873,N_2239,N_2264);
and U2874 (N_2874,N_2199,N_2241);
nor U2875 (N_2875,N_2470,N_2320);
or U2876 (N_2876,N_2452,N_2367);
xnor U2877 (N_2877,N_2472,N_2463);
nand U2878 (N_2878,N_2400,N_2384);
xor U2879 (N_2879,N_2159,N_2200);
xor U2880 (N_2880,N_2376,N_2448);
nor U2881 (N_2881,N_2405,N_2067);
xor U2882 (N_2882,N_2481,N_2373);
or U2883 (N_2883,N_2422,N_2254);
xnor U2884 (N_2884,N_2367,N_2471);
nor U2885 (N_2885,N_2362,N_2252);
xor U2886 (N_2886,N_2208,N_2224);
nor U2887 (N_2887,N_2122,N_2137);
or U2888 (N_2888,N_2311,N_2262);
xnor U2889 (N_2889,N_2098,N_2221);
nor U2890 (N_2890,N_2122,N_2246);
nor U2891 (N_2891,N_2246,N_2166);
nand U2892 (N_2892,N_2402,N_2116);
xnor U2893 (N_2893,N_2128,N_2388);
nor U2894 (N_2894,N_2259,N_2271);
or U2895 (N_2895,N_2377,N_2491);
or U2896 (N_2896,N_2139,N_2000);
or U2897 (N_2897,N_2356,N_2064);
nand U2898 (N_2898,N_2427,N_2043);
and U2899 (N_2899,N_2101,N_2425);
and U2900 (N_2900,N_2267,N_2051);
nand U2901 (N_2901,N_2288,N_2216);
nand U2902 (N_2902,N_2440,N_2409);
nand U2903 (N_2903,N_2196,N_2303);
nor U2904 (N_2904,N_2384,N_2223);
nand U2905 (N_2905,N_2233,N_2485);
or U2906 (N_2906,N_2497,N_2286);
or U2907 (N_2907,N_2176,N_2178);
xnor U2908 (N_2908,N_2483,N_2143);
and U2909 (N_2909,N_2286,N_2492);
nor U2910 (N_2910,N_2466,N_2139);
nor U2911 (N_2911,N_2211,N_2007);
and U2912 (N_2912,N_2144,N_2421);
nor U2913 (N_2913,N_2172,N_2216);
nand U2914 (N_2914,N_2091,N_2259);
xor U2915 (N_2915,N_2493,N_2340);
or U2916 (N_2916,N_2274,N_2008);
xor U2917 (N_2917,N_2044,N_2198);
or U2918 (N_2918,N_2195,N_2332);
and U2919 (N_2919,N_2418,N_2174);
nand U2920 (N_2920,N_2396,N_2480);
nand U2921 (N_2921,N_2151,N_2276);
and U2922 (N_2922,N_2226,N_2248);
xnor U2923 (N_2923,N_2295,N_2317);
nand U2924 (N_2924,N_2207,N_2348);
xor U2925 (N_2925,N_2057,N_2165);
or U2926 (N_2926,N_2328,N_2289);
nor U2927 (N_2927,N_2374,N_2290);
and U2928 (N_2928,N_2384,N_2381);
nor U2929 (N_2929,N_2238,N_2254);
xor U2930 (N_2930,N_2356,N_2299);
xor U2931 (N_2931,N_2037,N_2008);
xnor U2932 (N_2932,N_2129,N_2198);
xnor U2933 (N_2933,N_2110,N_2361);
nor U2934 (N_2934,N_2135,N_2083);
or U2935 (N_2935,N_2019,N_2145);
or U2936 (N_2936,N_2193,N_2274);
nor U2937 (N_2937,N_2121,N_2404);
or U2938 (N_2938,N_2435,N_2254);
xor U2939 (N_2939,N_2130,N_2028);
and U2940 (N_2940,N_2494,N_2224);
xnor U2941 (N_2941,N_2122,N_2000);
xnor U2942 (N_2942,N_2132,N_2486);
nand U2943 (N_2943,N_2165,N_2287);
or U2944 (N_2944,N_2068,N_2182);
and U2945 (N_2945,N_2249,N_2030);
and U2946 (N_2946,N_2003,N_2186);
nand U2947 (N_2947,N_2232,N_2234);
xnor U2948 (N_2948,N_2235,N_2211);
nand U2949 (N_2949,N_2063,N_2465);
xor U2950 (N_2950,N_2011,N_2430);
nand U2951 (N_2951,N_2209,N_2473);
xor U2952 (N_2952,N_2354,N_2231);
and U2953 (N_2953,N_2241,N_2242);
nand U2954 (N_2954,N_2424,N_2062);
and U2955 (N_2955,N_2483,N_2039);
or U2956 (N_2956,N_2024,N_2199);
nor U2957 (N_2957,N_2457,N_2219);
nand U2958 (N_2958,N_2065,N_2010);
nor U2959 (N_2959,N_2282,N_2212);
nand U2960 (N_2960,N_2234,N_2011);
xor U2961 (N_2961,N_2139,N_2027);
or U2962 (N_2962,N_2366,N_2399);
xor U2963 (N_2963,N_2216,N_2268);
nand U2964 (N_2964,N_2176,N_2415);
xor U2965 (N_2965,N_2425,N_2238);
nand U2966 (N_2966,N_2485,N_2117);
nor U2967 (N_2967,N_2344,N_2035);
xnor U2968 (N_2968,N_2379,N_2057);
xnor U2969 (N_2969,N_2413,N_2416);
xor U2970 (N_2970,N_2395,N_2447);
xnor U2971 (N_2971,N_2206,N_2460);
xor U2972 (N_2972,N_2476,N_2218);
nand U2973 (N_2973,N_2054,N_2443);
and U2974 (N_2974,N_2358,N_2418);
nand U2975 (N_2975,N_2464,N_2469);
nor U2976 (N_2976,N_2136,N_2010);
and U2977 (N_2977,N_2495,N_2192);
nor U2978 (N_2978,N_2284,N_2171);
nand U2979 (N_2979,N_2309,N_2240);
or U2980 (N_2980,N_2227,N_2285);
nor U2981 (N_2981,N_2095,N_2436);
or U2982 (N_2982,N_2295,N_2002);
or U2983 (N_2983,N_2475,N_2148);
nor U2984 (N_2984,N_2040,N_2074);
or U2985 (N_2985,N_2496,N_2402);
nor U2986 (N_2986,N_2301,N_2310);
or U2987 (N_2987,N_2066,N_2057);
nor U2988 (N_2988,N_2209,N_2097);
nor U2989 (N_2989,N_2072,N_2468);
and U2990 (N_2990,N_2402,N_2309);
nor U2991 (N_2991,N_2200,N_2193);
and U2992 (N_2992,N_2445,N_2358);
nand U2993 (N_2993,N_2448,N_2303);
nor U2994 (N_2994,N_2306,N_2047);
and U2995 (N_2995,N_2143,N_2479);
or U2996 (N_2996,N_2075,N_2231);
xor U2997 (N_2997,N_2313,N_2277);
nor U2998 (N_2998,N_2047,N_2054);
or U2999 (N_2999,N_2334,N_2375);
nand UO_0 (O_0,N_2717,N_2737);
nand UO_1 (O_1,N_2688,N_2881);
or UO_2 (O_2,N_2646,N_2832);
nand UO_3 (O_3,N_2740,N_2641);
xor UO_4 (O_4,N_2566,N_2665);
nand UO_5 (O_5,N_2957,N_2711);
nor UO_6 (O_6,N_2515,N_2622);
or UO_7 (O_7,N_2917,N_2735);
and UO_8 (O_8,N_2989,N_2828);
and UO_9 (O_9,N_2897,N_2605);
xnor UO_10 (O_10,N_2676,N_2528);
nand UO_11 (O_11,N_2818,N_2943);
nand UO_12 (O_12,N_2777,N_2513);
or UO_13 (O_13,N_2656,N_2783);
or UO_14 (O_14,N_2601,N_2847);
xor UO_15 (O_15,N_2744,N_2823);
xor UO_16 (O_16,N_2529,N_2853);
xor UO_17 (O_17,N_2638,N_2830);
nor UO_18 (O_18,N_2617,N_2597);
and UO_19 (O_19,N_2563,N_2634);
or UO_20 (O_20,N_2501,N_2964);
nand UO_21 (O_21,N_2826,N_2752);
nor UO_22 (O_22,N_2922,N_2535);
nor UO_23 (O_23,N_2559,N_2785);
or UO_24 (O_24,N_2863,N_2558);
xnor UO_25 (O_25,N_2631,N_2836);
or UO_26 (O_26,N_2886,N_2739);
or UO_27 (O_27,N_2759,N_2707);
nand UO_28 (O_28,N_2817,N_2754);
nor UO_29 (O_29,N_2627,N_2802);
or UO_30 (O_30,N_2702,N_2969);
or UO_31 (O_31,N_2545,N_2531);
or UO_32 (O_32,N_2693,N_2990);
and UO_33 (O_33,N_2858,N_2787);
or UO_34 (O_34,N_2774,N_2846);
or UO_35 (O_35,N_2937,N_2584);
nor UO_36 (O_36,N_2507,N_2512);
nor UO_37 (O_37,N_2751,N_2961);
nor UO_38 (O_38,N_2644,N_2636);
nor UO_39 (O_39,N_2632,N_2748);
xnor UO_40 (O_40,N_2872,N_2508);
and UO_41 (O_41,N_2966,N_2546);
nand UO_42 (O_42,N_2903,N_2661);
nor UO_43 (O_43,N_2649,N_2583);
nand UO_44 (O_44,N_2762,N_2851);
and UO_45 (O_45,N_2600,N_2991);
xnor UO_46 (O_46,N_2557,N_2988);
and UO_47 (O_47,N_2521,N_2875);
xnor UO_48 (O_48,N_2891,N_2782);
nand UO_49 (O_49,N_2664,N_2596);
xor UO_50 (O_50,N_2797,N_2935);
and UO_51 (O_51,N_2995,N_2861);
xor UO_52 (O_52,N_2930,N_2526);
and UO_53 (O_53,N_2610,N_2723);
nor UO_54 (O_54,N_2540,N_2948);
or UO_55 (O_55,N_2510,N_2806);
or UO_56 (O_56,N_2997,N_2962);
and UO_57 (O_57,N_2727,N_2831);
nor UO_58 (O_58,N_2895,N_2800);
nor UO_59 (O_59,N_2811,N_2522);
nand UO_60 (O_60,N_2733,N_2586);
nand UO_61 (O_61,N_2950,N_2538);
or UO_62 (O_62,N_2657,N_2843);
nand UO_63 (O_63,N_2712,N_2708);
nand UO_64 (O_64,N_2992,N_2899);
nand UO_65 (O_65,N_2536,N_2652);
and UO_66 (O_66,N_2852,N_2793);
or UO_67 (O_67,N_2923,N_2690);
xnor UO_68 (O_68,N_2869,N_2682);
nand UO_69 (O_69,N_2790,N_2591);
or UO_70 (O_70,N_2564,N_2603);
or UO_71 (O_71,N_2896,N_2683);
and UO_72 (O_72,N_2942,N_2635);
nand UO_73 (O_73,N_2813,N_2946);
nand UO_74 (O_74,N_2810,N_2890);
nand UO_75 (O_75,N_2505,N_2833);
xor UO_76 (O_76,N_2854,N_2868);
nor UO_77 (O_77,N_2541,N_2678);
or UO_78 (O_78,N_2927,N_2855);
or UO_79 (O_79,N_2542,N_2721);
and UO_80 (O_80,N_2919,N_2822);
nor UO_81 (O_81,N_2898,N_2829);
xor UO_82 (O_82,N_2604,N_2933);
and UO_83 (O_83,N_2756,N_2953);
xor UO_84 (O_84,N_2550,N_2906);
xnor UO_85 (O_85,N_2567,N_2674);
xnor UO_86 (O_86,N_2889,N_2675);
and UO_87 (O_87,N_2620,N_2952);
xor UO_88 (O_88,N_2925,N_2523);
nand UO_89 (O_89,N_2956,N_2862);
or UO_90 (O_90,N_2812,N_2555);
and UO_91 (O_91,N_2849,N_2938);
nand UO_92 (O_92,N_2581,N_2981);
or UO_93 (O_93,N_2970,N_2517);
and UO_94 (O_94,N_2928,N_2659);
or UO_95 (O_95,N_2500,N_2742);
nor UO_96 (O_96,N_2568,N_2667);
nand UO_97 (O_97,N_2570,N_2893);
and UO_98 (O_98,N_2730,N_2619);
xnor UO_99 (O_99,N_2578,N_2613);
and UO_100 (O_100,N_2986,N_2609);
or UO_101 (O_101,N_2985,N_2954);
or UO_102 (O_102,N_2771,N_2960);
and UO_103 (O_103,N_2808,N_2718);
xnor UO_104 (O_104,N_2967,N_2788);
and UO_105 (O_105,N_2686,N_2687);
xor UO_106 (O_106,N_2900,N_2874);
or UO_107 (O_107,N_2894,N_2587);
xnor UO_108 (O_108,N_2731,N_2845);
xor UO_109 (O_109,N_2743,N_2647);
or UO_110 (O_110,N_2719,N_2639);
or UO_111 (O_111,N_2537,N_2792);
and UO_112 (O_112,N_2746,N_2525);
nand UO_113 (O_113,N_2625,N_2856);
or UO_114 (O_114,N_2629,N_2553);
nor UO_115 (O_115,N_2776,N_2554);
nand UO_116 (O_116,N_2716,N_2694);
nor UO_117 (O_117,N_2565,N_2901);
nor UO_118 (O_118,N_2544,N_2769);
and UO_119 (O_119,N_2663,N_2916);
and UO_120 (O_120,N_2685,N_2679);
nand UO_121 (O_121,N_2918,N_2527);
or UO_122 (O_122,N_2574,N_2931);
xor UO_123 (O_123,N_2978,N_2572);
and UO_124 (O_124,N_2670,N_2908);
nor UO_125 (O_125,N_2871,N_2884);
nor UO_126 (O_126,N_2623,N_2640);
nand UO_127 (O_127,N_2653,N_2791);
or UO_128 (O_128,N_2971,N_2532);
xor UO_129 (O_129,N_2681,N_2509);
and UO_130 (O_130,N_2616,N_2786);
and UO_131 (O_131,N_2765,N_2804);
or UO_132 (O_132,N_2691,N_2745);
nand UO_133 (O_133,N_2936,N_2904);
nand UO_134 (O_134,N_2562,N_2556);
nor UO_135 (O_135,N_2585,N_2924);
xor UO_136 (O_136,N_2710,N_2779);
nor UO_137 (O_137,N_2520,N_2741);
nand UO_138 (O_138,N_2980,N_2867);
or UO_139 (O_139,N_2949,N_2909);
and UO_140 (O_140,N_2534,N_2977);
xnor UO_141 (O_141,N_2883,N_2669);
nand UO_142 (O_142,N_2816,N_2848);
nand UO_143 (O_143,N_2673,N_2589);
or UO_144 (O_144,N_2524,N_2758);
or UO_145 (O_145,N_2579,N_2994);
xnor UO_146 (O_146,N_2934,N_2713);
nor UO_147 (O_147,N_2511,N_2614);
nor UO_148 (O_148,N_2955,N_2945);
or UO_149 (O_149,N_2866,N_2795);
and UO_150 (O_150,N_2618,N_2963);
nand UO_151 (O_151,N_2607,N_2888);
xor UO_152 (O_152,N_2926,N_2819);
or UO_153 (O_153,N_2764,N_2502);
and UO_154 (O_154,N_2680,N_2975);
nand UO_155 (O_155,N_2877,N_2753);
nor UO_156 (O_156,N_2914,N_2569);
xor UO_157 (O_157,N_2770,N_2666);
and UO_158 (O_158,N_2857,N_2767);
nor UO_159 (O_159,N_2865,N_2689);
and UO_160 (O_160,N_2518,N_2654);
or UO_161 (O_161,N_2630,N_2701);
xnor UO_162 (O_162,N_2593,N_2533);
nand UO_163 (O_163,N_2504,N_2803);
or UO_164 (O_164,N_2575,N_2728);
and UO_165 (O_165,N_2706,N_2850);
nand UO_166 (O_166,N_2703,N_2968);
nor UO_167 (O_167,N_2608,N_2696);
and UO_168 (O_168,N_2506,N_2996);
xnor UO_169 (O_169,N_2825,N_2621);
and UO_170 (O_170,N_2606,N_2648);
nand UO_171 (O_171,N_2870,N_2951);
and UO_172 (O_172,N_2514,N_2805);
and UO_173 (O_173,N_2913,N_2539);
nor UO_174 (O_174,N_2809,N_2842);
and UO_175 (O_175,N_2880,N_2543);
or UO_176 (O_176,N_2503,N_2976);
and UO_177 (O_177,N_2892,N_2768);
nand UO_178 (O_178,N_2612,N_2658);
or UO_179 (O_179,N_2965,N_2755);
and UO_180 (O_180,N_2775,N_2705);
nor UO_181 (O_181,N_2582,N_2726);
and UO_182 (O_182,N_2835,N_2983);
and UO_183 (O_183,N_2982,N_2530);
or UO_184 (O_184,N_2915,N_2902);
nor UO_185 (O_185,N_2637,N_2650);
nor UO_186 (O_186,N_2672,N_2761);
and UO_187 (O_187,N_2885,N_2662);
nor UO_188 (O_188,N_2939,N_2973);
and UO_189 (O_189,N_2827,N_2911);
nand UO_190 (O_190,N_2590,N_2715);
or UO_191 (O_191,N_2692,N_2729);
and UO_192 (O_192,N_2592,N_2594);
and UO_193 (O_193,N_2552,N_2910);
or UO_194 (O_194,N_2974,N_2738);
nor UO_195 (O_195,N_2611,N_2912);
xor UO_196 (O_196,N_2709,N_2781);
nand UO_197 (O_197,N_2814,N_2615);
nor UO_198 (O_198,N_2876,N_2516);
or UO_199 (O_199,N_2519,N_2628);
nor UO_200 (O_200,N_2920,N_2879);
xor UO_201 (O_201,N_2560,N_2887);
xor UO_202 (O_202,N_2633,N_2598);
xor UO_203 (O_203,N_2780,N_2671);
nand UO_204 (O_204,N_2704,N_2736);
nand UO_205 (O_205,N_2643,N_2750);
or UO_206 (O_206,N_2841,N_2757);
nor UO_207 (O_207,N_2747,N_2760);
nand UO_208 (O_208,N_2944,N_2749);
and UO_209 (O_209,N_2815,N_2838);
and UO_210 (O_210,N_2801,N_2837);
or UO_211 (O_211,N_2784,N_2548);
and UO_212 (O_212,N_2698,N_2722);
nor UO_213 (O_213,N_2668,N_2571);
nand UO_214 (O_214,N_2772,N_2547);
nor UO_215 (O_215,N_2860,N_2799);
xor UO_216 (O_216,N_2844,N_2882);
or UO_217 (O_217,N_2645,N_2700);
nor UO_218 (O_218,N_2905,N_2834);
nand UO_219 (O_219,N_2684,N_2873);
or UO_220 (O_220,N_2839,N_2807);
or UO_221 (O_221,N_2626,N_2660);
nand UO_222 (O_222,N_2766,N_2984);
nor UO_223 (O_223,N_2824,N_2714);
nor UO_224 (O_224,N_2624,N_2699);
and UO_225 (O_225,N_2789,N_2878);
nand UO_226 (O_226,N_2724,N_2958);
nor UO_227 (O_227,N_2773,N_2821);
or UO_228 (O_228,N_2642,N_2778);
nand UO_229 (O_229,N_2561,N_2820);
nand UO_230 (O_230,N_2677,N_2695);
xor UO_231 (O_231,N_2864,N_2921);
nor UO_232 (O_232,N_2573,N_2993);
nor UO_233 (O_233,N_2720,N_2987);
nor UO_234 (O_234,N_2655,N_2763);
nor UO_235 (O_235,N_2549,N_2551);
and UO_236 (O_236,N_2940,N_2580);
or UO_237 (O_237,N_2796,N_2979);
xnor UO_238 (O_238,N_2959,N_2932);
nand UO_239 (O_239,N_2725,N_2929);
and UO_240 (O_240,N_2599,N_2697);
or UO_241 (O_241,N_2732,N_2794);
nand UO_242 (O_242,N_2840,N_2588);
or UO_243 (O_243,N_2941,N_2798);
nor UO_244 (O_244,N_2999,N_2998);
and UO_245 (O_245,N_2947,N_2907);
xnor UO_246 (O_246,N_2576,N_2595);
and UO_247 (O_247,N_2651,N_2972);
xor UO_248 (O_248,N_2859,N_2577);
or UO_249 (O_249,N_2602,N_2734);
nand UO_250 (O_250,N_2961,N_2900);
xor UO_251 (O_251,N_2785,N_2881);
or UO_252 (O_252,N_2820,N_2532);
nand UO_253 (O_253,N_2867,N_2944);
nor UO_254 (O_254,N_2685,N_2510);
nand UO_255 (O_255,N_2572,N_2780);
xnor UO_256 (O_256,N_2631,N_2964);
xor UO_257 (O_257,N_2529,N_2952);
nand UO_258 (O_258,N_2807,N_2664);
xnor UO_259 (O_259,N_2525,N_2602);
nand UO_260 (O_260,N_2949,N_2600);
nor UO_261 (O_261,N_2729,N_2940);
and UO_262 (O_262,N_2976,N_2993);
nor UO_263 (O_263,N_2727,N_2607);
and UO_264 (O_264,N_2909,N_2535);
or UO_265 (O_265,N_2827,N_2720);
and UO_266 (O_266,N_2789,N_2920);
nor UO_267 (O_267,N_2943,N_2921);
and UO_268 (O_268,N_2748,N_2929);
or UO_269 (O_269,N_2625,N_2660);
xor UO_270 (O_270,N_2759,N_2650);
nor UO_271 (O_271,N_2705,N_2628);
nor UO_272 (O_272,N_2697,N_2732);
or UO_273 (O_273,N_2814,N_2748);
xnor UO_274 (O_274,N_2966,N_2918);
nor UO_275 (O_275,N_2653,N_2793);
and UO_276 (O_276,N_2680,N_2869);
xor UO_277 (O_277,N_2735,N_2567);
nand UO_278 (O_278,N_2588,N_2896);
nand UO_279 (O_279,N_2672,N_2833);
nor UO_280 (O_280,N_2778,N_2987);
or UO_281 (O_281,N_2504,N_2544);
xor UO_282 (O_282,N_2849,N_2977);
nor UO_283 (O_283,N_2884,N_2619);
xor UO_284 (O_284,N_2930,N_2756);
and UO_285 (O_285,N_2793,N_2914);
xor UO_286 (O_286,N_2953,N_2917);
xnor UO_287 (O_287,N_2860,N_2965);
xor UO_288 (O_288,N_2995,N_2651);
and UO_289 (O_289,N_2572,N_2522);
xnor UO_290 (O_290,N_2603,N_2619);
and UO_291 (O_291,N_2506,N_2647);
and UO_292 (O_292,N_2693,N_2837);
nor UO_293 (O_293,N_2836,N_2513);
or UO_294 (O_294,N_2743,N_2955);
nor UO_295 (O_295,N_2705,N_2850);
and UO_296 (O_296,N_2745,N_2741);
nand UO_297 (O_297,N_2571,N_2775);
xor UO_298 (O_298,N_2853,N_2594);
nand UO_299 (O_299,N_2506,N_2688);
and UO_300 (O_300,N_2851,N_2751);
and UO_301 (O_301,N_2913,N_2841);
nand UO_302 (O_302,N_2598,N_2848);
nand UO_303 (O_303,N_2897,N_2765);
nor UO_304 (O_304,N_2542,N_2973);
xor UO_305 (O_305,N_2514,N_2662);
or UO_306 (O_306,N_2536,N_2667);
xnor UO_307 (O_307,N_2860,N_2667);
or UO_308 (O_308,N_2879,N_2667);
nand UO_309 (O_309,N_2952,N_2839);
nor UO_310 (O_310,N_2636,N_2756);
xor UO_311 (O_311,N_2675,N_2847);
xor UO_312 (O_312,N_2973,N_2527);
or UO_313 (O_313,N_2942,N_2507);
and UO_314 (O_314,N_2789,N_2703);
xor UO_315 (O_315,N_2547,N_2672);
or UO_316 (O_316,N_2506,N_2944);
or UO_317 (O_317,N_2958,N_2947);
and UO_318 (O_318,N_2866,N_2701);
and UO_319 (O_319,N_2537,N_2699);
nand UO_320 (O_320,N_2577,N_2753);
nor UO_321 (O_321,N_2876,N_2787);
nand UO_322 (O_322,N_2567,N_2534);
nor UO_323 (O_323,N_2809,N_2733);
xnor UO_324 (O_324,N_2983,N_2825);
xor UO_325 (O_325,N_2749,N_2798);
nor UO_326 (O_326,N_2871,N_2595);
nand UO_327 (O_327,N_2903,N_2918);
xor UO_328 (O_328,N_2904,N_2568);
xor UO_329 (O_329,N_2794,N_2740);
and UO_330 (O_330,N_2569,N_2617);
xnor UO_331 (O_331,N_2965,N_2744);
xor UO_332 (O_332,N_2779,N_2882);
xnor UO_333 (O_333,N_2739,N_2570);
or UO_334 (O_334,N_2996,N_2857);
nor UO_335 (O_335,N_2898,N_2686);
nand UO_336 (O_336,N_2987,N_2892);
nand UO_337 (O_337,N_2565,N_2755);
nand UO_338 (O_338,N_2645,N_2874);
nand UO_339 (O_339,N_2754,N_2998);
nor UO_340 (O_340,N_2950,N_2741);
nor UO_341 (O_341,N_2881,N_2514);
and UO_342 (O_342,N_2523,N_2924);
and UO_343 (O_343,N_2948,N_2906);
or UO_344 (O_344,N_2789,N_2819);
nand UO_345 (O_345,N_2589,N_2786);
nand UO_346 (O_346,N_2573,N_2895);
xor UO_347 (O_347,N_2864,N_2715);
or UO_348 (O_348,N_2712,N_2517);
xor UO_349 (O_349,N_2630,N_2611);
or UO_350 (O_350,N_2861,N_2531);
nor UO_351 (O_351,N_2525,N_2652);
or UO_352 (O_352,N_2986,N_2977);
or UO_353 (O_353,N_2673,N_2732);
nor UO_354 (O_354,N_2571,N_2598);
nand UO_355 (O_355,N_2758,N_2882);
or UO_356 (O_356,N_2717,N_2695);
and UO_357 (O_357,N_2953,N_2713);
nor UO_358 (O_358,N_2668,N_2640);
xnor UO_359 (O_359,N_2883,N_2901);
xor UO_360 (O_360,N_2910,N_2525);
nor UO_361 (O_361,N_2789,N_2717);
nand UO_362 (O_362,N_2852,N_2900);
nand UO_363 (O_363,N_2592,N_2711);
nand UO_364 (O_364,N_2625,N_2713);
and UO_365 (O_365,N_2530,N_2538);
or UO_366 (O_366,N_2527,N_2906);
nand UO_367 (O_367,N_2964,N_2740);
nor UO_368 (O_368,N_2794,N_2514);
and UO_369 (O_369,N_2720,N_2994);
nand UO_370 (O_370,N_2717,N_2593);
xor UO_371 (O_371,N_2977,N_2677);
nor UO_372 (O_372,N_2694,N_2702);
and UO_373 (O_373,N_2612,N_2963);
nor UO_374 (O_374,N_2940,N_2675);
or UO_375 (O_375,N_2907,N_2677);
xnor UO_376 (O_376,N_2762,N_2591);
xnor UO_377 (O_377,N_2840,N_2841);
or UO_378 (O_378,N_2794,N_2738);
xnor UO_379 (O_379,N_2704,N_2752);
nand UO_380 (O_380,N_2538,N_2779);
or UO_381 (O_381,N_2521,N_2680);
nor UO_382 (O_382,N_2621,N_2635);
and UO_383 (O_383,N_2857,N_2919);
and UO_384 (O_384,N_2676,N_2713);
or UO_385 (O_385,N_2789,N_2891);
nand UO_386 (O_386,N_2894,N_2933);
nor UO_387 (O_387,N_2679,N_2922);
nor UO_388 (O_388,N_2859,N_2607);
and UO_389 (O_389,N_2925,N_2675);
and UO_390 (O_390,N_2579,N_2993);
nor UO_391 (O_391,N_2891,N_2931);
or UO_392 (O_392,N_2879,N_2932);
nor UO_393 (O_393,N_2822,N_2943);
xor UO_394 (O_394,N_2743,N_2782);
nand UO_395 (O_395,N_2634,N_2895);
or UO_396 (O_396,N_2928,N_2877);
nand UO_397 (O_397,N_2691,N_2774);
nand UO_398 (O_398,N_2604,N_2714);
xor UO_399 (O_399,N_2945,N_2962);
or UO_400 (O_400,N_2603,N_2726);
or UO_401 (O_401,N_2523,N_2885);
nand UO_402 (O_402,N_2650,N_2730);
nor UO_403 (O_403,N_2813,N_2918);
or UO_404 (O_404,N_2618,N_2874);
and UO_405 (O_405,N_2505,N_2609);
or UO_406 (O_406,N_2909,N_2646);
nand UO_407 (O_407,N_2845,N_2722);
xor UO_408 (O_408,N_2601,N_2727);
nand UO_409 (O_409,N_2872,N_2692);
or UO_410 (O_410,N_2713,N_2949);
xor UO_411 (O_411,N_2837,N_2833);
xnor UO_412 (O_412,N_2681,N_2697);
nor UO_413 (O_413,N_2846,N_2883);
xor UO_414 (O_414,N_2745,N_2936);
or UO_415 (O_415,N_2758,N_2666);
nand UO_416 (O_416,N_2718,N_2591);
or UO_417 (O_417,N_2590,N_2972);
and UO_418 (O_418,N_2912,N_2824);
nor UO_419 (O_419,N_2563,N_2835);
xor UO_420 (O_420,N_2881,N_2991);
nand UO_421 (O_421,N_2932,N_2600);
or UO_422 (O_422,N_2585,N_2915);
and UO_423 (O_423,N_2686,N_2670);
xor UO_424 (O_424,N_2511,N_2553);
nor UO_425 (O_425,N_2878,N_2507);
xor UO_426 (O_426,N_2828,N_2815);
nor UO_427 (O_427,N_2622,N_2829);
or UO_428 (O_428,N_2582,N_2986);
nor UO_429 (O_429,N_2703,N_2781);
or UO_430 (O_430,N_2778,N_2886);
nor UO_431 (O_431,N_2680,N_2755);
or UO_432 (O_432,N_2556,N_2730);
and UO_433 (O_433,N_2545,N_2912);
xnor UO_434 (O_434,N_2856,N_2590);
nor UO_435 (O_435,N_2755,N_2916);
nand UO_436 (O_436,N_2928,N_2931);
nand UO_437 (O_437,N_2796,N_2505);
and UO_438 (O_438,N_2592,N_2732);
and UO_439 (O_439,N_2601,N_2607);
nor UO_440 (O_440,N_2599,N_2765);
nand UO_441 (O_441,N_2864,N_2639);
xor UO_442 (O_442,N_2799,N_2930);
and UO_443 (O_443,N_2826,N_2554);
or UO_444 (O_444,N_2752,N_2766);
and UO_445 (O_445,N_2984,N_2770);
and UO_446 (O_446,N_2626,N_2899);
and UO_447 (O_447,N_2830,N_2972);
or UO_448 (O_448,N_2613,N_2900);
or UO_449 (O_449,N_2662,N_2552);
nor UO_450 (O_450,N_2889,N_2981);
xnor UO_451 (O_451,N_2622,N_2743);
xor UO_452 (O_452,N_2773,N_2769);
xnor UO_453 (O_453,N_2823,N_2869);
and UO_454 (O_454,N_2873,N_2894);
and UO_455 (O_455,N_2787,N_2770);
xor UO_456 (O_456,N_2863,N_2923);
xor UO_457 (O_457,N_2933,N_2783);
nor UO_458 (O_458,N_2547,N_2606);
or UO_459 (O_459,N_2902,N_2553);
xnor UO_460 (O_460,N_2714,N_2869);
and UO_461 (O_461,N_2696,N_2664);
xor UO_462 (O_462,N_2848,N_2717);
xnor UO_463 (O_463,N_2788,N_2972);
nor UO_464 (O_464,N_2620,N_2759);
nand UO_465 (O_465,N_2643,N_2557);
and UO_466 (O_466,N_2797,N_2689);
nand UO_467 (O_467,N_2580,N_2748);
nand UO_468 (O_468,N_2733,N_2768);
xor UO_469 (O_469,N_2873,N_2586);
or UO_470 (O_470,N_2880,N_2928);
nand UO_471 (O_471,N_2968,N_2706);
nor UO_472 (O_472,N_2632,N_2803);
and UO_473 (O_473,N_2889,N_2820);
nand UO_474 (O_474,N_2651,N_2617);
xnor UO_475 (O_475,N_2744,N_2993);
or UO_476 (O_476,N_2789,N_2868);
nor UO_477 (O_477,N_2826,N_2673);
or UO_478 (O_478,N_2834,N_2614);
or UO_479 (O_479,N_2973,N_2504);
xor UO_480 (O_480,N_2518,N_2752);
xnor UO_481 (O_481,N_2808,N_2702);
nand UO_482 (O_482,N_2943,N_2598);
or UO_483 (O_483,N_2512,N_2976);
or UO_484 (O_484,N_2670,N_2801);
and UO_485 (O_485,N_2817,N_2925);
nand UO_486 (O_486,N_2904,N_2785);
xnor UO_487 (O_487,N_2939,N_2753);
nand UO_488 (O_488,N_2861,N_2596);
or UO_489 (O_489,N_2537,N_2737);
and UO_490 (O_490,N_2800,N_2964);
or UO_491 (O_491,N_2794,N_2888);
xor UO_492 (O_492,N_2755,N_2563);
or UO_493 (O_493,N_2961,N_2608);
and UO_494 (O_494,N_2578,N_2921);
nand UO_495 (O_495,N_2553,N_2513);
or UO_496 (O_496,N_2754,N_2936);
nor UO_497 (O_497,N_2501,N_2644);
or UO_498 (O_498,N_2621,N_2734);
or UO_499 (O_499,N_2626,N_2591);
endmodule