module basic_1500_15000_2000_10_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_1048,In_57);
and U1 (N_1,In_423,In_719);
nor U2 (N_2,In_156,In_1331);
or U3 (N_3,In_916,In_304);
or U4 (N_4,In_662,In_1216);
xor U5 (N_5,In_1051,In_1499);
nand U6 (N_6,In_257,In_90);
nor U7 (N_7,In_788,In_914);
or U8 (N_8,In_1245,In_1463);
xor U9 (N_9,In_297,In_572);
and U10 (N_10,In_626,In_814);
and U11 (N_11,In_220,In_1104);
nor U12 (N_12,In_376,In_1050);
and U13 (N_13,In_1456,In_7);
nor U14 (N_14,In_1070,In_86);
or U15 (N_15,In_146,In_601);
nor U16 (N_16,In_1040,In_236);
nor U17 (N_17,In_1186,In_91);
nor U18 (N_18,In_591,In_1052);
nor U19 (N_19,In_1262,In_1253);
nor U20 (N_20,In_960,In_1238);
and U21 (N_21,In_312,In_1315);
and U22 (N_22,In_1351,In_647);
nor U23 (N_23,In_1251,In_231);
nor U24 (N_24,In_93,In_673);
and U25 (N_25,In_1483,In_393);
and U26 (N_26,In_1311,In_167);
nand U27 (N_27,In_1254,In_912);
or U28 (N_28,In_819,In_1343);
nor U29 (N_29,In_770,In_1289);
nor U30 (N_30,In_1386,In_1191);
or U31 (N_31,In_1210,In_1031);
or U32 (N_32,In_616,In_9);
or U33 (N_33,In_1105,In_964);
or U34 (N_34,In_735,In_1223);
nand U35 (N_35,In_507,In_858);
nand U36 (N_36,In_820,In_535);
and U37 (N_37,In_479,In_141);
nor U38 (N_38,In_642,In_1482);
and U39 (N_39,In_1076,In_1379);
xor U40 (N_40,In_557,In_965);
nor U41 (N_41,In_768,In_459);
nor U42 (N_42,In_802,In_751);
and U43 (N_43,In_1441,In_1298);
xor U44 (N_44,In_1147,In_119);
and U45 (N_45,In_358,In_1064);
or U46 (N_46,In_1329,In_546);
nor U47 (N_47,In_585,In_1222);
and U48 (N_48,In_1106,In_1145);
or U49 (N_49,In_1137,In_746);
and U50 (N_50,In_136,In_273);
and U51 (N_51,In_314,In_335);
and U52 (N_52,In_799,In_643);
xnor U53 (N_53,In_668,In_339);
nor U54 (N_54,In_1266,In_0);
and U55 (N_55,In_1382,In_1178);
and U56 (N_56,In_102,In_1131);
nand U57 (N_57,In_340,In_478);
nand U58 (N_58,In_827,In_1055);
xnor U59 (N_59,In_1065,In_1268);
and U60 (N_60,In_1190,In_785);
or U61 (N_61,In_945,In_1009);
or U62 (N_62,In_1108,In_696);
xor U63 (N_63,In_1330,In_260);
xnor U64 (N_64,In_1276,In_428);
and U65 (N_65,In_1209,In_515);
nand U66 (N_66,In_679,In_851);
nand U67 (N_67,In_503,In_75);
nand U68 (N_68,In_1470,In_889);
nand U69 (N_69,In_1007,In_1172);
nor U70 (N_70,In_112,In_812);
nor U71 (N_71,In_1487,In_382);
nor U72 (N_72,In_23,In_589);
and U73 (N_73,In_1024,In_961);
xor U74 (N_74,In_439,In_565);
nor U75 (N_75,In_1368,In_950);
and U76 (N_76,In_1449,In_494);
nand U77 (N_77,In_243,In_160);
and U78 (N_78,In_189,In_874);
or U79 (N_79,In_847,In_648);
nor U80 (N_80,In_975,In_1087);
nor U81 (N_81,In_850,In_372);
nor U82 (N_82,In_1498,In_794);
xor U83 (N_83,In_473,In_427);
or U84 (N_84,In_1119,In_1090);
xnor U85 (N_85,In_1317,In_158);
and U86 (N_86,In_1139,In_629);
xor U87 (N_87,In_1225,In_226);
and U88 (N_88,In_467,In_947);
or U89 (N_89,In_300,In_1165);
nor U90 (N_90,In_868,In_654);
nor U91 (N_91,In_952,In_837);
and U92 (N_92,In_398,In_1241);
nor U93 (N_93,In_957,In_993);
nor U94 (N_94,In_1468,In_869);
nor U95 (N_95,In_1492,In_415);
nand U96 (N_96,In_94,In_1120);
and U97 (N_97,In_468,In_717);
nor U98 (N_98,In_1391,In_1022);
and U99 (N_99,In_1229,In_342);
or U100 (N_100,In_53,In_476);
nor U101 (N_101,In_1306,In_1063);
xnor U102 (N_102,In_852,In_1479);
nor U103 (N_103,In_1219,In_140);
nand U104 (N_104,In_603,In_407);
xnor U105 (N_105,In_1142,In_653);
xnor U106 (N_106,In_1406,In_229);
nor U107 (N_107,In_153,In_1019);
nand U108 (N_108,In_491,In_677);
nor U109 (N_109,In_1061,In_622);
nand U110 (N_110,In_397,In_996);
or U111 (N_111,In_967,In_161);
xor U112 (N_112,In_5,In_1237);
nor U113 (N_113,In_1316,In_729);
nand U114 (N_114,In_646,In_1109);
nor U115 (N_115,In_330,In_1335);
xor U116 (N_116,In_442,In_1114);
or U117 (N_117,In_937,In_378);
xor U118 (N_118,In_337,In_587);
or U119 (N_119,In_1025,In_63);
xor U120 (N_120,In_877,In_324);
nor U121 (N_121,In_402,In_988);
and U122 (N_122,In_1123,In_1404);
xor U123 (N_123,In_1326,In_216);
or U124 (N_124,In_1297,In_309);
or U125 (N_125,In_660,In_1246);
xor U126 (N_126,In_1086,In_1193);
and U127 (N_127,In_292,In_1304);
or U128 (N_128,In_1028,In_1454);
or U129 (N_129,In_730,In_897);
nand U130 (N_130,In_495,In_1081);
nor U131 (N_131,In_1160,In_791);
or U132 (N_132,In_82,In_1320);
or U133 (N_133,In_892,In_1159);
nand U134 (N_134,In_365,In_544);
nor U135 (N_135,In_1486,In_1224);
nor U136 (N_136,In_835,In_1126);
or U137 (N_137,In_282,In_935);
xnor U138 (N_138,In_87,In_984);
and U139 (N_139,In_919,In_1097);
and U140 (N_140,In_526,In_240);
xor U141 (N_141,In_1099,In_702);
and U142 (N_142,In_1365,In_28);
xor U143 (N_143,In_39,In_180);
or U144 (N_144,In_361,In_1014);
or U145 (N_145,In_1157,In_833);
or U146 (N_146,In_804,In_1407);
xor U147 (N_147,In_285,In_1107);
nand U148 (N_148,In_215,In_55);
nor U149 (N_149,In_1079,In_334);
xnor U150 (N_150,In_1039,In_755);
nand U151 (N_151,In_554,In_264);
and U152 (N_152,In_560,In_21);
xnor U153 (N_153,In_253,In_1006);
nand U154 (N_154,In_512,In_172);
xor U155 (N_155,In_1041,In_567);
xnor U156 (N_156,In_1103,In_516);
xor U157 (N_157,In_661,In_981);
xnor U158 (N_158,In_883,In_840);
nor U159 (N_159,In_1258,In_1008);
nor U160 (N_160,In_1162,In_485);
xor U161 (N_161,In_807,In_448);
xor U162 (N_162,In_121,In_1452);
or U163 (N_163,In_199,In_724);
or U164 (N_164,In_898,In_1427);
nor U165 (N_165,In_70,In_1236);
xnor U166 (N_166,In_217,In_1445);
or U167 (N_167,In_1220,In_1464);
and U168 (N_168,In_839,In_1084);
and U169 (N_169,In_484,In_742);
nor U170 (N_170,In_813,In_893);
and U171 (N_171,In_523,In_737);
and U172 (N_172,In_1042,In_720);
and U173 (N_173,In_604,In_98);
nor U174 (N_174,In_612,In_1488);
or U175 (N_175,In_1455,In_1334);
nor U176 (N_176,In_1321,In_1332);
and U177 (N_177,In_88,In_227);
and U178 (N_178,In_1451,In_1425);
or U179 (N_179,In_1124,In_1066);
xnor U180 (N_180,In_345,In_1416);
and U181 (N_181,In_1462,In_771);
or U182 (N_182,In_1327,In_563);
xor U183 (N_183,In_671,In_1232);
nor U184 (N_184,In_821,In_1493);
xor U185 (N_185,In_1197,In_1323);
xnor U186 (N_186,In_1352,In_1442);
or U187 (N_187,In_235,In_997);
or U188 (N_188,In_1440,In_636);
xor U189 (N_189,In_1432,In_20);
xor U190 (N_190,In_287,In_162);
nor U191 (N_191,In_1111,In_913);
xnor U192 (N_192,In_1319,In_1211);
or U193 (N_193,In_774,In_188);
nand U194 (N_194,In_441,In_691);
nor U195 (N_195,In_205,In_645);
or U196 (N_196,In_1181,In_509);
or U197 (N_197,In_347,In_944);
and U198 (N_198,In_187,In_808);
nor U199 (N_199,In_741,In_1100);
and U200 (N_200,In_1378,In_296);
xor U201 (N_201,In_518,In_1077);
and U202 (N_202,In_886,In_1308);
xnor U203 (N_203,In_350,In_1281);
xnor U204 (N_204,In_795,In_811);
nor U205 (N_205,In_866,In_1001);
nand U206 (N_206,In_1200,In_191);
xnor U207 (N_207,In_941,In_1143);
xnor U208 (N_208,In_1011,In_530);
nand U209 (N_209,In_756,In_313);
or U210 (N_210,In_1047,In_793);
and U211 (N_211,In_1239,In_193);
or U212 (N_212,In_245,In_288);
and U213 (N_213,In_664,In_890);
nor U214 (N_214,In_711,In_1122);
and U215 (N_215,In_454,In_634);
nand U216 (N_216,In_558,In_790);
or U217 (N_217,In_1495,In_715);
nand U218 (N_218,In_1138,In_764);
or U219 (N_219,In_579,In_464);
nand U220 (N_220,In_832,In_66);
or U221 (N_221,In_129,In_765);
xnor U222 (N_222,In_888,In_954);
or U223 (N_223,In_1093,In_594);
and U224 (N_224,In_685,In_1096);
nor U225 (N_225,In_1476,In_1372);
nor U226 (N_226,In_614,In_34);
and U227 (N_227,In_991,In_627);
and U228 (N_228,In_480,In_1473);
xnor U229 (N_229,In_1152,In_1385);
and U230 (N_230,In_1265,In_413);
nor U231 (N_231,In_58,In_1337);
and U232 (N_232,In_578,In_766);
nor U233 (N_233,In_806,In_274);
nand U234 (N_234,In_628,In_761);
or U235 (N_235,In_435,In_905);
nor U236 (N_236,In_963,In_605);
nand U237 (N_237,In_1213,In_37);
or U238 (N_238,In_1448,In_708);
xnor U239 (N_239,In_1085,In_537);
nand U240 (N_240,In_79,In_1261);
xor U241 (N_241,In_303,In_564);
nand U242 (N_242,In_966,In_689);
or U243 (N_243,In_573,In_328);
nand U244 (N_244,In_584,In_598);
nand U245 (N_245,In_1046,In_989);
and U246 (N_246,In_922,In_316);
or U247 (N_247,In_475,In_1349);
and U248 (N_248,In_716,In_381);
nor U249 (N_249,In_182,In_453);
and U250 (N_250,In_203,In_657);
and U251 (N_251,In_1279,In_987);
or U252 (N_252,In_1023,In_780);
nand U253 (N_253,In_99,In_154);
nand U254 (N_254,In_105,In_817);
nand U255 (N_255,In_895,In_424);
nor U256 (N_256,In_778,In_500);
and U257 (N_257,In_1156,In_686);
xnor U258 (N_258,In_1285,In_1089);
nand U259 (N_259,In_867,In_49);
xor U260 (N_260,In_602,In_71);
or U261 (N_261,In_131,In_700);
and U262 (N_262,In_994,In_592);
nand U263 (N_263,In_504,In_450);
and U264 (N_264,In_1299,In_763);
xor U265 (N_265,In_1194,In_1328);
or U266 (N_266,In_531,In_1421);
nand U267 (N_267,In_1068,In_597);
nand U268 (N_268,In_1059,In_394);
xnor U269 (N_269,In_524,In_138);
nor U270 (N_270,In_803,In_1313);
or U271 (N_271,In_25,In_678);
and U272 (N_272,In_1417,In_1402);
or U273 (N_273,In_672,In_942);
nand U274 (N_274,In_1187,In_698);
xor U275 (N_275,In_797,In_45);
and U276 (N_276,In_1405,In_33);
nor U277 (N_277,In_444,In_218);
xor U278 (N_278,In_32,In_1158);
nand U279 (N_279,In_655,In_401);
nor U280 (N_280,In_792,In_81);
and U281 (N_281,In_1003,In_1430);
xor U282 (N_282,In_1133,In_165);
nor U283 (N_283,In_62,In_985);
nand U284 (N_284,In_1287,In_13);
or U285 (N_285,In_123,In_1243);
nor U286 (N_286,In_1384,In_48);
nor U287 (N_287,In_291,In_380);
and U288 (N_288,In_624,In_781);
nand U289 (N_289,In_122,In_465);
or U290 (N_290,In_590,In_968);
nor U291 (N_291,In_2,In_1370);
nor U292 (N_292,In_901,In_200);
xor U293 (N_293,In_667,In_437);
and U294 (N_294,In_574,In_980);
nand U295 (N_295,In_586,In_1004);
or U296 (N_296,In_1307,In_899);
or U297 (N_297,In_1339,In_175);
or U298 (N_298,In_1078,In_1350);
xor U299 (N_299,In_72,In_411);
xnor U300 (N_300,In_1242,In_1244);
and U301 (N_301,In_658,In_1249);
or U302 (N_302,In_387,In_1457);
xnor U303 (N_303,In_1188,In_214);
xnor U304 (N_304,In_1309,In_266);
or U305 (N_305,In_630,In_1175);
nand U306 (N_306,In_346,In_1098);
nand U307 (N_307,In_1393,In_593);
or U308 (N_308,In_61,In_1177);
nand U309 (N_309,In_1480,In_4);
or U310 (N_310,In_545,In_1214);
nor U311 (N_311,In_871,In_1082);
nor U312 (N_312,In_1037,In_341);
nand U313 (N_313,In_618,In_1458);
nor U314 (N_314,In_962,In_223);
nor U315 (N_315,In_894,In_1227);
nand U316 (N_316,In_1010,In_1288);
and U317 (N_317,In_1459,In_221);
and U318 (N_318,In_232,In_496);
or U319 (N_319,In_67,In_252);
nand U320 (N_320,In_1263,In_242);
nor U321 (N_321,In_1198,In_209);
nor U322 (N_322,In_1101,In_782);
nor U323 (N_323,In_492,In_404);
and U324 (N_324,In_306,In_463);
nor U325 (N_325,In_528,In_1259);
and U326 (N_326,In_1149,In_16);
or U327 (N_327,In_1020,In_390);
nand U328 (N_328,In_733,In_757);
nand U329 (N_329,In_280,In_457);
xnor U330 (N_330,In_436,In_955);
nand U331 (N_331,In_452,In_426);
xnor U332 (N_332,In_1389,In_576);
nand U333 (N_333,In_352,In_219);
xor U334 (N_334,In_1163,In_836);
xor U335 (N_335,In_329,In_1380);
nand U336 (N_336,In_1154,In_270);
or U337 (N_337,In_349,In_1234);
nand U338 (N_338,In_522,In_1208);
and U339 (N_339,In_619,In_860);
nor U340 (N_340,In_521,In_1044);
nand U341 (N_341,In_1282,In_1233);
xor U342 (N_342,In_174,In_106);
nand U343 (N_343,In_1409,In_1127);
nand U344 (N_344,In_1121,In_769);
and U345 (N_345,In_934,In_1112);
nor U346 (N_346,In_1102,In_145);
nand U347 (N_347,In_391,In_936);
or U348 (N_348,In_878,In_1400);
nor U349 (N_349,In_1490,In_115);
xnor U350 (N_350,In_451,In_320);
xor U351 (N_351,In_838,In_652);
nor U352 (N_352,In_255,In_1424);
nand U353 (N_353,In_1415,In_256);
or U354 (N_354,In_460,In_959);
nor U355 (N_355,In_1002,In_305);
or U356 (N_356,In_97,In_370);
and U357 (N_357,In_1255,In_732);
nor U358 (N_358,In_331,In_675);
nor U359 (N_359,In_853,In_826);
or U360 (N_360,In_1284,In_14);
nor U361 (N_361,In_1000,In_1141);
or U362 (N_362,In_447,In_1256);
and U363 (N_363,In_932,In_420);
nand U364 (N_364,In_114,In_117);
nor U365 (N_365,In_670,In_120);
nor U366 (N_366,In_754,In_1412);
nand U367 (N_367,In_699,In_1390);
and U368 (N_368,In_904,In_543);
nand U369 (N_369,In_1355,In_130);
and U370 (N_370,In_779,In_176);
xnor U371 (N_371,In_723,In_1305);
xnor U372 (N_372,In_1286,In_80);
and U373 (N_373,In_1273,In_855);
nor U374 (N_374,In_1179,In_879);
nor U375 (N_375,In_1168,In_24);
or U376 (N_376,In_953,In_1132);
nor U377 (N_377,In_322,In_1322);
and U378 (N_378,In_684,In_1377);
nor U379 (N_379,In_508,In_731);
xor U380 (N_380,In_635,In_929);
xor U381 (N_381,In_46,In_1074);
xnor U382 (N_382,In_1212,In_613);
or U383 (N_383,In_870,In_1477);
or U384 (N_384,In_179,In_164);
nor U385 (N_385,In_992,In_805);
and U386 (N_386,In_1032,In_1472);
nor U387 (N_387,In_1341,In_307);
nand U388 (N_388,In_38,In_17);
nor U389 (N_389,In_1036,In_360);
and U390 (N_390,In_293,In_862);
or U391 (N_391,In_422,In_1302);
nor U392 (N_392,In_621,In_30);
or U393 (N_393,In_1429,In_1240);
nand U394 (N_394,In_786,In_713);
nand U395 (N_395,In_816,In_308);
nand U396 (N_396,In_1228,In_326);
nand U397 (N_397,In_363,In_721);
and U398 (N_398,In_111,In_1460);
and U399 (N_399,In_1371,In_233);
and U400 (N_400,In_728,In_1344);
nor U401 (N_401,In_1401,In_656);
xor U402 (N_402,In_29,In_566);
nand U403 (N_403,In_828,In_84);
or U404 (N_404,In_810,In_611);
nand U405 (N_405,In_386,In_250);
or U406 (N_406,In_738,In_1413);
nand U407 (N_407,In_418,In_801);
nand U408 (N_408,In_623,In_1364);
nand U409 (N_409,In_789,In_1095);
nor U410 (N_410,In_607,In_758);
or U411 (N_411,In_863,In_178);
or U412 (N_412,In_1403,In_571);
nand U413 (N_413,In_343,In_752);
or U414 (N_414,In_267,In_10);
and U415 (N_415,In_1342,In_246);
and U416 (N_416,In_1312,In_784);
nor U417 (N_417,In_924,In_384);
or U418 (N_418,In_798,In_1248);
or U419 (N_419,In_1395,In_400);
nand U420 (N_420,In_744,In_95);
and U421 (N_421,In_555,In_44);
nor U422 (N_422,In_1235,In_1176);
nand U423 (N_423,In_1161,In_669);
nand U424 (N_424,In_829,In_318);
and U425 (N_425,In_157,In_1438);
nand U426 (N_426,In_562,In_481);
and U427 (N_427,In_1035,In_396);
and U428 (N_428,In_1129,In_1295);
or U429 (N_429,In_625,In_469);
xnor U430 (N_430,In_633,In_1428);
nor U431 (N_431,In_213,In_995);
xnor U432 (N_432,In_455,In_408);
nand U433 (N_433,In_323,In_375);
and U434 (N_434,In_1434,In_903);
nor U435 (N_435,In_1073,In_228);
or U436 (N_436,In_1414,In_1144);
nand U437 (N_437,In_948,In_1057);
or U438 (N_438,In_1481,In_529);
nand U439 (N_439,In_978,In_859);
nor U440 (N_440,In_186,In_1115);
nand U441 (N_441,In_1067,In_1450);
nand U442 (N_442,In_709,In_920);
or U443 (N_443,In_1475,In_1180);
and U444 (N_444,In_815,In_1189);
or U445 (N_445,In_973,In_854);
xor U446 (N_446,In_135,In_759);
or U447 (N_447,In_1366,In_1466);
or U448 (N_448,In_1336,In_550);
or U449 (N_449,In_527,In_1088);
xnor U450 (N_450,In_753,In_1484);
nand U451 (N_451,In_238,In_520);
and U452 (N_452,In_263,In_449);
and U453 (N_453,In_581,In_1361);
and U454 (N_454,In_353,In_665);
nand U455 (N_455,In_359,In_943);
nand U456 (N_456,In_1363,In_1345);
nor U457 (N_457,In_999,In_276);
and U458 (N_458,In_712,In_1267);
and U459 (N_459,In_1231,In_1423);
or U460 (N_460,In_1196,In_224);
xor U461 (N_461,In_928,In_173);
xnor U462 (N_462,In_762,In_727);
or U463 (N_463,In_971,In_1094);
and U464 (N_464,In_321,In_265);
and U465 (N_465,In_1062,In_1206);
nand U466 (N_466,In_1280,In_487);
xnor U467 (N_467,In_1376,In_680);
nand U468 (N_468,In_1069,In_775);
nor U469 (N_469,In_410,In_362);
nand U470 (N_470,In_338,In_101);
nor U471 (N_471,In_823,In_54);
nor U472 (N_472,In_534,In_1260);
nor U473 (N_473,In_979,In_659);
and U474 (N_474,In_818,In_1291);
xnor U475 (N_475,In_983,In_990);
xnor U476 (N_476,In_385,In_1174);
xor U477 (N_477,In_848,In_861);
and U478 (N_478,In_374,In_1408);
and U479 (N_479,In_891,In_525);
or U480 (N_480,In_974,In_703);
or U481 (N_481,In_1118,In_204);
or U482 (N_482,In_1347,In_906);
nor U483 (N_483,In_1348,In_290);
or U484 (N_484,In_1230,In_68);
xor U485 (N_485,In_262,In_1269);
or U486 (N_486,In_506,In_405);
nor U487 (N_487,In_644,In_750);
nand U488 (N_488,In_1381,In_1420);
nor U489 (N_489,In_725,In_1443);
and U490 (N_490,In_556,In_1060);
and U491 (N_491,In_251,In_921);
and U492 (N_492,In_1290,In_896);
nand U493 (N_493,In_748,In_1277);
xnor U494 (N_494,In_1387,In_726);
nor U495 (N_495,In_1354,In_225);
and U496 (N_496,In_809,In_139);
or U497 (N_497,In_110,In_159);
and U498 (N_498,In_170,In_864);
nor U499 (N_499,In_1013,In_632);
and U500 (N_500,In_1444,In_77);
and U501 (N_501,In_551,In_1043);
nor U502 (N_502,In_986,In_580);
and U503 (N_503,In_641,In_409);
nor U504 (N_504,In_369,In_278);
xnor U505 (N_505,In_517,In_379);
nand U506 (N_506,In_59,In_1447);
nand U507 (N_507,In_277,In_1226);
and U508 (N_508,In_295,In_104);
xor U509 (N_509,In_96,In_1092);
and U510 (N_510,In_946,In_332);
xnor U511 (N_511,In_900,In_1049);
nand U512 (N_512,In_933,In_514);
and U513 (N_513,In_583,In_1314);
xor U514 (N_514,In_1016,In_438);
and U515 (N_515,In_541,In_196);
xor U516 (N_516,In_1374,In_89);
xnor U517 (N_517,In_743,In_144);
and U518 (N_518,In_268,In_399);
xor U519 (N_519,In_505,In_1075);
nor U520 (N_520,In_902,In_760);
xor U521 (N_521,In_1026,In_461);
nor U522 (N_522,In_1439,In_976);
or U523 (N_523,In_132,In_687);
nand U524 (N_524,In_1310,In_969);
xnor U525 (N_525,In_283,In_796);
nand U526 (N_526,In_958,In_183);
or U527 (N_527,In_1091,In_650);
nor U528 (N_528,In_244,In_1296);
or U529 (N_529,In_317,In_800);
and U530 (N_530,In_190,In_315);
xnor U531 (N_531,In_234,In_458);
or U532 (N_532,In_849,In_207);
nand U533 (N_533,In_1205,In_1474);
nand U534 (N_534,In_876,In_78);
xor U535 (N_535,In_1030,In_406);
and U536 (N_536,In_1446,In_462);
or U537 (N_537,In_887,In_1017);
nand U538 (N_538,In_872,In_615);
and U539 (N_539,In_511,In_620);
or U540 (N_540,In_383,In_116);
xnor U541 (N_541,In_367,In_606);
nand U542 (N_542,In_1293,In_676);
nor U543 (N_543,In_777,In_1369);
or U544 (N_544,In_65,In_683);
nor U545 (N_545,In_1140,In_513);
or U546 (N_546,In_237,In_1155);
nand U547 (N_547,In_956,In_222);
xor U548 (N_548,In_134,In_666);
nand U549 (N_549,In_1171,In_42);
or U550 (N_550,In_553,In_1394);
or U551 (N_551,In_210,In_171);
xnor U552 (N_552,In_1362,In_843);
xor U553 (N_553,In_1058,In_1333);
nor U554 (N_554,In_1467,In_502);
nor U555 (N_555,In_249,In_610);
or U556 (N_556,In_181,In_1469);
or U557 (N_557,In_510,In_64);
or U558 (N_558,In_885,In_881);
nor U559 (N_559,In_289,In_198);
xnor U560 (N_560,In_1151,In_125);
or U561 (N_561,In_772,In_1436);
nor U562 (N_562,In_1183,In_575);
xnor U563 (N_563,In_206,In_831);
nor U564 (N_564,In_1325,In_1083);
and U565 (N_565,In_1426,In_127);
nor U566 (N_566,In_128,In_561);
nor U567 (N_567,In_1117,In_364);
or U568 (N_568,In_1125,In_416);
nor U569 (N_569,In_429,In_825);
and U570 (N_570,In_133,In_298);
nor U571 (N_571,In_472,In_76);
and U572 (N_572,In_1471,In_395);
or U573 (N_573,In_1461,In_970);
or U574 (N_574,In_1398,In_1038);
and U575 (N_575,In_1034,In_22);
and U576 (N_576,In_26,In_582);
and U577 (N_577,In_357,In_184);
xnor U578 (N_578,In_1278,In_705);
xnor U579 (N_579,In_498,In_163);
nand U580 (N_580,In_1410,In_907);
or U581 (N_581,In_1029,In_1437);
nor U582 (N_582,In_1113,In_663);
and U583 (N_583,In_1399,In_466);
and U584 (N_584,In_588,In_43);
xnor U585 (N_585,In_241,In_532);
or U586 (N_586,In_51,In_747);
and U587 (N_587,In_834,In_1359);
or U588 (N_588,In_830,In_690);
or U589 (N_589,In_301,In_1173);
or U590 (N_590,In_1489,In_739);
or U591 (N_591,In_841,In_927);
or U592 (N_592,In_445,In_1358);
nor U593 (N_593,In_166,In_417);
nor U594 (N_594,In_595,In_354);
nor U595 (N_595,In_373,In_208);
xnor U596 (N_596,In_325,In_882);
nor U597 (N_597,In_577,In_552);
nand U598 (N_598,In_1274,In_11);
and U599 (N_599,In_1164,In_599);
and U600 (N_600,In_177,In_740);
nor U601 (N_601,In_701,In_477);
xor U602 (N_602,In_880,In_923);
and U603 (N_603,In_272,In_842);
nand U604 (N_604,In_3,In_142);
or U605 (N_605,In_1465,In_540);
xor U606 (N_606,In_100,In_239);
xor U607 (N_607,In_1292,In_27);
or U608 (N_608,In_931,In_344);
xor U609 (N_609,In_403,In_682);
xor U610 (N_610,In_714,In_1146);
or U611 (N_611,In_490,In_143);
xor U612 (N_612,In_776,In_1202);
xnor U613 (N_613,In_147,In_1392);
xor U614 (N_614,In_1135,In_169);
nand U615 (N_615,In_824,In_275);
or U616 (N_616,In_471,In_1080);
and U617 (N_617,In_1045,In_431);
nand U618 (N_618,In_8,In_1411);
nand U619 (N_619,In_1116,In_1453);
nand U620 (N_620,In_486,In_938);
or U621 (N_621,In_1419,In_559);
or U622 (N_622,In_609,In_1167);
and U623 (N_623,In_1203,In_548);
and U624 (N_624,In_1217,In_40);
and U625 (N_625,In_536,In_1272);
and U626 (N_626,In_773,In_197);
xor U627 (N_627,In_425,In_474);
and U628 (N_628,In_875,In_1271);
xor U629 (N_629,In_918,In_631);
nand U630 (N_630,In_150,In_1134);
or U631 (N_631,In_1166,In_547);
nand U632 (N_632,In_734,In_706);
and U633 (N_633,In_1264,In_499);
nand U634 (N_634,In_1340,In_56);
or U635 (N_635,In_185,In_638);
and U636 (N_636,In_168,In_355);
xor U637 (N_637,In_1491,In_1207);
nor U638 (N_638,In_412,In_19);
nand U639 (N_639,In_1218,In_1054);
xor U640 (N_640,In_940,In_600);
nand U641 (N_641,In_542,In_749);
nand U642 (N_642,In_389,In_908);
or U643 (N_643,In_36,In_430);
nor U644 (N_644,In_1012,In_421);
and U645 (N_645,In_845,In_284);
and U646 (N_646,In_688,In_1357);
nor U647 (N_647,In_1303,In_47);
or U648 (N_648,In_18,In_1072);
nor U649 (N_649,In_917,In_651);
xnor U650 (N_650,In_15,In_254);
nand U651 (N_651,In_1497,In_1033);
nor U652 (N_652,In_1275,In_568);
and U653 (N_653,In_1170,In_951);
nor U654 (N_654,In_911,In_148);
xnor U655 (N_655,In_1318,In_483);
nor U656 (N_656,In_368,In_538);
xnor U657 (N_657,In_279,In_1396);
or U658 (N_658,In_259,In_1360);
nor U659 (N_659,In_12,In_137);
nor U660 (N_660,In_1247,In_704);
and U661 (N_661,In_1201,In_443);
nand U662 (N_662,In_73,In_41);
and U663 (N_663,In_1148,In_1324);
and U664 (N_664,In_1005,In_549);
xnor U665 (N_665,In_1294,In_718);
and U666 (N_666,In_6,In_649);
xor U667 (N_667,In_201,In_118);
and U668 (N_668,In_52,In_533);
xor U669 (N_669,In_617,In_637);
xnor U670 (N_670,In_1494,In_972);
or U671 (N_671,In_351,In_92);
nor U672 (N_672,In_501,In_783);
and U673 (N_673,In_1300,In_1128);
and U674 (N_674,In_432,In_909);
xnor U675 (N_675,In_261,In_440);
and U676 (N_676,In_433,In_865);
nand U677 (N_677,In_258,In_195);
xnor U678 (N_678,In_767,In_419);
or U679 (N_679,In_1431,In_103);
xnor U680 (N_680,In_745,In_356);
and U681 (N_681,In_1353,In_248);
or U682 (N_682,In_1185,In_1182);
nor U683 (N_683,In_570,In_846);
xor U684 (N_684,In_1283,In_1346);
or U685 (N_685,In_1195,In_1027);
nand U686 (N_686,In_1250,In_977);
nand U687 (N_687,In_493,In_211);
and U688 (N_688,In_269,In_1136);
or U689 (N_689,In_539,In_1257);
and U690 (N_690,In_707,In_695);
nand U691 (N_691,In_470,In_247);
and U692 (N_692,In_1204,In_1130);
nor U693 (N_693,In_640,In_1071);
nand U694 (N_694,In_608,In_884);
nor U695 (N_695,In_488,In_1485);
nor U696 (N_696,In_310,In_69);
xnor U697 (N_697,In_856,In_915);
and U698 (N_698,In_155,In_1388);
xor U699 (N_699,In_319,In_74);
nand U700 (N_700,In_519,In_392);
or U701 (N_701,In_1367,In_939);
or U702 (N_702,In_1015,In_1435);
nand U703 (N_703,In_388,In_446);
and U704 (N_704,In_1199,In_1169);
nor U705 (N_705,In_1192,In_1270);
nor U706 (N_706,In_697,In_1383);
xor U707 (N_707,In_1397,In_1221);
and U708 (N_708,In_569,In_194);
and U709 (N_709,In_1301,In_126);
nor U710 (N_710,In_1018,In_844);
xor U711 (N_711,In_982,In_1478);
or U712 (N_712,In_1375,In_1150);
and U713 (N_713,In_1184,In_31);
nand U714 (N_714,In_1215,In_910);
or U715 (N_715,In_124,In_926);
or U716 (N_716,In_311,In_333);
and U717 (N_717,In_482,In_925);
and U718 (N_718,In_83,In_377);
xnor U719 (N_719,In_1433,In_736);
nand U720 (N_720,In_1053,In_639);
and U721 (N_721,In_1373,In_109);
nor U722 (N_722,In_348,In_302);
and U723 (N_723,In_35,In_692);
xnor U724 (N_724,In_50,In_1496);
and U725 (N_725,In_1422,In_998);
nand U726 (N_726,In_930,In_674);
nand U727 (N_727,In_286,In_694);
and U728 (N_728,In_710,In_299);
or U729 (N_729,In_1110,In_212);
nor U730 (N_730,In_857,In_822);
nor U731 (N_731,In_873,In_108);
nor U732 (N_732,In_151,In_192);
or U733 (N_733,In_1056,In_371);
xor U734 (N_734,In_85,In_434);
or U735 (N_735,In_456,In_1338);
and U736 (N_736,In_1252,In_107);
and U737 (N_737,In_202,In_489);
nand U738 (N_738,In_366,In_113);
or U739 (N_739,In_681,In_281);
nor U740 (N_740,In_230,In_1);
or U741 (N_741,In_596,In_722);
nor U742 (N_742,In_787,In_336);
and U743 (N_743,In_1356,In_60);
or U744 (N_744,In_152,In_1418);
or U745 (N_745,In_949,In_271);
nor U746 (N_746,In_414,In_327);
and U747 (N_747,In_497,In_1153);
or U748 (N_748,In_294,In_693);
nor U749 (N_749,In_1021,In_149);
xnor U750 (N_750,In_689,In_258);
xnor U751 (N_751,In_1375,In_1175);
and U752 (N_752,In_19,In_592);
and U753 (N_753,In_1077,In_106);
and U754 (N_754,In_836,In_1402);
xnor U755 (N_755,In_1289,In_947);
and U756 (N_756,In_266,In_244);
nand U757 (N_757,In_371,In_1227);
or U758 (N_758,In_1174,In_66);
nor U759 (N_759,In_968,In_1406);
xnor U760 (N_760,In_773,In_1105);
nor U761 (N_761,In_406,In_456);
xnor U762 (N_762,In_1373,In_1269);
and U763 (N_763,In_961,In_315);
nor U764 (N_764,In_149,In_1295);
xnor U765 (N_765,In_1255,In_54);
or U766 (N_766,In_193,In_846);
or U767 (N_767,In_1279,In_81);
and U768 (N_768,In_1464,In_583);
xnor U769 (N_769,In_178,In_296);
nand U770 (N_770,In_1246,In_127);
nand U771 (N_771,In_410,In_749);
or U772 (N_772,In_497,In_707);
xnor U773 (N_773,In_981,In_248);
xor U774 (N_774,In_121,In_451);
xnor U775 (N_775,In_960,In_573);
nor U776 (N_776,In_2,In_961);
or U777 (N_777,In_241,In_1440);
nand U778 (N_778,In_799,In_1143);
or U779 (N_779,In_744,In_1479);
nor U780 (N_780,In_1078,In_1296);
or U781 (N_781,In_1113,In_1033);
nand U782 (N_782,In_1112,In_688);
or U783 (N_783,In_1062,In_83);
nor U784 (N_784,In_27,In_565);
nand U785 (N_785,In_1234,In_1357);
and U786 (N_786,In_681,In_103);
or U787 (N_787,In_27,In_178);
nand U788 (N_788,In_857,In_348);
nand U789 (N_789,In_173,In_789);
or U790 (N_790,In_1396,In_710);
xor U791 (N_791,In_635,In_14);
nor U792 (N_792,In_851,In_253);
xnor U793 (N_793,In_832,In_309);
and U794 (N_794,In_1316,In_1220);
xnor U795 (N_795,In_862,In_268);
nor U796 (N_796,In_279,In_1477);
or U797 (N_797,In_151,In_1367);
xor U798 (N_798,In_506,In_261);
nor U799 (N_799,In_560,In_1468);
nand U800 (N_800,In_1254,In_1470);
xor U801 (N_801,In_252,In_709);
or U802 (N_802,In_801,In_97);
and U803 (N_803,In_1115,In_740);
and U804 (N_804,In_1089,In_992);
nor U805 (N_805,In_771,In_46);
xor U806 (N_806,In_1215,In_1274);
and U807 (N_807,In_682,In_843);
xor U808 (N_808,In_191,In_773);
and U809 (N_809,In_1297,In_1277);
and U810 (N_810,In_192,In_152);
or U811 (N_811,In_1389,In_1157);
nand U812 (N_812,In_315,In_816);
nor U813 (N_813,In_513,In_782);
and U814 (N_814,In_9,In_945);
or U815 (N_815,In_11,In_869);
nor U816 (N_816,In_347,In_930);
and U817 (N_817,In_176,In_1360);
xnor U818 (N_818,In_234,In_926);
or U819 (N_819,In_842,In_677);
nand U820 (N_820,In_778,In_406);
and U821 (N_821,In_755,In_1228);
xor U822 (N_822,In_1265,In_863);
and U823 (N_823,In_199,In_298);
and U824 (N_824,In_1138,In_1409);
nor U825 (N_825,In_1006,In_991);
nand U826 (N_826,In_882,In_615);
nor U827 (N_827,In_1262,In_531);
or U828 (N_828,In_1356,In_645);
nand U829 (N_829,In_1375,In_1047);
nor U830 (N_830,In_188,In_1395);
xnor U831 (N_831,In_297,In_776);
or U832 (N_832,In_677,In_728);
nand U833 (N_833,In_879,In_1216);
and U834 (N_834,In_392,In_470);
and U835 (N_835,In_90,In_1086);
nand U836 (N_836,In_1269,In_1125);
and U837 (N_837,In_1379,In_1166);
nor U838 (N_838,In_385,In_1330);
or U839 (N_839,In_1122,In_89);
nand U840 (N_840,In_338,In_1023);
nand U841 (N_841,In_404,In_625);
and U842 (N_842,In_1203,In_117);
xor U843 (N_843,In_345,In_739);
nor U844 (N_844,In_685,In_350);
xor U845 (N_845,In_1213,In_855);
nor U846 (N_846,In_244,In_1417);
and U847 (N_847,In_1052,In_703);
xnor U848 (N_848,In_417,In_846);
xnor U849 (N_849,In_1429,In_577);
and U850 (N_850,In_174,In_1485);
nand U851 (N_851,In_1034,In_163);
xor U852 (N_852,In_272,In_222);
and U853 (N_853,In_871,In_1151);
nand U854 (N_854,In_1484,In_1223);
nand U855 (N_855,In_214,In_167);
nand U856 (N_856,In_0,In_1154);
xor U857 (N_857,In_3,In_951);
xor U858 (N_858,In_1489,In_1476);
xor U859 (N_859,In_1253,In_602);
nor U860 (N_860,In_1077,In_684);
or U861 (N_861,In_548,In_626);
nand U862 (N_862,In_1096,In_1283);
and U863 (N_863,In_1499,In_885);
nand U864 (N_864,In_1220,In_1038);
xnor U865 (N_865,In_761,In_1412);
nand U866 (N_866,In_1379,In_430);
xnor U867 (N_867,In_1499,In_374);
xnor U868 (N_868,In_986,In_664);
xor U869 (N_869,In_116,In_461);
xor U870 (N_870,In_442,In_743);
nor U871 (N_871,In_526,In_608);
xor U872 (N_872,In_561,In_758);
or U873 (N_873,In_524,In_1163);
or U874 (N_874,In_1301,In_138);
nor U875 (N_875,In_887,In_255);
or U876 (N_876,In_172,In_635);
nor U877 (N_877,In_302,In_968);
or U878 (N_878,In_130,In_1480);
or U879 (N_879,In_695,In_777);
nand U880 (N_880,In_363,In_828);
nand U881 (N_881,In_1446,In_1003);
nand U882 (N_882,In_54,In_279);
xor U883 (N_883,In_662,In_763);
or U884 (N_884,In_464,In_1048);
nand U885 (N_885,In_70,In_383);
or U886 (N_886,In_158,In_544);
or U887 (N_887,In_5,In_314);
xnor U888 (N_888,In_617,In_1430);
xor U889 (N_889,In_1383,In_1081);
xnor U890 (N_890,In_1127,In_325);
and U891 (N_891,In_623,In_321);
and U892 (N_892,In_374,In_433);
xor U893 (N_893,In_765,In_805);
xor U894 (N_894,In_808,In_102);
nor U895 (N_895,In_84,In_937);
nor U896 (N_896,In_514,In_276);
nand U897 (N_897,In_575,In_1313);
nor U898 (N_898,In_505,In_1378);
and U899 (N_899,In_171,In_666);
and U900 (N_900,In_880,In_1018);
or U901 (N_901,In_937,In_920);
nor U902 (N_902,In_596,In_1235);
nand U903 (N_903,In_441,In_774);
xor U904 (N_904,In_230,In_1386);
nand U905 (N_905,In_449,In_1289);
nor U906 (N_906,In_172,In_1274);
nand U907 (N_907,In_1358,In_1283);
nand U908 (N_908,In_43,In_1489);
xnor U909 (N_909,In_1018,In_374);
xnor U910 (N_910,In_677,In_298);
xnor U911 (N_911,In_1276,In_286);
or U912 (N_912,In_652,In_988);
and U913 (N_913,In_204,In_861);
nand U914 (N_914,In_653,In_1403);
and U915 (N_915,In_1253,In_164);
nor U916 (N_916,In_270,In_844);
nand U917 (N_917,In_372,In_1280);
and U918 (N_918,In_1491,In_105);
nand U919 (N_919,In_246,In_334);
xor U920 (N_920,In_913,In_1205);
or U921 (N_921,In_335,In_61);
and U922 (N_922,In_705,In_529);
xor U923 (N_923,In_623,In_967);
and U924 (N_924,In_47,In_890);
and U925 (N_925,In_660,In_114);
and U926 (N_926,In_860,In_1129);
nor U927 (N_927,In_616,In_6);
and U928 (N_928,In_483,In_261);
xor U929 (N_929,In_845,In_1233);
and U930 (N_930,In_1382,In_1018);
nor U931 (N_931,In_961,In_1192);
and U932 (N_932,In_875,In_538);
nor U933 (N_933,In_1227,In_1083);
and U934 (N_934,In_596,In_1385);
nand U935 (N_935,In_1027,In_1363);
nor U936 (N_936,In_324,In_1183);
and U937 (N_937,In_803,In_600);
nand U938 (N_938,In_1434,In_1311);
and U939 (N_939,In_38,In_1431);
xnor U940 (N_940,In_497,In_111);
nand U941 (N_941,In_1113,In_1484);
nand U942 (N_942,In_1489,In_153);
or U943 (N_943,In_273,In_291);
xnor U944 (N_944,In_48,In_151);
nand U945 (N_945,In_1303,In_89);
xor U946 (N_946,In_514,In_683);
and U947 (N_947,In_888,In_750);
or U948 (N_948,In_1021,In_575);
nor U949 (N_949,In_878,In_554);
nor U950 (N_950,In_740,In_238);
xnor U951 (N_951,In_96,In_1354);
nand U952 (N_952,In_145,In_144);
or U953 (N_953,In_828,In_922);
nand U954 (N_954,In_1118,In_823);
nand U955 (N_955,In_954,In_784);
nor U956 (N_956,In_179,In_1332);
and U957 (N_957,In_49,In_1498);
nor U958 (N_958,In_1012,In_63);
and U959 (N_959,In_878,In_459);
nor U960 (N_960,In_23,In_1122);
nor U961 (N_961,In_175,In_929);
nand U962 (N_962,In_44,In_0);
xnor U963 (N_963,In_962,In_1366);
nand U964 (N_964,In_144,In_1020);
xor U965 (N_965,In_1323,In_504);
or U966 (N_966,In_984,In_729);
xnor U967 (N_967,In_637,In_1097);
nand U968 (N_968,In_1055,In_24);
nor U969 (N_969,In_1224,In_355);
xnor U970 (N_970,In_90,In_724);
or U971 (N_971,In_384,In_400);
nor U972 (N_972,In_962,In_381);
nand U973 (N_973,In_810,In_187);
nor U974 (N_974,In_1079,In_792);
xnor U975 (N_975,In_847,In_44);
nand U976 (N_976,In_824,In_1069);
nor U977 (N_977,In_92,In_828);
or U978 (N_978,In_781,In_272);
and U979 (N_979,In_412,In_851);
or U980 (N_980,In_146,In_297);
or U981 (N_981,In_638,In_1001);
nor U982 (N_982,In_1165,In_448);
nand U983 (N_983,In_145,In_488);
nor U984 (N_984,In_1270,In_345);
nand U985 (N_985,In_1278,In_792);
nand U986 (N_986,In_335,In_1025);
or U987 (N_987,In_354,In_1235);
xor U988 (N_988,In_673,In_642);
nand U989 (N_989,In_753,In_1249);
nor U990 (N_990,In_914,In_860);
xor U991 (N_991,In_410,In_240);
or U992 (N_992,In_795,In_440);
nand U993 (N_993,In_119,In_1346);
and U994 (N_994,In_899,In_0);
and U995 (N_995,In_364,In_82);
or U996 (N_996,In_1138,In_1381);
or U997 (N_997,In_459,In_539);
xor U998 (N_998,In_124,In_1286);
xor U999 (N_999,In_143,In_1248);
and U1000 (N_1000,In_1196,In_411);
xnor U1001 (N_1001,In_1009,In_937);
nor U1002 (N_1002,In_1264,In_903);
xnor U1003 (N_1003,In_153,In_519);
and U1004 (N_1004,In_201,In_306);
or U1005 (N_1005,In_803,In_461);
xnor U1006 (N_1006,In_1097,In_53);
nand U1007 (N_1007,In_846,In_1035);
xnor U1008 (N_1008,In_286,In_736);
and U1009 (N_1009,In_281,In_355);
xnor U1010 (N_1010,In_58,In_180);
xor U1011 (N_1011,In_407,In_616);
nand U1012 (N_1012,In_497,In_1489);
or U1013 (N_1013,In_964,In_113);
or U1014 (N_1014,In_119,In_896);
nor U1015 (N_1015,In_685,In_1422);
xnor U1016 (N_1016,In_1190,In_913);
xnor U1017 (N_1017,In_1098,In_1086);
nand U1018 (N_1018,In_78,In_1110);
nor U1019 (N_1019,In_349,In_12);
xnor U1020 (N_1020,In_110,In_1401);
nor U1021 (N_1021,In_39,In_1288);
or U1022 (N_1022,In_305,In_650);
nor U1023 (N_1023,In_835,In_908);
or U1024 (N_1024,In_892,In_295);
nand U1025 (N_1025,In_1395,In_850);
or U1026 (N_1026,In_1005,In_327);
or U1027 (N_1027,In_39,In_182);
xnor U1028 (N_1028,In_163,In_434);
and U1029 (N_1029,In_170,In_258);
and U1030 (N_1030,In_569,In_1239);
nor U1031 (N_1031,In_1350,In_767);
nor U1032 (N_1032,In_126,In_503);
nand U1033 (N_1033,In_69,In_1394);
nor U1034 (N_1034,In_1006,In_208);
nand U1035 (N_1035,In_714,In_702);
and U1036 (N_1036,In_390,In_756);
and U1037 (N_1037,In_1281,In_1437);
or U1038 (N_1038,In_441,In_384);
or U1039 (N_1039,In_1488,In_1317);
nor U1040 (N_1040,In_1237,In_244);
and U1041 (N_1041,In_78,In_1272);
nand U1042 (N_1042,In_1455,In_171);
and U1043 (N_1043,In_1014,In_969);
and U1044 (N_1044,In_104,In_1389);
xnor U1045 (N_1045,In_1294,In_365);
xor U1046 (N_1046,In_154,In_686);
and U1047 (N_1047,In_737,In_26);
or U1048 (N_1048,In_259,In_1026);
xor U1049 (N_1049,In_448,In_519);
or U1050 (N_1050,In_851,In_1224);
and U1051 (N_1051,In_164,In_974);
and U1052 (N_1052,In_724,In_725);
nand U1053 (N_1053,In_1453,In_29);
or U1054 (N_1054,In_703,In_616);
nor U1055 (N_1055,In_1070,In_413);
nor U1056 (N_1056,In_1078,In_329);
nor U1057 (N_1057,In_1495,In_672);
and U1058 (N_1058,In_1212,In_232);
nand U1059 (N_1059,In_199,In_1292);
nand U1060 (N_1060,In_75,In_817);
nand U1061 (N_1061,In_486,In_638);
and U1062 (N_1062,In_1228,In_34);
nand U1063 (N_1063,In_612,In_970);
or U1064 (N_1064,In_0,In_883);
or U1065 (N_1065,In_1362,In_769);
or U1066 (N_1066,In_361,In_1203);
nand U1067 (N_1067,In_154,In_548);
xor U1068 (N_1068,In_638,In_1447);
or U1069 (N_1069,In_1190,In_587);
xnor U1070 (N_1070,In_1078,In_434);
xor U1071 (N_1071,In_1393,In_1100);
and U1072 (N_1072,In_346,In_910);
or U1073 (N_1073,In_621,In_168);
nor U1074 (N_1074,In_1191,In_166);
nor U1075 (N_1075,In_676,In_1100);
and U1076 (N_1076,In_473,In_1372);
and U1077 (N_1077,In_301,In_723);
nand U1078 (N_1078,In_1346,In_729);
nor U1079 (N_1079,In_743,In_290);
nand U1080 (N_1080,In_1034,In_78);
and U1081 (N_1081,In_1212,In_660);
nor U1082 (N_1082,In_51,In_429);
nand U1083 (N_1083,In_184,In_1090);
xor U1084 (N_1084,In_46,In_1291);
and U1085 (N_1085,In_79,In_793);
nor U1086 (N_1086,In_1411,In_1419);
nor U1087 (N_1087,In_766,In_937);
nor U1088 (N_1088,In_1260,In_1466);
xor U1089 (N_1089,In_149,In_1088);
xnor U1090 (N_1090,In_852,In_1306);
nor U1091 (N_1091,In_1318,In_1194);
xnor U1092 (N_1092,In_1241,In_1490);
nand U1093 (N_1093,In_800,In_1071);
nand U1094 (N_1094,In_82,In_1181);
nor U1095 (N_1095,In_1342,In_2);
or U1096 (N_1096,In_507,In_40);
and U1097 (N_1097,In_208,In_15);
xnor U1098 (N_1098,In_727,In_408);
or U1099 (N_1099,In_411,In_515);
or U1100 (N_1100,In_1234,In_688);
nor U1101 (N_1101,In_485,In_769);
xnor U1102 (N_1102,In_7,In_641);
xnor U1103 (N_1103,In_122,In_718);
nand U1104 (N_1104,In_658,In_830);
xor U1105 (N_1105,In_904,In_181);
and U1106 (N_1106,In_341,In_629);
nor U1107 (N_1107,In_1419,In_1318);
or U1108 (N_1108,In_1065,In_133);
nand U1109 (N_1109,In_399,In_544);
nor U1110 (N_1110,In_955,In_732);
nor U1111 (N_1111,In_661,In_929);
xor U1112 (N_1112,In_289,In_1373);
and U1113 (N_1113,In_1291,In_596);
xnor U1114 (N_1114,In_308,In_268);
xor U1115 (N_1115,In_1163,In_722);
xor U1116 (N_1116,In_543,In_1072);
xnor U1117 (N_1117,In_13,In_656);
and U1118 (N_1118,In_83,In_390);
nor U1119 (N_1119,In_832,In_243);
nor U1120 (N_1120,In_0,In_1428);
or U1121 (N_1121,In_1000,In_607);
xnor U1122 (N_1122,In_1085,In_1071);
nor U1123 (N_1123,In_98,In_1481);
xnor U1124 (N_1124,In_125,In_446);
xor U1125 (N_1125,In_805,In_243);
or U1126 (N_1126,In_541,In_1268);
nor U1127 (N_1127,In_1337,In_518);
and U1128 (N_1128,In_742,In_1472);
xnor U1129 (N_1129,In_1419,In_35);
and U1130 (N_1130,In_0,In_1131);
or U1131 (N_1131,In_540,In_831);
and U1132 (N_1132,In_836,In_1467);
and U1133 (N_1133,In_1098,In_192);
and U1134 (N_1134,In_273,In_292);
nor U1135 (N_1135,In_654,In_338);
nor U1136 (N_1136,In_457,In_311);
xor U1137 (N_1137,In_613,In_1416);
nor U1138 (N_1138,In_1002,In_919);
or U1139 (N_1139,In_2,In_688);
and U1140 (N_1140,In_292,In_625);
nor U1141 (N_1141,In_263,In_6);
nor U1142 (N_1142,In_1264,In_425);
and U1143 (N_1143,In_1007,In_258);
and U1144 (N_1144,In_1477,In_1240);
or U1145 (N_1145,In_34,In_938);
nand U1146 (N_1146,In_633,In_845);
and U1147 (N_1147,In_1470,In_774);
or U1148 (N_1148,In_55,In_575);
and U1149 (N_1149,In_284,In_1462);
and U1150 (N_1150,In_502,In_36);
nor U1151 (N_1151,In_34,In_1359);
or U1152 (N_1152,In_38,In_956);
and U1153 (N_1153,In_883,In_1412);
xnor U1154 (N_1154,In_142,In_1448);
xnor U1155 (N_1155,In_1472,In_890);
or U1156 (N_1156,In_919,In_1179);
or U1157 (N_1157,In_579,In_1179);
xnor U1158 (N_1158,In_1300,In_159);
or U1159 (N_1159,In_1180,In_241);
nor U1160 (N_1160,In_868,In_929);
and U1161 (N_1161,In_1226,In_1454);
xnor U1162 (N_1162,In_713,In_955);
nand U1163 (N_1163,In_1405,In_1169);
xnor U1164 (N_1164,In_102,In_1407);
and U1165 (N_1165,In_1452,In_1015);
or U1166 (N_1166,In_1401,In_431);
nand U1167 (N_1167,In_1148,In_1202);
or U1168 (N_1168,In_499,In_963);
or U1169 (N_1169,In_1480,In_1382);
nand U1170 (N_1170,In_199,In_797);
nand U1171 (N_1171,In_615,In_33);
and U1172 (N_1172,In_569,In_1039);
and U1173 (N_1173,In_793,In_678);
nand U1174 (N_1174,In_736,In_1081);
nor U1175 (N_1175,In_1173,In_575);
xor U1176 (N_1176,In_294,In_199);
and U1177 (N_1177,In_1179,In_1113);
or U1178 (N_1178,In_1228,In_769);
or U1179 (N_1179,In_60,In_858);
and U1180 (N_1180,In_887,In_835);
and U1181 (N_1181,In_483,In_775);
or U1182 (N_1182,In_416,In_1071);
nor U1183 (N_1183,In_393,In_88);
or U1184 (N_1184,In_757,In_16);
nor U1185 (N_1185,In_1206,In_240);
nor U1186 (N_1186,In_1358,In_400);
xnor U1187 (N_1187,In_56,In_688);
and U1188 (N_1188,In_1267,In_350);
xnor U1189 (N_1189,In_1064,In_991);
nand U1190 (N_1190,In_980,In_1290);
nand U1191 (N_1191,In_74,In_46);
or U1192 (N_1192,In_582,In_633);
nor U1193 (N_1193,In_324,In_1385);
nand U1194 (N_1194,In_106,In_406);
nand U1195 (N_1195,In_778,In_1206);
xnor U1196 (N_1196,In_1244,In_894);
nor U1197 (N_1197,In_1221,In_311);
and U1198 (N_1198,In_637,In_702);
and U1199 (N_1199,In_223,In_322);
xor U1200 (N_1200,In_1163,In_1226);
and U1201 (N_1201,In_857,In_1321);
and U1202 (N_1202,In_1030,In_823);
xnor U1203 (N_1203,In_681,In_1447);
and U1204 (N_1204,In_1292,In_554);
or U1205 (N_1205,In_1062,In_863);
and U1206 (N_1206,In_229,In_449);
nand U1207 (N_1207,In_675,In_274);
nand U1208 (N_1208,In_463,In_102);
xor U1209 (N_1209,In_74,In_1171);
and U1210 (N_1210,In_578,In_296);
nand U1211 (N_1211,In_1360,In_889);
xnor U1212 (N_1212,In_1075,In_63);
and U1213 (N_1213,In_1124,In_202);
xnor U1214 (N_1214,In_1022,In_1310);
nand U1215 (N_1215,In_118,In_1069);
or U1216 (N_1216,In_528,In_834);
nor U1217 (N_1217,In_432,In_1310);
and U1218 (N_1218,In_584,In_553);
and U1219 (N_1219,In_1101,In_762);
and U1220 (N_1220,In_789,In_823);
xor U1221 (N_1221,In_682,In_1013);
or U1222 (N_1222,In_801,In_54);
or U1223 (N_1223,In_145,In_502);
xor U1224 (N_1224,In_1043,In_119);
xnor U1225 (N_1225,In_740,In_245);
nand U1226 (N_1226,In_1002,In_953);
or U1227 (N_1227,In_358,In_699);
xnor U1228 (N_1228,In_1461,In_19);
and U1229 (N_1229,In_206,In_122);
nor U1230 (N_1230,In_772,In_600);
xor U1231 (N_1231,In_904,In_832);
xnor U1232 (N_1232,In_985,In_1058);
and U1233 (N_1233,In_1417,In_1052);
and U1234 (N_1234,In_897,In_236);
or U1235 (N_1235,In_476,In_1182);
and U1236 (N_1236,In_1021,In_1487);
or U1237 (N_1237,In_665,In_982);
nand U1238 (N_1238,In_874,In_578);
nor U1239 (N_1239,In_1229,In_1344);
nand U1240 (N_1240,In_667,In_1273);
nand U1241 (N_1241,In_706,In_417);
or U1242 (N_1242,In_621,In_285);
nor U1243 (N_1243,In_107,In_1308);
nand U1244 (N_1244,In_1485,In_1064);
nor U1245 (N_1245,In_914,In_63);
nor U1246 (N_1246,In_1358,In_640);
nor U1247 (N_1247,In_1497,In_722);
and U1248 (N_1248,In_423,In_959);
xnor U1249 (N_1249,In_1168,In_52);
or U1250 (N_1250,In_472,In_812);
and U1251 (N_1251,In_1071,In_463);
or U1252 (N_1252,In_1199,In_925);
nor U1253 (N_1253,In_1427,In_315);
or U1254 (N_1254,In_1221,In_197);
xnor U1255 (N_1255,In_1444,In_543);
or U1256 (N_1256,In_255,In_1396);
nor U1257 (N_1257,In_949,In_1456);
nor U1258 (N_1258,In_1448,In_481);
or U1259 (N_1259,In_407,In_12);
nand U1260 (N_1260,In_700,In_159);
nor U1261 (N_1261,In_1252,In_506);
xnor U1262 (N_1262,In_825,In_326);
nor U1263 (N_1263,In_22,In_1483);
nor U1264 (N_1264,In_1085,In_866);
and U1265 (N_1265,In_1208,In_1011);
nand U1266 (N_1266,In_298,In_1087);
and U1267 (N_1267,In_1183,In_29);
xnor U1268 (N_1268,In_907,In_311);
and U1269 (N_1269,In_873,In_91);
nand U1270 (N_1270,In_742,In_21);
nor U1271 (N_1271,In_1168,In_185);
and U1272 (N_1272,In_74,In_484);
and U1273 (N_1273,In_872,In_818);
and U1274 (N_1274,In_590,In_172);
nor U1275 (N_1275,In_1050,In_887);
nor U1276 (N_1276,In_826,In_117);
nor U1277 (N_1277,In_316,In_111);
nor U1278 (N_1278,In_1033,In_1405);
or U1279 (N_1279,In_11,In_178);
nor U1280 (N_1280,In_433,In_707);
nand U1281 (N_1281,In_314,In_1137);
or U1282 (N_1282,In_857,In_643);
nor U1283 (N_1283,In_280,In_328);
xnor U1284 (N_1284,In_1186,In_317);
nor U1285 (N_1285,In_228,In_1281);
or U1286 (N_1286,In_949,In_920);
xor U1287 (N_1287,In_188,In_50);
nand U1288 (N_1288,In_1476,In_1379);
or U1289 (N_1289,In_178,In_199);
or U1290 (N_1290,In_572,In_879);
nor U1291 (N_1291,In_1428,In_931);
or U1292 (N_1292,In_828,In_508);
xor U1293 (N_1293,In_670,In_817);
xnor U1294 (N_1294,In_1297,In_1089);
nand U1295 (N_1295,In_486,In_387);
nand U1296 (N_1296,In_33,In_351);
nand U1297 (N_1297,In_1331,In_1329);
xnor U1298 (N_1298,In_757,In_1462);
xor U1299 (N_1299,In_360,In_83);
nand U1300 (N_1300,In_570,In_170);
nor U1301 (N_1301,In_282,In_1004);
or U1302 (N_1302,In_1172,In_233);
or U1303 (N_1303,In_1039,In_1374);
nand U1304 (N_1304,In_32,In_641);
nand U1305 (N_1305,In_1286,In_1231);
nor U1306 (N_1306,In_939,In_1213);
nor U1307 (N_1307,In_1319,In_511);
and U1308 (N_1308,In_207,In_394);
nor U1309 (N_1309,In_1237,In_132);
nor U1310 (N_1310,In_941,In_615);
nand U1311 (N_1311,In_681,In_389);
or U1312 (N_1312,In_1232,In_1215);
or U1313 (N_1313,In_66,In_1151);
and U1314 (N_1314,In_960,In_831);
or U1315 (N_1315,In_813,In_1195);
or U1316 (N_1316,In_850,In_1469);
nor U1317 (N_1317,In_305,In_541);
and U1318 (N_1318,In_146,In_46);
and U1319 (N_1319,In_143,In_1385);
nand U1320 (N_1320,In_567,In_456);
or U1321 (N_1321,In_187,In_172);
xor U1322 (N_1322,In_42,In_828);
nor U1323 (N_1323,In_433,In_980);
nand U1324 (N_1324,In_151,In_870);
nor U1325 (N_1325,In_667,In_446);
nand U1326 (N_1326,In_999,In_167);
and U1327 (N_1327,In_288,In_834);
xnor U1328 (N_1328,In_633,In_807);
and U1329 (N_1329,In_969,In_878);
xnor U1330 (N_1330,In_542,In_1153);
or U1331 (N_1331,In_1474,In_609);
xor U1332 (N_1332,In_1020,In_309);
nand U1333 (N_1333,In_317,In_1421);
xor U1334 (N_1334,In_541,In_1389);
nor U1335 (N_1335,In_1108,In_571);
nor U1336 (N_1336,In_416,In_390);
nor U1337 (N_1337,In_465,In_615);
and U1338 (N_1338,In_711,In_470);
or U1339 (N_1339,In_533,In_1389);
nand U1340 (N_1340,In_9,In_1049);
and U1341 (N_1341,In_1077,In_1146);
and U1342 (N_1342,In_751,In_1013);
xnor U1343 (N_1343,In_559,In_843);
xnor U1344 (N_1344,In_1149,In_1209);
nor U1345 (N_1345,In_476,In_320);
or U1346 (N_1346,In_1464,In_79);
xor U1347 (N_1347,In_705,In_1362);
nor U1348 (N_1348,In_1286,In_49);
nand U1349 (N_1349,In_72,In_535);
nand U1350 (N_1350,In_298,In_839);
xor U1351 (N_1351,In_961,In_1359);
xnor U1352 (N_1352,In_127,In_1468);
xnor U1353 (N_1353,In_1438,In_507);
xor U1354 (N_1354,In_260,In_1416);
nor U1355 (N_1355,In_969,In_887);
or U1356 (N_1356,In_56,In_476);
xor U1357 (N_1357,In_276,In_1469);
nor U1358 (N_1358,In_116,In_314);
or U1359 (N_1359,In_378,In_347);
or U1360 (N_1360,In_1499,In_1471);
and U1361 (N_1361,In_370,In_417);
nor U1362 (N_1362,In_668,In_172);
or U1363 (N_1363,In_184,In_56);
nor U1364 (N_1364,In_1430,In_1351);
or U1365 (N_1365,In_88,In_538);
and U1366 (N_1366,In_408,In_23);
nor U1367 (N_1367,In_1098,In_1495);
nand U1368 (N_1368,In_583,In_535);
and U1369 (N_1369,In_537,In_1447);
nand U1370 (N_1370,In_1121,In_1470);
nor U1371 (N_1371,In_53,In_1441);
nor U1372 (N_1372,In_1093,In_1364);
nor U1373 (N_1373,In_1347,In_1371);
nand U1374 (N_1374,In_703,In_797);
xnor U1375 (N_1375,In_1347,In_1225);
or U1376 (N_1376,In_125,In_646);
nand U1377 (N_1377,In_1057,In_1194);
and U1378 (N_1378,In_1209,In_97);
or U1379 (N_1379,In_1055,In_188);
xor U1380 (N_1380,In_665,In_1086);
or U1381 (N_1381,In_1275,In_1264);
nor U1382 (N_1382,In_209,In_373);
nand U1383 (N_1383,In_779,In_1200);
and U1384 (N_1384,In_607,In_1483);
or U1385 (N_1385,In_631,In_1176);
nor U1386 (N_1386,In_857,In_604);
nand U1387 (N_1387,In_42,In_860);
xor U1388 (N_1388,In_161,In_35);
nor U1389 (N_1389,In_1432,In_309);
nor U1390 (N_1390,In_139,In_892);
nand U1391 (N_1391,In_290,In_782);
nand U1392 (N_1392,In_589,In_694);
nand U1393 (N_1393,In_678,In_681);
nand U1394 (N_1394,In_23,In_966);
or U1395 (N_1395,In_13,In_28);
and U1396 (N_1396,In_168,In_9);
and U1397 (N_1397,In_268,In_594);
or U1398 (N_1398,In_757,In_377);
or U1399 (N_1399,In_298,In_244);
nand U1400 (N_1400,In_685,In_1086);
nor U1401 (N_1401,In_666,In_1183);
and U1402 (N_1402,In_1218,In_12);
and U1403 (N_1403,In_280,In_606);
nand U1404 (N_1404,In_770,In_314);
nor U1405 (N_1405,In_1251,In_375);
nor U1406 (N_1406,In_505,In_847);
nand U1407 (N_1407,In_358,In_558);
or U1408 (N_1408,In_1373,In_713);
nor U1409 (N_1409,In_931,In_1424);
and U1410 (N_1410,In_1414,In_1201);
or U1411 (N_1411,In_18,In_464);
or U1412 (N_1412,In_828,In_1009);
xnor U1413 (N_1413,In_93,In_403);
xor U1414 (N_1414,In_466,In_748);
or U1415 (N_1415,In_430,In_1346);
and U1416 (N_1416,In_336,In_534);
xnor U1417 (N_1417,In_608,In_23);
xor U1418 (N_1418,In_374,In_104);
or U1419 (N_1419,In_1316,In_1060);
or U1420 (N_1420,In_1277,In_931);
xnor U1421 (N_1421,In_1433,In_176);
xnor U1422 (N_1422,In_427,In_138);
or U1423 (N_1423,In_891,In_209);
nor U1424 (N_1424,In_1302,In_1313);
nor U1425 (N_1425,In_670,In_19);
nor U1426 (N_1426,In_1468,In_1208);
or U1427 (N_1427,In_1040,In_480);
or U1428 (N_1428,In_12,In_1203);
xnor U1429 (N_1429,In_1279,In_1080);
nor U1430 (N_1430,In_1419,In_1056);
or U1431 (N_1431,In_54,In_889);
and U1432 (N_1432,In_62,In_548);
or U1433 (N_1433,In_463,In_838);
xor U1434 (N_1434,In_1191,In_1051);
xnor U1435 (N_1435,In_871,In_511);
or U1436 (N_1436,In_144,In_1152);
nand U1437 (N_1437,In_1379,In_1194);
xor U1438 (N_1438,In_142,In_837);
xnor U1439 (N_1439,In_1375,In_767);
nand U1440 (N_1440,In_1046,In_1390);
nor U1441 (N_1441,In_687,In_1198);
xnor U1442 (N_1442,In_939,In_784);
nand U1443 (N_1443,In_1238,In_359);
nand U1444 (N_1444,In_211,In_1088);
or U1445 (N_1445,In_271,In_36);
and U1446 (N_1446,In_724,In_960);
xnor U1447 (N_1447,In_726,In_572);
xnor U1448 (N_1448,In_1350,In_938);
xor U1449 (N_1449,In_995,In_1320);
nand U1450 (N_1450,In_1475,In_93);
xnor U1451 (N_1451,In_1046,In_676);
nor U1452 (N_1452,In_772,In_807);
xor U1453 (N_1453,In_462,In_1125);
nand U1454 (N_1454,In_1091,In_9);
and U1455 (N_1455,In_1319,In_174);
and U1456 (N_1456,In_1184,In_10);
nor U1457 (N_1457,In_762,In_1385);
xor U1458 (N_1458,In_579,In_504);
nand U1459 (N_1459,In_85,In_484);
or U1460 (N_1460,In_1282,In_331);
or U1461 (N_1461,In_934,In_1237);
nand U1462 (N_1462,In_1096,In_1099);
or U1463 (N_1463,In_158,In_58);
and U1464 (N_1464,In_1036,In_26);
xnor U1465 (N_1465,In_1289,In_140);
xnor U1466 (N_1466,In_580,In_431);
and U1467 (N_1467,In_1442,In_421);
nor U1468 (N_1468,In_1314,In_317);
or U1469 (N_1469,In_253,In_1231);
nor U1470 (N_1470,In_785,In_1048);
nand U1471 (N_1471,In_493,In_344);
and U1472 (N_1472,In_1283,In_390);
xor U1473 (N_1473,In_1404,In_1283);
nand U1474 (N_1474,In_938,In_301);
or U1475 (N_1475,In_606,In_1457);
xor U1476 (N_1476,In_1458,In_1001);
nand U1477 (N_1477,In_1466,In_429);
nand U1478 (N_1478,In_1386,In_1249);
or U1479 (N_1479,In_1427,In_1085);
nand U1480 (N_1480,In_983,In_467);
or U1481 (N_1481,In_1147,In_1115);
nand U1482 (N_1482,In_148,In_958);
nor U1483 (N_1483,In_1444,In_1169);
xnor U1484 (N_1484,In_1147,In_1333);
xnor U1485 (N_1485,In_888,In_301);
xnor U1486 (N_1486,In_602,In_730);
and U1487 (N_1487,In_1106,In_133);
or U1488 (N_1488,In_587,In_1297);
and U1489 (N_1489,In_79,In_831);
xor U1490 (N_1490,In_757,In_899);
nand U1491 (N_1491,In_24,In_1379);
xor U1492 (N_1492,In_61,In_297);
nor U1493 (N_1493,In_217,In_189);
nand U1494 (N_1494,In_357,In_459);
nor U1495 (N_1495,In_515,In_202);
or U1496 (N_1496,In_899,In_333);
and U1497 (N_1497,In_817,In_93);
nand U1498 (N_1498,In_1475,In_1010);
nand U1499 (N_1499,In_556,In_1052);
xor U1500 (N_1500,N_204,N_1441);
or U1501 (N_1501,N_99,N_723);
nand U1502 (N_1502,N_719,N_1077);
or U1503 (N_1503,N_1280,N_937);
and U1504 (N_1504,N_1415,N_1294);
xor U1505 (N_1505,N_1495,N_61);
nand U1506 (N_1506,N_57,N_1424);
nand U1507 (N_1507,N_401,N_364);
nand U1508 (N_1508,N_358,N_690);
nor U1509 (N_1509,N_1497,N_1390);
xnor U1510 (N_1510,N_297,N_760);
nand U1511 (N_1511,N_1364,N_720);
nor U1512 (N_1512,N_1370,N_276);
and U1513 (N_1513,N_538,N_970);
xnor U1514 (N_1514,N_1314,N_1317);
xor U1515 (N_1515,N_118,N_783);
xor U1516 (N_1516,N_821,N_447);
nand U1517 (N_1517,N_901,N_740);
nand U1518 (N_1518,N_109,N_329);
nand U1519 (N_1519,N_1188,N_1339);
nand U1520 (N_1520,N_603,N_463);
nand U1521 (N_1521,N_1340,N_348);
nand U1522 (N_1522,N_1355,N_1422);
xor U1523 (N_1523,N_1050,N_751);
nand U1524 (N_1524,N_889,N_859);
xor U1525 (N_1525,N_0,N_1036);
xnor U1526 (N_1526,N_1300,N_2);
nand U1527 (N_1527,N_1047,N_707);
nor U1528 (N_1528,N_1200,N_1282);
or U1529 (N_1529,N_939,N_134);
xor U1530 (N_1530,N_1253,N_1167);
and U1531 (N_1531,N_808,N_1131);
nor U1532 (N_1532,N_211,N_1008);
or U1533 (N_1533,N_727,N_570);
or U1534 (N_1534,N_1134,N_749);
xor U1535 (N_1535,N_917,N_1315);
xor U1536 (N_1536,N_541,N_1025);
xnor U1537 (N_1537,N_1151,N_1046);
nor U1538 (N_1538,N_169,N_129);
xor U1539 (N_1539,N_1243,N_1160);
xor U1540 (N_1540,N_652,N_24);
xor U1541 (N_1541,N_346,N_738);
and U1542 (N_1542,N_590,N_746);
nor U1543 (N_1543,N_1003,N_170);
xor U1544 (N_1544,N_395,N_31);
and U1545 (N_1545,N_102,N_1069);
xor U1546 (N_1546,N_1092,N_174);
and U1547 (N_1547,N_934,N_950);
xor U1548 (N_1548,N_639,N_16);
and U1549 (N_1549,N_869,N_226);
or U1550 (N_1550,N_268,N_547);
or U1551 (N_1551,N_1186,N_1255);
xnor U1552 (N_1552,N_1017,N_993);
or U1553 (N_1553,N_112,N_38);
or U1554 (N_1554,N_1296,N_920);
or U1555 (N_1555,N_745,N_1499);
nor U1556 (N_1556,N_145,N_958);
xor U1557 (N_1557,N_155,N_218);
or U1558 (N_1558,N_1265,N_788);
or U1559 (N_1559,N_514,N_448);
or U1560 (N_1560,N_184,N_195);
or U1561 (N_1561,N_1018,N_1341);
or U1562 (N_1562,N_1348,N_55);
nand U1563 (N_1563,N_972,N_221);
and U1564 (N_1564,N_445,N_483);
xnor U1565 (N_1565,N_847,N_225);
xnor U1566 (N_1566,N_188,N_777);
xor U1567 (N_1567,N_1100,N_894);
or U1568 (N_1568,N_1041,N_1237);
nand U1569 (N_1569,N_799,N_905);
and U1570 (N_1570,N_78,N_177);
nor U1571 (N_1571,N_254,N_884);
xnor U1572 (N_1572,N_273,N_668);
nor U1573 (N_1573,N_1325,N_1185);
nor U1574 (N_1574,N_1454,N_571);
or U1575 (N_1575,N_864,N_655);
nand U1576 (N_1576,N_602,N_1079);
nand U1577 (N_1577,N_1274,N_667);
or U1578 (N_1578,N_1356,N_695);
and U1579 (N_1579,N_949,N_822);
nand U1580 (N_1580,N_451,N_1273);
nand U1581 (N_1581,N_604,N_191);
or U1582 (N_1582,N_1388,N_146);
nor U1583 (N_1583,N_1303,N_795);
nand U1584 (N_1584,N_1342,N_705);
xnor U1585 (N_1585,N_456,N_1106);
and U1586 (N_1586,N_614,N_510);
xor U1587 (N_1587,N_836,N_1035);
nand U1588 (N_1588,N_759,N_71);
or U1589 (N_1589,N_1074,N_637);
nor U1590 (N_1590,N_1085,N_730);
or U1591 (N_1591,N_1399,N_56);
or U1592 (N_1592,N_416,N_792);
nor U1593 (N_1593,N_13,N_1344);
or U1594 (N_1594,N_1235,N_1097);
and U1595 (N_1595,N_842,N_918);
nor U1596 (N_1596,N_1288,N_203);
nor U1597 (N_1597,N_820,N_1444);
or U1598 (N_1598,N_224,N_93);
nor U1599 (N_1599,N_839,N_167);
or U1600 (N_1600,N_1406,N_1216);
xor U1601 (N_1601,N_397,N_1128);
nand U1602 (N_1602,N_1164,N_527);
nor U1603 (N_1603,N_815,N_1467);
nor U1604 (N_1604,N_517,N_44);
or U1605 (N_1605,N_158,N_1051);
nand U1606 (N_1606,N_797,N_682);
and U1607 (N_1607,N_828,N_83);
or U1608 (N_1608,N_311,N_940);
and U1609 (N_1609,N_1391,N_1292);
or U1610 (N_1610,N_1295,N_328);
or U1611 (N_1611,N_744,N_278);
nor U1612 (N_1612,N_251,N_1335);
nor U1613 (N_1613,N_307,N_1439);
xor U1614 (N_1614,N_183,N_734);
or U1615 (N_1615,N_239,N_313);
nor U1616 (N_1616,N_59,N_953);
nand U1617 (N_1617,N_319,N_1385);
nor U1618 (N_1618,N_805,N_235);
xnor U1619 (N_1619,N_583,N_1081);
xor U1620 (N_1620,N_803,N_874);
nor U1621 (N_1621,N_1373,N_646);
nand U1622 (N_1622,N_504,N_561);
or U1623 (N_1623,N_1484,N_1456);
and U1624 (N_1624,N_539,N_84);
nor U1625 (N_1625,N_30,N_237);
and U1626 (N_1626,N_1459,N_241);
or U1627 (N_1627,N_114,N_1493);
xnor U1628 (N_1628,N_1175,N_1037);
and U1629 (N_1629,N_1223,N_1103);
nand U1630 (N_1630,N_1093,N_281);
or U1631 (N_1631,N_280,N_1011);
nand U1632 (N_1632,N_1065,N_710);
xnor U1633 (N_1633,N_338,N_645);
nand U1634 (N_1634,N_810,N_22);
nand U1635 (N_1635,N_689,N_989);
nor U1636 (N_1636,N_1016,N_932);
nor U1637 (N_1637,N_1154,N_1189);
and U1638 (N_1638,N_8,N_852);
nor U1639 (N_1639,N_677,N_524);
or U1640 (N_1640,N_1457,N_1451);
or U1641 (N_1641,N_574,N_706);
xor U1642 (N_1642,N_628,N_1268);
nor U1643 (N_1643,N_618,N_1118);
and U1644 (N_1644,N_1312,N_819);
nor U1645 (N_1645,N_1334,N_587);
nor U1646 (N_1646,N_496,N_107);
xnor U1647 (N_1647,N_493,N_785);
xor U1648 (N_1648,N_50,N_800);
and U1649 (N_1649,N_178,N_899);
nand U1650 (N_1650,N_1115,N_67);
nor U1651 (N_1651,N_398,N_1258);
nand U1652 (N_1652,N_79,N_1209);
nor U1653 (N_1653,N_1056,N_43);
nand U1654 (N_1654,N_1030,N_1172);
xor U1655 (N_1655,N_248,N_1453);
or U1656 (N_1656,N_906,N_190);
nand U1657 (N_1657,N_875,N_1326);
or U1658 (N_1658,N_314,N_522);
nand U1659 (N_1659,N_555,N_1087);
nand U1660 (N_1660,N_334,N_1313);
or U1661 (N_1661,N_1310,N_990);
xnor U1662 (N_1662,N_1020,N_530);
xnor U1663 (N_1663,N_635,N_217);
nand U1664 (N_1664,N_1032,N_912);
nor U1665 (N_1665,N_1187,N_1460);
and U1666 (N_1666,N_698,N_1381);
nand U1667 (N_1667,N_850,N_630);
and U1668 (N_1668,N_1483,N_392);
or U1669 (N_1669,N_176,N_680);
and U1670 (N_1670,N_975,N_1021);
nor U1671 (N_1671,N_1193,N_625);
nor U1672 (N_1672,N_500,N_888);
nor U1673 (N_1673,N_1336,N_1208);
xor U1674 (N_1674,N_1,N_263);
nor U1675 (N_1675,N_438,N_1099);
or U1676 (N_1676,N_110,N_141);
nor U1677 (N_1677,N_76,N_582);
and U1678 (N_1678,N_165,N_293);
or U1679 (N_1679,N_814,N_48);
xor U1680 (N_1680,N_87,N_215);
or U1681 (N_1681,N_37,N_1220);
or U1682 (N_1682,N_113,N_856);
nand U1683 (N_1683,N_283,N_1284);
nor U1684 (N_1684,N_351,N_536);
nand U1685 (N_1685,N_1307,N_1418);
xor U1686 (N_1686,N_41,N_753);
or U1687 (N_1687,N_647,N_11);
xnor U1688 (N_1688,N_1170,N_832);
and U1689 (N_1689,N_434,N_412);
nor U1690 (N_1690,N_432,N_1423);
and U1691 (N_1691,N_909,N_767);
nor U1692 (N_1692,N_429,N_757);
nand U1693 (N_1693,N_396,N_1133);
and U1694 (N_1694,N_1407,N_355);
nor U1695 (N_1695,N_75,N_830);
xor U1696 (N_1696,N_5,N_1114);
xor U1697 (N_1697,N_615,N_961);
or U1698 (N_1698,N_1014,N_378);
and U1699 (N_1699,N_1194,N_900);
nor U1700 (N_1700,N_361,N_954);
xor U1701 (N_1701,N_1205,N_763);
and U1702 (N_1702,N_755,N_729);
nor U1703 (N_1703,N_413,N_947);
nor U1704 (N_1704,N_229,N_1135);
xnor U1705 (N_1705,N_252,N_722);
and U1706 (N_1706,N_857,N_175);
nor U1707 (N_1707,N_1156,N_1171);
nor U1708 (N_1708,N_1318,N_528);
nor U1709 (N_1709,N_1221,N_60);
xnor U1710 (N_1710,N_1236,N_648);
nand U1711 (N_1711,N_736,N_501);
and U1712 (N_1712,N_966,N_1277);
xnor U1713 (N_1713,N_607,N_1083);
nor U1714 (N_1714,N_408,N_904);
nand U1715 (N_1715,N_851,N_272);
or U1716 (N_1716,N_593,N_39);
xor U1717 (N_1717,N_1230,N_1159);
xnor U1718 (N_1718,N_344,N_1143);
or U1719 (N_1719,N_312,N_521);
xnor U1720 (N_1720,N_131,N_216);
or U1721 (N_1721,N_207,N_1239);
nand U1722 (N_1722,N_27,N_266);
and U1723 (N_1723,N_168,N_622);
nand U1724 (N_1724,N_1094,N_1398);
nand U1725 (N_1725,N_1440,N_1420);
and U1726 (N_1726,N_249,N_465);
and U1727 (N_1727,N_925,N_1244);
or U1728 (N_1728,N_1110,N_936);
xor U1729 (N_1729,N_1007,N_1357);
nand U1730 (N_1730,N_1449,N_807);
and U1731 (N_1731,N_377,N_686);
xor U1732 (N_1732,N_988,N_236);
nand U1733 (N_1733,N_854,N_772);
nor U1734 (N_1734,N_985,N_509);
and U1735 (N_1735,N_1177,N_316);
nand U1736 (N_1736,N_1086,N_488);
nor U1737 (N_1737,N_212,N_101);
or U1738 (N_1738,N_127,N_605);
xor U1739 (N_1739,N_1199,N_879);
and U1740 (N_1740,N_654,N_437);
nor U1741 (N_1741,N_1071,N_1349);
xor U1742 (N_1742,N_1026,N_1168);
or U1743 (N_1743,N_208,N_1104);
and U1744 (N_1744,N_778,N_478);
and U1745 (N_1745,N_1252,N_1465);
or U1746 (N_1746,N_944,N_157);
and U1747 (N_1747,N_844,N_189);
nand U1748 (N_1748,N_1363,N_490);
or U1749 (N_1749,N_484,N_1322);
nand U1750 (N_1750,N_161,N_773);
and U1751 (N_1751,N_994,N_1138);
xnor U1752 (N_1752,N_711,N_595);
xor U1753 (N_1753,N_81,N_731);
nor U1754 (N_1754,N_264,N_223);
nand U1755 (N_1755,N_568,N_846);
nand U1756 (N_1756,N_634,N_997);
nand U1757 (N_1757,N_424,N_1090);
xnor U1758 (N_1758,N_943,N_880);
and U1759 (N_1759,N_640,N_505);
nand U1760 (N_1760,N_942,N_3);
nand U1761 (N_1761,N_90,N_86);
xnor U1762 (N_1762,N_1147,N_1320);
or U1763 (N_1763,N_182,N_386);
nand U1764 (N_1764,N_633,N_467);
xnor U1765 (N_1765,N_716,N_1414);
and U1766 (N_1766,N_829,N_578);
or U1767 (N_1767,N_750,N_368);
and U1768 (N_1768,N_1436,N_882);
xor U1769 (N_1769,N_580,N_1468);
xnor U1770 (N_1770,N_153,N_956);
xor U1771 (N_1771,N_597,N_119);
xnor U1772 (N_1772,N_739,N_1287);
and U1773 (N_1773,N_480,N_643);
and U1774 (N_1774,N_331,N_627);
and U1775 (N_1775,N_1345,N_552);
and U1776 (N_1776,N_1000,N_173);
xor U1777 (N_1777,N_291,N_585);
nand U1778 (N_1778,N_411,N_601);
and U1779 (N_1779,N_572,N_135);
and U1780 (N_1780,N_310,N_1019);
or U1781 (N_1781,N_1263,N_369);
nor U1782 (N_1782,N_1217,N_964);
and U1783 (N_1783,N_42,N_1197);
and U1784 (N_1784,N_733,N_1149);
nand U1785 (N_1785,N_573,N_147);
xnor U1786 (N_1786,N_325,N_515);
nor U1787 (N_1787,N_1376,N_330);
and U1788 (N_1788,N_352,N_1285);
or U1789 (N_1789,N_980,N_339);
or U1790 (N_1790,N_518,N_532);
and U1791 (N_1791,N_1266,N_219);
nand U1792 (N_1792,N_1247,N_1129);
and U1793 (N_1793,N_206,N_1224);
or U1794 (N_1794,N_1359,N_609);
or U1795 (N_1795,N_124,N_679);
xnor U1796 (N_1796,N_712,N_337);
xor U1797 (N_1797,N_370,N_1146);
or U1798 (N_1798,N_1137,N_1121);
nand U1799 (N_1799,N_271,N_1222);
xor U1800 (N_1800,N_477,N_1347);
or U1801 (N_1801,N_475,N_274);
and U1802 (N_1802,N_360,N_567);
and U1803 (N_1803,N_611,N_40);
or U1804 (N_1804,N_741,N_1487);
or U1805 (N_1805,N_775,N_696);
nand U1806 (N_1806,N_959,N_560);
xor U1807 (N_1807,N_426,N_1397);
xnor U1808 (N_1808,N_479,N_952);
or U1809 (N_1809,N_95,N_315);
and U1810 (N_1810,N_529,N_1181);
xnor U1811 (N_1811,N_1157,N_1057);
nand U1812 (N_1812,N_1067,N_70);
xnor U1813 (N_1813,N_623,N_1203);
xnor U1814 (N_1814,N_94,N_304);
nand U1815 (N_1815,N_833,N_1232);
nor U1816 (N_1816,N_793,N_402);
nand U1817 (N_1817,N_1346,N_809);
nor U1818 (N_1818,N_559,N_659);
or U1819 (N_1819,N_1338,N_902);
xor U1820 (N_1820,N_1212,N_1384);
or U1821 (N_1821,N_1276,N_452);
nand U1822 (N_1822,N_631,N_1109);
nand U1823 (N_1823,N_1429,N_1098);
xor U1824 (N_1824,N_1176,N_1096);
and U1825 (N_1825,N_1202,N_495);
xnor U1826 (N_1826,N_1492,N_813);
or U1827 (N_1827,N_979,N_747);
or U1828 (N_1828,N_63,N_841);
and U1829 (N_1829,N_1053,N_636);
or U1830 (N_1830,N_460,N_503);
xor U1831 (N_1831,N_1078,N_100);
or U1832 (N_1832,N_1257,N_258);
nand U1833 (N_1833,N_1219,N_861);
and U1834 (N_1834,N_1264,N_592);
xnor U1835 (N_1835,N_1015,N_485);
xnor U1836 (N_1836,N_928,N_117);
and U1837 (N_1837,N_752,N_49);
xor U1838 (N_1838,N_149,N_929);
xor U1839 (N_1839,N_796,N_1089);
nor U1840 (N_1840,N_692,N_1042);
or U1841 (N_1841,N_789,N_1238);
or U1842 (N_1842,N_921,N_1293);
xnor U1843 (N_1843,N_366,N_1463);
nand U1844 (N_1844,N_382,N_758);
and U1845 (N_1845,N_853,N_1437);
or U1846 (N_1846,N_1366,N_1102);
and U1847 (N_1847,N_265,N_768);
and U1848 (N_1848,N_581,N_193);
xnor U1849 (N_1849,N_210,N_951);
or U1850 (N_1850,N_825,N_380);
nand U1851 (N_1851,N_1240,N_694);
and U1852 (N_1852,N_728,N_1228);
or U1853 (N_1853,N_976,N_1301);
and U1854 (N_1854,N_761,N_1445);
or U1855 (N_1855,N_130,N_1153);
or U1856 (N_1856,N_1248,N_660);
nor U1857 (N_1857,N_446,N_1330);
and U1858 (N_1858,N_1408,N_253);
nand U1859 (N_1859,N_688,N_23);
nand U1860 (N_1860,N_1361,N_69);
and U1861 (N_1861,N_473,N_244);
xnor U1862 (N_1862,N_1319,N_405);
and U1863 (N_1863,N_642,N_626);
nand U1864 (N_1864,N_250,N_306);
xor U1865 (N_1865,N_946,N_1179);
and U1866 (N_1866,N_790,N_267);
or U1867 (N_1867,N_556,N_665);
nor U1868 (N_1868,N_1464,N_1490);
xor U1869 (N_1869,N_1485,N_897);
or U1870 (N_1870,N_128,N_19);
or U1871 (N_1871,N_666,N_1082);
or U1872 (N_1872,N_323,N_748);
and U1873 (N_1873,N_663,N_1062);
xnor U1874 (N_1874,N_1141,N_1365);
xor U1875 (N_1875,N_624,N_1117);
and U1876 (N_1876,N_1132,N_1058);
and U1877 (N_1877,N_1120,N_476);
and U1878 (N_1878,N_58,N_1417);
xor U1879 (N_1879,N_919,N_298);
nor U1880 (N_1880,N_1479,N_550);
or U1881 (N_1881,N_343,N_1059);
xor U1882 (N_1882,N_120,N_1161);
or U1883 (N_1883,N_908,N_471);
nand U1884 (N_1884,N_1350,N_82);
and U1885 (N_1885,N_1169,N_322);
nor U1886 (N_1886,N_213,N_1130);
xor U1887 (N_1887,N_983,N_340);
nor U1888 (N_1888,N_542,N_292);
nand U1889 (N_1889,N_1155,N_1486);
or U1890 (N_1890,N_357,N_629);
nand U1891 (N_1891,N_1375,N_1111);
nand U1892 (N_1892,N_923,N_974);
nor U1893 (N_1893,N_1358,N_735);
and U1894 (N_1894,N_1329,N_669);
nor U1895 (N_1895,N_1494,N_511);
or U1896 (N_1896,N_1060,N_1038);
xor U1897 (N_1897,N_46,N_1166);
xnor U1898 (N_1898,N_98,N_286);
and U1899 (N_1899,N_1070,N_898);
or U1900 (N_1900,N_1144,N_222);
nand U1901 (N_1901,N_1412,N_599);
xor U1902 (N_1902,N_1040,N_1045);
or U1903 (N_1903,N_1229,N_324);
xor U1904 (N_1904,N_890,N_726);
and U1905 (N_1905,N_649,N_867);
nand U1906 (N_1906,N_610,N_776);
xor U1907 (N_1907,N_1165,N_289);
or U1908 (N_1908,N_1068,N_415);
and U1909 (N_1909,N_474,N_658);
xnor U1910 (N_1910,N_116,N_986);
nor U1911 (N_1911,N_246,N_673);
or U1912 (N_1912,N_1427,N_29);
xnor U1913 (N_1913,N_1409,N_638);
and U1914 (N_1914,N_1369,N_240);
xor U1915 (N_1915,N_417,N_442);
or U1916 (N_1916,N_1249,N_926);
nand U1917 (N_1917,N_896,N_73);
and U1918 (N_1918,N_259,N_591);
xor U1919 (N_1919,N_25,N_742);
and U1920 (N_1920,N_754,N_1489);
and U1921 (N_1921,N_179,N_598);
or U1922 (N_1922,N_718,N_523);
nand U1923 (N_1923,N_1145,N_227);
and U1924 (N_1924,N_927,N_1148);
and U1925 (N_1925,N_576,N_714);
nor U1926 (N_1926,N_469,N_1190);
or U1927 (N_1927,N_1225,N_535);
and U1928 (N_1928,N_1446,N_1316);
nor U1929 (N_1929,N_519,N_423);
or U1930 (N_1930,N_1475,N_1251);
or U1931 (N_1931,N_356,N_1072);
or U1932 (N_1932,N_1289,N_481);
and U1933 (N_1933,N_765,N_992);
xnor U1934 (N_1934,N_1231,N_1480);
nand U1935 (N_1935,N_999,N_770);
and U1936 (N_1936,N_685,N_577);
and U1937 (N_1937,N_945,N_136);
and U1938 (N_1938,N_1001,N_430);
or U1939 (N_1939,N_342,N_389);
and U1940 (N_1940,N_365,N_892);
or U1941 (N_1941,N_641,N_418);
nor U1942 (N_1942,N_1075,N_687);
nor U1943 (N_1943,N_1393,N_612);
nand U1944 (N_1944,N_1004,N_732);
nand U1945 (N_1945,N_657,N_871);
and U1946 (N_1946,N_1142,N_52);
nor U1947 (N_1947,N_893,N_166);
or U1948 (N_1948,N_589,N_327);
and U1949 (N_1949,N_384,N_1386);
and U1950 (N_1950,N_103,N_10);
xor U1951 (N_1951,N_619,N_1088);
nor U1952 (N_1952,N_150,N_1351);
xor U1953 (N_1953,N_834,N_911);
xnor U1954 (N_1954,N_584,N_724);
nor U1955 (N_1955,N_385,N_6);
or U1956 (N_1956,N_1076,N_1174);
nand U1957 (N_1957,N_1191,N_320);
xnor U1958 (N_1958,N_968,N_1262);
and U1959 (N_1959,N_279,N_1401);
xnor U1960 (N_1960,N_1182,N_1196);
nor U1961 (N_1961,N_1419,N_74);
and U1962 (N_1962,N_1291,N_1474);
xor U1963 (N_1963,N_457,N_681);
and U1964 (N_1964,N_363,N_895);
or U1965 (N_1965,N_562,N_1461);
xor U1966 (N_1966,N_1064,N_440);
or U1967 (N_1967,N_996,N_88);
xnor U1968 (N_1968,N_1337,N_1308);
nor U1969 (N_1969,N_769,N_1234);
nand U1970 (N_1970,N_491,N_957);
nor U1971 (N_1971,N_1471,N_439);
nor U1972 (N_1972,N_421,N_713);
nor U1973 (N_1973,N_762,N_349);
and U1974 (N_1974,N_1302,N_1044);
nor U1975 (N_1975,N_450,N_656);
or U1976 (N_1976,N_849,N_1416);
nand U1977 (N_1977,N_743,N_353);
nand U1978 (N_1978,N_444,N_1389);
xor U1979 (N_1979,N_162,N_1210);
nand U1980 (N_1980,N_1362,N_1421);
and U1981 (N_1981,N_817,N_302);
and U1982 (N_1982,N_115,N_209);
and U1983 (N_1983,N_1105,N_461);
nand U1984 (N_1984,N_717,N_818);
nand U1985 (N_1985,N_332,N_156);
or U1986 (N_1986,N_1178,N_1180);
and U1987 (N_1987,N_948,N_816);
xnor U1988 (N_1988,N_1242,N_454);
and U1989 (N_1989,N_1091,N_534);
nand U1990 (N_1990,N_410,N_1084);
or U1991 (N_1991,N_1010,N_1290);
nand U1992 (N_1992,N_105,N_699);
nand U1993 (N_1993,N_878,N_290);
nor U1994 (N_1994,N_373,N_987);
nand U1995 (N_1995,N_228,N_1029);
nand U1996 (N_1996,N_1256,N_725);
and U1997 (N_1997,N_531,N_870);
nand U1998 (N_1998,N_1279,N_492);
nand U1999 (N_1999,N_407,N_201);
or U2000 (N_2000,N_171,N_935);
and U2001 (N_2001,N_670,N_866);
xor U2002 (N_2002,N_1452,N_1278);
nor U2003 (N_2003,N_125,N_21);
nand U2004 (N_2004,N_375,N_843);
and U2005 (N_2005,N_1066,N_487);
or U2006 (N_2006,N_801,N_431);
nand U2007 (N_2007,N_564,N_886);
or U2008 (N_2008,N_941,N_554);
nand U2009 (N_2009,N_1428,N_984);
nand U2010 (N_2010,N_826,N_1403);
xnor U2011 (N_2011,N_1458,N_766);
or U2012 (N_2012,N_1039,N_1473);
and U2013 (N_2013,N_4,N_381);
nand U2014 (N_2014,N_881,N_1028);
and U2015 (N_2015,N_498,N_1405);
or U2016 (N_2016,N_163,N_420);
nor U2017 (N_2017,N_620,N_220);
nand U2018 (N_2018,N_309,N_1119);
nor U2019 (N_2019,N_419,N_703);
and U2020 (N_2020,N_931,N_1214);
and U2021 (N_2021,N_15,N_781);
and U2022 (N_2022,N_12,N_811);
xnor U2023 (N_2023,N_701,N_1324);
or U2024 (N_2024,N_594,N_981);
nand U2025 (N_2025,N_350,N_780);
and U2026 (N_2026,N_910,N_1043);
nor U2027 (N_2027,N_1204,N_106);
and U2028 (N_2028,N_231,N_1233);
or U2029 (N_2029,N_159,N_525);
nand U2030 (N_2030,N_661,N_428);
or U2031 (N_2031,N_1080,N_34);
or U2032 (N_2032,N_466,N_1126);
xnor U2033 (N_2033,N_192,N_284);
and U2034 (N_2034,N_376,N_1367);
xnor U2035 (N_2035,N_1434,N_1033);
nor U2036 (N_2036,N_1101,N_557);
nand U2037 (N_2037,N_684,N_443);
nor U2038 (N_2038,N_435,N_489);
or U2039 (N_2039,N_756,N_1395);
and U2040 (N_2040,N_260,N_139);
or U2041 (N_2041,N_194,N_449);
nand U2042 (N_2042,N_1073,N_17);
or U2043 (N_2043,N_414,N_92);
nand U2044 (N_2044,N_1443,N_606);
nand U2045 (N_2045,N_1152,N_1211);
xor U2046 (N_2046,N_1246,N_827);
or U2047 (N_2047,N_891,N_65);
xnor U2048 (N_2048,N_388,N_233);
xnor U2049 (N_2049,N_1472,N_7);
or U2050 (N_2050,N_537,N_1127);
or U2051 (N_2051,N_186,N_1476);
and U2052 (N_2052,N_1163,N_1378);
nor U2053 (N_2053,N_1413,N_245);
and U2054 (N_2054,N_512,N_998);
nor U2055 (N_2055,N_185,N_1267);
and U2056 (N_2056,N_977,N_963);
nor U2057 (N_2057,N_1430,N_1283);
nor U2058 (N_2058,N_257,N_678);
xnor U2059 (N_2059,N_1192,N_513);
nand U2060 (N_2060,N_1404,N_1162);
xnor U2061 (N_2061,N_427,N_347);
xor U2062 (N_2062,N_409,N_704);
or U2063 (N_2063,N_1195,N_143);
nand U2064 (N_2064,N_1150,N_123);
and U2065 (N_2065,N_1306,N_1482);
xnor U2066 (N_2066,N_160,N_971);
nand U2067 (N_2067,N_812,N_916);
xnor U2068 (N_2068,N_270,N_367);
or U2069 (N_2069,N_199,N_784);
xor U2070 (N_2070,N_1012,N_1425);
or U2071 (N_2071,N_1140,N_1269);
nor U2072 (N_2072,N_462,N_45);
xnor U2073 (N_2073,N_269,N_566);
nor U2074 (N_2074,N_1438,N_544);
nand U2075 (N_2075,N_464,N_1392);
nand U2076 (N_2076,N_565,N_1379);
xor U2077 (N_2077,N_36,N_28);
xor U2078 (N_2078,N_372,N_1123);
nand U2079 (N_2079,N_406,N_1207);
and U2080 (N_2080,N_96,N_806);
nand U2081 (N_2081,N_674,N_520);
and U2082 (N_2082,N_132,N_205);
xnor U2083 (N_2083,N_277,N_526);
xor U2084 (N_2084,N_1275,N_617);
xor U2085 (N_2085,N_72,N_672);
nor U2086 (N_2086,N_108,N_831);
or U2087 (N_2087,N_262,N_14);
or U2088 (N_2088,N_533,N_1498);
xor U2089 (N_2089,N_1354,N_1491);
xor U2090 (N_2090,N_335,N_354);
nand U2091 (N_2091,N_502,N_876);
xor U2092 (N_2092,N_786,N_991);
and U2093 (N_2093,N_336,N_973);
or U2094 (N_2094,N_133,N_1108);
or U2095 (N_2095,N_774,N_181);
nor U2096 (N_2096,N_823,N_296);
xnor U2097 (N_2097,N_436,N_197);
nor U2098 (N_2098,N_390,N_697);
xnor U2099 (N_2099,N_391,N_80);
nand U2100 (N_2100,N_588,N_1198);
nand U2101 (N_2101,N_1009,N_1023);
nand U2102 (N_2102,N_1206,N_794);
or U2103 (N_2103,N_305,N_691);
and U2104 (N_2104,N_196,N_671);
xnor U2105 (N_2105,N_458,N_453);
nor U2106 (N_2106,N_144,N_543);
or U2107 (N_2107,N_499,N_1470);
xnor U2108 (N_2108,N_804,N_468);
nand U2109 (N_2109,N_285,N_1402);
nor U2110 (N_2110,N_32,N_1113);
and U2111 (N_2111,N_1478,N_662);
nand U2112 (N_2112,N_579,N_89);
and U2113 (N_2113,N_802,N_1368);
xor U2114 (N_2114,N_967,N_18);
xor U2115 (N_2115,N_1496,N_1352);
or U2116 (N_2116,N_138,N_1005);
xor U2117 (N_2117,N_1063,N_955);
nor U2118 (N_2118,N_1353,N_1433);
nor U2119 (N_2119,N_938,N_608);
nor U2120 (N_2120,N_482,N_1447);
nand U2121 (N_2121,N_791,N_1332);
nor U2122 (N_2122,N_551,N_425);
nor U2123 (N_2123,N_708,N_676);
nor U2124 (N_2124,N_913,N_387);
or U2125 (N_2125,N_122,N_362);
nand U2126 (N_2126,N_914,N_345);
xor U2127 (N_2127,N_933,N_172);
or U2128 (N_2128,N_1002,N_1173);
or U2129 (N_2129,N_1410,N_1112);
nor U2130 (N_2130,N_865,N_653);
nand U2131 (N_2131,N_1311,N_1013);
and U2132 (N_2132,N_152,N_317);
nor U2133 (N_2133,N_1450,N_403);
and U2134 (N_2134,N_1213,N_1298);
xnor U2135 (N_2135,N_1299,N_374);
or U2136 (N_2136,N_787,N_137);
xor U2137 (N_2137,N_151,N_693);
nor U2138 (N_2138,N_1380,N_1006);
or U2139 (N_2139,N_294,N_1383);
nor U2140 (N_2140,N_969,N_982);
nor U2141 (N_2141,N_66,N_1061);
nand U2142 (N_2142,N_64,N_333);
nor U2143 (N_2143,N_569,N_600);
nor U2144 (N_2144,N_1116,N_1343);
or U2145 (N_2145,N_140,N_824);
xor U2146 (N_2146,N_154,N_1331);
nor U2147 (N_2147,N_613,N_885);
nand U2148 (N_2148,N_721,N_1215);
nor U2149 (N_2149,N_1477,N_1241);
or U2150 (N_2150,N_295,N_1261);
or U2151 (N_2151,N_546,N_187);
and U2152 (N_2152,N_616,N_164);
or U2153 (N_2153,N_621,N_472);
or U2154 (N_2154,N_1462,N_540);
nand U2155 (N_2155,N_255,N_1360);
nand U2156 (N_2156,N_995,N_877);
or U2157 (N_2157,N_1024,N_214);
xor U2158 (N_2158,N_1400,N_771);
nand U2159 (N_2159,N_1139,N_198);
or U2160 (N_2160,N_1448,N_779);
xnor U2161 (N_2161,N_632,N_1124);
nand U2162 (N_2162,N_282,N_1281);
nor U2163 (N_2163,N_68,N_855);
nand U2164 (N_2164,N_907,N_26);
xnor U2165 (N_2165,N_1411,N_924);
nor U2166 (N_2166,N_664,N_85);
nand U2167 (N_2167,N_1136,N_359);
and U2168 (N_2168,N_301,N_930);
or U2169 (N_2169,N_1328,N_596);
and U2170 (N_2170,N_860,N_142);
nand U2171 (N_2171,N_202,N_256);
or U2172 (N_2172,N_455,N_303);
xor U2173 (N_2173,N_1304,N_121);
xor U2174 (N_2174,N_441,N_1054);
and U2175 (N_2175,N_53,N_862);
and U2176 (N_2176,N_700,N_200);
nand U2177 (N_2177,N_300,N_1442);
xnor U2178 (N_2178,N_371,N_508);
and U2179 (N_2179,N_1305,N_1309);
nand U2180 (N_2180,N_234,N_1259);
or U2181 (N_2181,N_232,N_20);
or U2182 (N_2182,N_1226,N_1254);
or U2183 (N_2183,N_575,N_308);
nand U2184 (N_2184,N_1125,N_1321);
nor U2185 (N_2185,N_1377,N_1055);
nor U2186 (N_2186,N_903,N_404);
xor U2187 (N_2187,N_126,N_318);
nor U2188 (N_2188,N_683,N_230);
nand U2189 (N_2189,N_1260,N_650);
and U2190 (N_2190,N_715,N_299);
and U2191 (N_2191,N_104,N_1469);
nor U2192 (N_2192,N_243,N_675);
nand U2193 (N_2193,N_1107,N_965);
and U2194 (N_2194,N_1049,N_62);
nor U2195 (N_2195,N_516,N_326);
xor U2196 (N_2196,N_422,N_1031);
nand U2197 (N_2197,N_962,N_321);
xnor U2198 (N_2198,N_1052,N_858);
and U2199 (N_2199,N_548,N_586);
and U2200 (N_2200,N_399,N_1394);
nor U2201 (N_2201,N_1333,N_960);
nor U2202 (N_2202,N_180,N_486);
xor U2203 (N_2203,N_1432,N_1466);
nor U2204 (N_2204,N_837,N_702);
nand U2205 (N_2205,N_1270,N_553);
nand U2206 (N_2206,N_77,N_287);
nor U2207 (N_2207,N_433,N_1271);
nand U2208 (N_2208,N_393,N_1387);
nand U2209 (N_2209,N_91,N_1488);
nand U2210 (N_2210,N_394,N_1372);
and U2211 (N_2211,N_1027,N_47);
nand U2212 (N_2212,N_494,N_148);
or U2213 (N_2213,N_497,N_54);
nor U2214 (N_2214,N_1297,N_1218);
nor U2215 (N_2215,N_1201,N_764);
nor U2216 (N_2216,N_737,N_1327);
and U2217 (N_2217,N_709,N_400);
and U2218 (N_2218,N_275,N_238);
xnor U2219 (N_2219,N_111,N_506);
nand U2220 (N_2220,N_1396,N_863);
or U2221 (N_2221,N_563,N_840);
nand U2222 (N_2222,N_651,N_1048);
nand U2223 (N_2223,N_1183,N_459);
nor U2224 (N_2224,N_545,N_1122);
nor U2225 (N_2225,N_261,N_978);
or U2226 (N_2226,N_379,N_848);
and U2227 (N_2227,N_1371,N_97);
or U2228 (N_2228,N_341,N_835);
nor U2229 (N_2229,N_1245,N_1431);
xnor U2230 (N_2230,N_35,N_887);
nor U2231 (N_2231,N_915,N_1184);
and U2232 (N_2232,N_1227,N_1481);
nand U2233 (N_2233,N_1374,N_1455);
nor U2234 (N_2234,N_1286,N_798);
nor U2235 (N_2235,N_242,N_1022);
xor U2236 (N_2236,N_288,N_873);
xor U2237 (N_2237,N_838,N_868);
and U2238 (N_2238,N_883,N_51);
xnor U2239 (N_2239,N_782,N_1250);
or U2240 (N_2240,N_33,N_1095);
nand U2241 (N_2241,N_922,N_507);
or U2242 (N_2242,N_1158,N_549);
and U2243 (N_2243,N_1034,N_558);
nor U2244 (N_2244,N_845,N_247);
and U2245 (N_2245,N_9,N_644);
and U2246 (N_2246,N_1323,N_1382);
or U2247 (N_2247,N_470,N_1426);
nand U2248 (N_2248,N_383,N_1435);
and U2249 (N_2249,N_872,N_1272);
and U2250 (N_2250,N_482,N_1272);
nor U2251 (N_2251,N_762,N_638);
xor U2252 (N_2252,N_1356,N_394);
xnor U2253 (N_2253,N_1497,N_963);
nand U2254 (N_2254,N_873,N_86);
nand U2255 (N_2255,N_1299,N_79);
nor U2256 (N_2256,N_1349,N_923);
xnor U2257 (N_2257,N_1027,N_48);
nor U2258 (N_2258,N_1393,N_376);
xnor U2259 (N_2259,N_1371,N_1217);
nor U2260 (N_2260,N_1227,N_62);
nand U2261 (N_2261,N_1385,N_743);
and U2262 (N_2262,N_1205,N_458);
and U2263 (N_2263,N_786,N_493);
nor U2264 (N_2264,N_227,N_289);
xor U2265 (N_2265,N_456,N_478);
and U2266 (N_2266,N_1068,N_620);
xor U2267 (N_2267,N_1064,N_591);
or U2268 (N_2268,N_616,N_68);
or U2269 (N_2269,N_1048,N_1065);
and U2270 (N_2270,N_1493,N_1037);
nand U2271 (N_2271,N_880,N_1184);
and U2272 (N_2272,N_465,N_879);
or U2273 (N_2273,N_567,N_1381);
xnor U2274 (N_2274,N_237,N_1399);
or U2275 (N_2275,N_516,N_392);
nand U2276 (N_2276,N_158,N_629);
nor U2277 (N_2277,N_156,N_808);
or U2278 (N_2278,N_708,N_1101);
and U2279 (N_2279,N_166,N_926);
xor U2280 (N_2280,N_704,N_11);
nand U2281 (N_2281,N_432,N_1381);
xor U2282 (N_2282,N_50,N_916);
or U2283 (N_2283,N_1024,N_223);
nand U2284 (N_2284,N_369,N_629);
or U2285 (N_2285,N_1273,N_16);
or U2286 (N_2286,N_890,N_333);
nor U2287 (N_2287,N_958,N_68);
or U2288 (N_2288,N_1365,N_91);
or U2289 (N_2289,N_37,N_1402);
xnor U2290 (N_2290,N_284,N_368);
xor U2291 (N_2291,N_1398,N_186);
nand U2292 (N_2292,N_1390,N_1291);
or U2293 (N_2293,N_1468,N_541);
and U2294 (N_2294,N_247,N_1107);
xnor U2295 (N_2295,N_635,N_760);
nor U2296 (N_2296,N_583,N_688);
nand U2297 (N_2297,N_1002,N_101);
and U2298 (N_2298,N_950,N_669);
nor U2299 (N_2299,N_721,N_746);
nand U2300 (N_2300,N_1420,N_900);
or U2301 (N_2301,N_1252,N_754);
nand U2302 (N_2302,N_523,N_81);
or U2303 (N_2303,N_393,N_1044);
nor U2304 (N_2304,N_633,N_1112);
and U2305 (N_2305,N_1317,N_1187);
nand U2306 (N_2306,N_1122,N_380);
nor U2307 (N_2307,N_194,N_273);
or U2308 (N_2308,N_780,N_1266);
and U2309 (N_2309,N_938,N_1291);
or U2310 (N_2310,N_249,N_282);
xnor U2311 (N_2311,N_1370,N_116);
or U2312 (N_2312,N_564,N_1070);
nand U2313 (N_2313,N_1324,N_794);
nor U2314 (N_2314,N_1488,N_1011);
nand U2315 (N_2315,N_263,N_564);
nand U2316 (N_2316,N_930,N_176);
nand U2317 (N_2317,N_1195,N_779);
nand U2318 (N_2318,N_818,N_1334);
or U2319 (N_2319,N_1394,N_621);
and U2320 (N_2320,N_470,N_1240);
xnor U2321 (N_2321,N_411,N_1311);
xor U2322 (N_2322,N_420,N_1001);
nand U2323 (N_2323,N_386,N_466);
and U2324 (N_2324,N_1130,N_8);
xor U2325 (N_2325,N_1267,N_197);
nand U2326 (N_2326,N_612,N_249);
nand U2327 (N_2327,N_444,N_202);
nor U2328 (N_2328,N_1230,N_94);
or U2329 (N_2329,N_1375,N_155);
or U2330 (N_2330,N_77,N_391);
or U2331 (N_2331,N_382,N_955);
nand U2332 (N_2332,N_1089,N_320);
xnor U2333 (N_2333,N_1414,N_127);
or U2334 (N_2334,N_1197,N_938);
nor U2335 (N_2335,N_148,N_1183);
or U2336 (N_2336,N_1067,N_581);
xor U2337 (N_2337,N_1064,N_574);
nand U2338 (N_2338,N_626,N_156);
nor U2339 (N_2339,N_1312,N_144);
or U2340 (N_2340,N_551,N_1326);
nand U2341 (N_2341,N_148,N_1045);
and U2342 (N_2342,N_995,N_445);
nor U2343 (N_2343,N_478,N_178);
and U2344 (N_2344,N_511,N_594);
and U2345 (N_2345,N_893,N_499);
xor U2346 (N_2346,N_99,N_803);
xnor U2347 (N_2347,N_881,N_1489);
and U2348 (N_2348,N_452,N_1433);
or U2349 (N_2349,N_503,N_12);
and U2350 (N_2350,N_962,N_1320);
or U2351 (N_2351,N_785,N_912);
nor U2352 (N_2352,N_698,N_715);
nand U2353 (N_2353,N_1359,N_1425);
nand U2354 (N_2354,N_245,N_462);
and U2355 (N_2355,N_833,N_688);
nor U2356 (N_2356,N_1256,N_1300);
or U2357 (N_2357,N_1269,N_580);
or U2358 (N_2358,N_426,N_705);
or U2359 (N_2359,N_99,N_980);
or U2360 (N_2360,N_1439,N_85);
nor U2361 (N_2361,N_973,N_1499);
nor U2362 (N_2362,N_1292,N_1285);
nor U2363 (N_2363,N_108,N_85);
or U2364 (N_2364,N_76,N_569);
or U2365 (N_2365,N_194,N_1315);
or U2366 (N_2366,N_1485,N_774);
nor U2367 (N_2367,N_794,N_1218);
nor U2368 (N_2368,N_202,N_868);
and U2369 (N_2369,N_56,N_5);
nand U2370 (N_2370,N_1336,N_899);
xnor U2371 (N_2371,N_1066,N_1496);
or U2372 (N_2372,N_1472,N_806);
nand U2373 (N_2373,N_518,N_1275);
and U2374 (N_2374,N_355,N_990);
and U2375 (N_2375,N_650,N_950);
or U2376 (N_2376,N_1262,N_361);
xor U2377 (N_2377,N_70,N_1363);
nor U2378 (N_2378,N_782,N_545);
and U2379 (N_2379,N_1007,N_259);
and U2380 (N_2380,N_1422,N_976);
xnor U2381 (N_2381,N_1024,N_246);
and U2382 (N_2382,N_562,N_900);
xnor U2383 (N_2383,N_883,N_199);
or U2384 (N_2384,N_1170,N_778);
or U2385 (N_2385,N_1107,N_401);
or U2386 (N_2386,N_1155,N_979);
xnor U2387 (N_2387,N_485,N_685);
nand U2388 (N_2388,N_1144,N_680);
or U2389 (N_2389,N_416,N_835);
and U2390 (N_2390,N_681,N_949);
xor U2391 (N_2391,N_1149,N_960);
and U2392 (N_2392,N_1452,N_417);
nand U2393 (N_2393,N_458,N_1337);
nand U2394 (N_2394,N_608,N_1024);
nand U2395 (N_2395,N_181,N_820);
nor U2396 (N_2396,N_303,N_882);
nor U2397 (N_2397,N_1489,N_1154);
or U2398 (N_2398,N_1389,N_1027);
and U2399 (N_2399,N_404,N_989);
xor U2400 (N_2400,N_424,N_669);
or U2401 (N_2401,N_294,N_948);
and U2402 (N_2402,N_755,N_1049);
nor U2403 (N_2403,N_271,N_485);
nor U2404 (N_2404,N_1279,N_1010);
or U2405 (N_2405,N_1141,N_1435);
or U2406 (N_2406,N_1453,N_1297);
nor U2407 (N_2407,N_555,N_114);
or U2408 (N_2408,N_353,N_511);
or U2409 (N_2409,N_659,N_353);
nor U2410 (N_2410,N_867,N_1408);
nand U2411 (N_2411,N_768,N_899);
or U2412 (N_2412,N_1443,N_453);
or U2413 (N_2413,N_1007,N_1440);
and U2414 (N_2414,N_151,N_965);
or U2415 (N_2415,N_1377,N_922);
xor U2416 (N_2416,N_68,N_219);
xor U2417 (N_2417,N_1394,N_276);
nor U2418 (N_2418,N_518,N_1252);
or U2419 (N_2419,N_1246,N_1264);
nand U2420 (N_2420,N_607,N_1254);
nand U2421 (N_2421,N_873,N_1204);
xnor U2422 (N_2422,N_260,N_545);
and U2423 (N_2423,N_833,N_592);
and U2424 (N_2424,N_1215,N_130);
and U2425 (N_2425,N_79,N_1065);
or U2426 (N_2426,N_769,N_558);
xnor U2427 (N_2427,N_1205,N_537);
nand U2428 (N_2428,N_1196,N_1160);
and U2429 (N_2429,N_915,N_32);
or U2430 (N_2430,N_160,N_896);
and U2431 (N_2431,N_706,N_594);
and U2432 (N_2432,N_667,N_517);
nor U2433 (N_2433,N_112,N_993);
nand U2434 (N_2434,N_819,N_1051);
xnor U2435 (N_2435,N_880,N_762);
and U2436 (N_2436,N_832,N_81);
or U2437 (N_2437,N_1472,N_1146);
and U2438 (N_2438,N_397,N_1022);
nor U2439 (N_2439,N_489,N_707);
or U2440 (N_2440,N_714,N_546);
and U2441 (N_2441,N_217,N_590);
and U2442 (N_2442,N_994,N_353);
and U2443 (N_2443,N_6,N_565);
or U2444 (N_2444,N_475,N_9);
or U2445 (N_2445,N_170,N_204);
nand U2446 (N_2446,N_388,N_1122);
nor U2447 (N_2447,N_906,N_1318);
or U2448 (N_2448,N_1334,N_691);
xor U2449 (N_2449,N_1196,N_743);
and U2450 (N_2450,N_943,N_622);
nor U2451 (N_2451,N_1171,N_927);
or U2452 (N_2452,N_38,N_622);
nand U2453 (N_2453,N_415,N_480);
nand U2454 (N_2454,N_1130,N_60);
and U2455 (N_2455,N_1162,N_1378);
xnor U2456 (N_2456,N_356,N_345);
and U2457 (N_2457,N_516,N_47);
or U2458 (N_2458,N_228,N_1426);
or U2459 (N_2459,N_387,N_1142);
xnor U2460 (N_2460,N_716,N_967);
nand U2461 (N_2461,N_371,N_91);
xor U2462 (N_2462,N_767,N_1445);
nor U2463 (N_2463,N_1367,N_408);
xor U2464 (N_2464,N_677,N_282);
nand U2465 (N_2465,N_741,N_538);
and U2466 (N_2466,N_363,N_1318);
and U2467 (N_2467,N_978,N_1410);
nand U2468 (N_2468,N_1258,N_923);
xor U2469 (N_2469,N_468,N_467);
xnor U2470 (N_2470,N_1263,N_958);
nand U2471 (N_2471,N_1118,N_136);
nand U2472 (N_2472,N_79,N_435);
and U2473 (N_2473,N_786,N_1182);
and U2474 (N_2474,N_74,N_248);
xnor U2475 (N_2475,N_1059,N_202);
nand U2476 (N_2476,N_559,N_1006);
nor U2477 (N_2477,N_1146,N_106);
xor U2478 (N_2478,N_739,N_30);
and U2479 (N_2479,N_700,N_696);
or U2480 (N_2480,N_14,N_1198);
and U2481 (N_2481,N_1136,N_873);
and U2482 (N_2482,N_199,N_1286);
xor U2483 (N_2483,N_285,N_518);
nand U2484 (N_2484,N_726,N_528);
and U2485 (N_2485,N_453,N_1044);
or U2486 (N_2486,N_508,N_1480);
nor U2487 (N_2487,N_784,N_197);
nor U2488 (N_2488,N_278,N_651);
nor U2489 (N_2489,N_688,N_69);
nor U2490 (N_2490,N_815,N_1090);
xnor U2491 (N_2491,N_882,N_264);
xor U2492 (N_2492,N_600,N_1456);
xnor U2493 (N_2493,N_1365,N_220);
and U2494 (N_2494,N_1169,N_310);
and U2495 (N_2495,N_475,N_1418);
xor U2496 (N_2496,N_362,N_1271);
xnor U2497 (N_2497,N_538,N_1449);
xor U2498 (N_2498,N_1131,N_481);
nor U2499 (N_2499,N_833,N_546);
nand U2500 (N_2500,N_1155,N_1122);
nor U2501 (N_2501,N_1310,N_850);
or U2502 (N_2502,N_338,N_781);
xnor U2503 (N_2503,N_766,N_116);
or U2504 (N_2504,N_740,N_253);
nand U2505 (N_2505,N_859,N_996);
and U2506 (N_2506,N_851,N_1008);
xor U2507 (N_2507,N_1148,N_1190);
nor U2508 (N_2508,N_295,N_956);
and U2509 (N_2509,N_287,N_394);
nand U2510 (N_2510,N_976,N_317);
or U2511 (N_2511,N_575,N_73);
xor U2512 (N_2512,N_1432,N_1084);
and U2513 (N_2513,N_149,N_575);
or U2514 (N_2514,N_165,N_655);
xor U2515 (N_2515,N_977,N_1350);
xnor U2516 (N_2516,N_708,N_707);
nor U2517 (N_2517,N_251,N_1392);
nor U2518 (N_2518,N_1484,N_455);
nand U2519 (N_2519,N_55,N_487);
and U2520 (N_2520,N_1077,N_722);
xnor U2521 (N_2521,N_1286,N_551);
and U2522 (N_2522,N_347,N_513);
nor U2523 (N_2523,N_921,N_990);
xor U2524 (N_2524,N_581,N_1378);
nor U2525 (N_2525,N_1498,N_345);
nand U2526 (N_2526,N_870,N_410);
and U2527 (N_2527,N_856,N_575);
xnor U2528 (N_2528,N_1139,N_182);
nand U2529 (N_2529,N_983,N_534);
and U2530 (N_2530,N_429,N_574);
or U2531 (N_2531,N_731,N_783);
or U2532 (N_2532,N_726,N_1164);
nor U2533 (N_2533,N_854,N_1112);
or U2534 (N_2534,N_628,N_737);
xor U2535 (N_2535,N_937,N_1322);
nand U2536 (N_2536,N_729,N_490);
nor U2537 (N_2537,N_1422,N_23);
and U2538 (N_2538,N_1114,N_969);
or U2539 (N_2539,N_690,N_637);
xor U2540 (N_2540,N_789,N_412);
nor U2541 (N_2541,N_437,N_541);
and U2542 (N_2542,N_1194,N_504);
and U2543 (N_2543,N_1204,N_1488);
nor U2544 (N_2544,N_1476,N_175);
xor U2545 (N_2545,N_475,N_406);
or U2546 (N_2546,N_1312,N_760);
nand U2547 (N_2547,N_1212,N_423);
or U2548 (N_2548,N_1402,N_1114);
nand U2549 (N_2549,N_299,N_125);
xnor U2550 (N_2550,N_678,N_888);
nand U2551 (N_2551,N_1448,N_502);
and U2552 (N_2552,N_725,N_515);
nand U2553 (N_2553,N_694,N_980);
and U2554 (N_2554,N_25,N_264);
nor U2555 (N_2555,N_805,N_1353);
or U2556 (N_2556,N_1021,N_642);
nand U2557 (N_2557,N_581,N_1397);
nand U2558 (N_2558,N_1235,N_1304);
nand U2559 (N_2559,N_213,N_701);
xnor U2560 (N_2560,N_428,N_1262);
or U2561 (N_2561,N_1064,N_479);
or U2562 (N_2562,N_678,N_663);
and U2563 (N_2563,N_1326,N_833);
or U2564 (N_2564,N_340,N_329);
or U2565 (N_2565,N_1478,N_1214);
nor U2566 (N_2566,N_485,N_1084);
or U2567 (N_2567,N_983,N_334);
or U2568 (N_2568,N_1178,N_1383);
nand U2569 (N_2569,N_472,N_1144);
or U2570 (N_2570,N_1072,N_922);
nor U2571 (N_2571,N_1075,N_198);
nor U2572 (N_2572,N_205,N_150);
nor U2573 (N_2573,N_737,N_859);
nor U2574 (N_2574,N_1218,N_1404);
or U2575 (N_2575,N_907,N_53);
xor U2576 (N_2576,N_248,N_1219);
nor U2577 (N_2577,N_230,N_1175);
and U2578 (N_2578,N_696,N_502);
xor U2579 (N_2579,N_274,N_840);
xor U2580 (N_2580,N_253,N_68);
and U2581 (N_2581,N_593,N_1343);
and U2582 (N_2582,N_1004,N_765);
and U2583 (N_2583,N_343,N_1357);
nor U2584 (N_2584,N_511,N_479);
or U2585 (N_2585,N_524,N_1420);
xor U2586 (N_2586,N_1210,N_55);
xnor U2587 (N_2587,N_885,N_1149);
nor U2588 (N_2588,N_1269,N_590);
or U2589 (N_2589,N_1369,N_1012);
nor U2590 (N_2590,N_697,N_1307);
nand U2591 (N_2591,N_705,N_1000);
nor U2592 (N_2592,N_333,N_1465);
xnor U2593 (N_2593,N_1264,N_1275);
or U2594 (N_2594,N_886,N_1013);
and U2595 (N_2595,N_1203,N_109);
nor U2596 (N_2596,N_452,N_1430);
nor U2597 (N_2597,N_293,N_972);
xnor U2598 (N_2598,N_1274,N_869);
xor U2599 (N_2599,N_1241,N_1174);
and U2600 (N_2600,N_1130,N_662);
nor U2601 (N_2601,N_683,N_1011);
xor U2602 (N_2602,N_956,N_462);
or U2603 (N_2603,N_935,N_238);
xor U2604 (N_2604,N_1303,N_817);
nand U2605 (N_2605,N_1258,N_517);
and U2606 (N_2606,N_941,N_687);
or U2607 (N_2607,N_1374,N_613);
or U2608 (N_2608,N_1418,N_457);
xor U2609 (N_2609,N_992,N_1426);
or U2610 (N_2610,N_663,N_341);
xnor U2611 (N_2611,N_1033,N_1144);
and U2612 (N_2612,N_912,N_328);
and U2613 (N_2613,N_942,N_535);
and U2614 (N_2614,N_508,N_888);
and U2615 (N_2615,N_282,N_534);
or U2616 (N_2616,N_341,N_815);
xor U2617 (N_2617,N_612,N_1129);
nor U2618 (N_2618,N_600,N_1377);
or U2619 (N_2619,N_1399,N_1283);
or U2620 (N_2620,N_782,N_485);
nand U2621 (N_2621,N_224,N_40);
or U2622 (N_2622,N_1342,N_809);
and U2623 (N_2623,N_1350,N_873);
nor U2624 (N_2624,N_1457,N_1490);
nand U2625 (N_2625,N_752,N_1269);
or U2626 (N_2626,N_616,N_1195);
or U2627 (N_2627,N_361,N_281);
nand U2628 (N_2628,N_345,N_1295);
nand U2629 (N_2629,N_253,N_1451);
and U2630 (N_2630,N_911,N_856);
nand U2631 (N_2631,N_1215,N_243);
and U2632 (N_2632,N_219,N_577);
or U2633 (N_2633,N_17,N_1197);
nor U2634 (N_2634,N_926,N_815);
or U2635 (N_2635,N_1378,N_761);
or U2636 (N_2636,N_1404,N_1325);
nand U2637 (N_2637,N_416,N_868);
nor U2638 (N_2638,N_1003,N_59);
xnor U2639 (N_2639,N_965,N_330);
or U2640 (N_2640,N_1186,N_944);
nand U2641 (N_2641,N_1137,N_42);
nor U2642 (N_2642,N_639,N_1289);
and U2643 (N_2643,N_1260,N_728);
nor U2644 (N_2644,N_902,N_542);
and U2645 (N_2645,N_894,N_500);
nand U2646 (N_2646,N_1396,N_1192);
and U2647 (N_2647,N_256,N_548);
nand U2648 (N_2648,N_646,N_811);
nand U2649 (N_2649,N_10,N_398);
nor U2650 (N_2650,N_199,N_533);
xnor U2651 (N_2651,N_1401,N_1114);
and U2652 (N_2652,N_605,N_1474);
nand U2653 (N_2653,N_938,N_1069);
xnor U2654 (N_2654,N_1312,N_1158);
xnor U2655 (N_2655,N_1195,N_367);
or U2656 (N_2656,N_18,N_1203);
xnor U2657 (N_2657,N_436,N_1198);
xor U2658 (N_2658,N_1351,N_164);
or U2659 (N_2659,N_282,N_1268);
xnor U2660 (N_2660,N_746,N_502);
xnor U2661 (N_2661,N_949,N_1397);
nand U2662 (N_2662,N_68,N_249);
xnor U2663 (N_2663,N_982,N_1256);
xnor U2664 (N_2664,N_1250,N_1061);
and U2665 (N_2665,N_607,N_679);
nor U2666 (N_2666,N_1163,N_236);
xnor U2667 (N_2667,N_862,N_367);
nor U2668 (N_2668,N_1266,N_1087);
and U2669 (N_2669,N_428,N_1331);
and U2670 (N_2670,N_463,N_626);
and U2671 (N_2671,N_4,N_580);
and U2672 (N_2672,N_220,N_639);
or U2673 (N_2673,N_1407,N_1085);
nand U2674 (N_2674,N_267,N_303);
nor U2675 (N_2675,N_974,N_627);
nor U2676 (N_2676,N_666,N_1029);
and U2677 (N_2677,N_94,N_416);
or U2678 (N_2678,N_1165,N_1103);
xor U2679 (N_2679,N_140,N_662);
or U2680 (N_2680,N_1349,N_782);
nand U2681 (N_2681,N_639,N_76);
and U2682 (N_2682,N_480,N_111);
nand U2683 (N_2683,N_748,N_81);
xor U2684 (N_2684,N_775,N_1035);
nand U2685 (N_2685,N_76,N_783);
nor U2686 (N_2686,N_392,N_538);
and U2687 (N_2687,N_878,N_289);
or U2688 (N_2688,N_182,N_721);
or U2689 (N_2689,N_675,N_237);
xor U2690 (N_2690,N_1092,N_15);
xor U2691 (N_2691,N_1374,N_1180);
or U2692 (N_2692,N_487,N_1476);
and U2693 (N_2693,N_929,N_1453);
xnor U2694 (N_2694,N_1220,N_315);
or U2695 (N_2695,N_1316,N_389);
or U2696 (N_2696,N_1047,N_932);
xor U2697 (N_2697,N_1468,N_308);
xor U2698 (N_2698,N_1377,N_743);
or U2699 (N_2699,N_1075,N_1016);
nand U2700 (N_2700,N_492,N_188);
and U2701 (N_2701,N_338,N_1211);
or U2702 (N_2702,N_73,N_691);
and U2703 (N_2703,N_189,N_178);
nor U2704 (N_2704,N_339,N_636);
nor U2705 (N_2705,N_1465,N_436);
nor U2706 (N_2706,N_1436,N_1198);
nand U2707 (N_2707,N_204,N_1194);
nor U2708 (N_2708,N_331,N_409);
or U2709 (N_2709,N_339,N_646);
nand U2710 (N_2710,N_1219,N_701);
or U2711 (N_2711,N_861,N_1150);
and U2712 (N_2712,N_581,N_265);
and U2713 (N_2713,N_1194,N_1069);
and U2714 (N_2714,N_501,N_163);
xor U2715 (N_2715,N_144,N_50);
xor U2716 (N_2716,N_142,N_392);
and U2717 (N_2717,N_1412,N_1183);
nor U2718 (N_2718,N_1389,N_24);
xor U2719 (N_2719,N_150,N_1139);
or U2720 (N_2720,N_192,N_543);
xnor U2721 (N_2721,N_100,N_1243);
xnor U2722 (N_2722,N_616,N_1315);
xnor U2723 (N_2723,N_157,N_955);
xor U2724 (N_2724,N_165,N_876);
nor U2725 (N_2725,N_1418,N_168);
or U2726 (N_2726,N_547,N_22);
and U2727 (N_2727,N_344,N_340);
and U2728 (N_2728,N_1279,N_1403);
xnor U2729 (N_2729,N_122,N_1040);
xor U2730 (N_2730,N_57,N_319);
or U2731 (N_2731,N_77,N_1020);
and U2732 (N_2732,N_1150,N_924);
and U2733 (N_2733,N_142,N_1447);
nand U2734 (N_2734,N_843,N_1076);
nand U2735 (N_2735,N_240,N_1430);
or U2736 (N_2736,N_633,N_641);
nand U2737 (N_2737,N_186,N_752);
or U2738 (N_2738,N_838,N_292);
xnor U2739 (N_2739,N_498,N_206);
xor U2740 (N_2740,N_987,N_208);
and U2741 (N_2741,N_803,N_805);
nand U2742 (N_2742,N_1304,N_1362);
and U2743 (N_2743,N_100,N_959);
and U2744 (N_2744,N_210,N_1498);
nor U2745 (N_2745,N_1125,N_381);
or U2746 (N_2746,N_162,N_1499);
xor U2747 (N_2747,N_329,N_228);
nor U2748 (N_2748,N_26,N_403);
nor U2749 (N_2749,N_441,N_538);
and U2750 (N_2750,N_1072,N_1185);
xnor U2751 (N_2751,N_1328,N_503);
nand U2752 (N_2752,N_1124,N_576);
nor U2753 (N_2753,N_665,N_1427);
xor U2754 (N_2754,N_85,N_700);
xnor U2755 (N_2755,N_1297,N_1229);
or U2756 (N_2756,N_462,N_1243);
nand U2757 (N_2757,N_729,N_1281);
nor U2758 (N_2758,N_774,N_1407);
nand U2759 (N_2759,N_451,N_244);
nand U2760 (N_2760,N_921,N_945);
nand U2761 (N_2761,N_1435,N_172);
nand U2762 (N_2762,N_1496,N_676);
nand U2763 (N_2763,N_964,N_1042);
or U2764 (N_2764,N_1358,N_52);
or U2765 (N_2765,N_422,N_1213);
nand U2766 (N_2766,N_761,N_774);
nor U2767 (N_2767,N_1408,N_146);
or U2768 (N_2768,N_683,N_59);
and U2769 (N_2769,N_334,N_1154);
xnor U2770 (N_2770,N_929,N_537);
and U2771 (N_2771,N_306,N_1139);
or U2772 (N_2772,N_75,N_825);
nor U2773 (N_2773,N_744,N_351);
xor U2774 (N_2774,N_711,N_1358);
xnor U2775 (N_2775,N_573,N_148);
nor U2776 (N_2776,N_285,N_1195);
nand U2777 (N_2777,N_1242,N_713);
xnor U2778 (N_2778,N_990,N_1421);
xor U2779 (N_2779,N_696,N_398);
xnor U2780 (N_2780,N_272,N_865);
or U2781 (N_2781,N_1291,N_339);
or U2782 (N_2782,N_320,N_1373);
or U2783 (N_2783,N_595,N_1420);
xnor U2784 (N_2784,N_457,N_1295);
xor U2785 (N_2785,N_267,N_1407);
nand U2786 (N_2786,N_36,N_32);
nor U2787 (N_2787,N_541,N_243);
nor U2788 (N_2788,N_568,N_1114);
nor U2789 (N_2789,N_1284,N_1420);
xor U2790 (N_2790,N_1493,N_1128);
or U2791 (N_2791,N_98,N_791);
nand U2792 (N_2792,N_1315,N_226);
or U2793 (N_2793,N_933,N_1347);
or U2794 (N_2794,N_1474,N_582);
and U2795 (N_2795,N_717,N_439);
or U2796 (N_2796,N_443,N_1464);
and U2797 (N_2797,N_289,N_1034);
and U2798 (N_2798,N_651,N_1484);
and U2799 (N_2799,N_353,N_708);
nor U2800 (N_2800,N_931,N_34);
nor U2801 (N_2801,N_1308,N_380);
nor U2802 (N_2802,N_1343,N_399);
and U2803 (N_2803,N_264,N_537);
xor U2804 (N_2804,N_1244,N_360);
nor U2805 (N_2805,N_1460,N_1058);
and U2806 (N_2806,N_1452,N_1260);
and U2807 (N_2807,N_1031,N_798);
nand U2808 (N_2808,N_1308,N_459);
nor U2809 (N_2809,N_1218,N_981);
xor U2810 (N_2810,N_1300,N_600);
xnor U2811 (N_2811,N_458,N_861);
or U2812 (N_2812,N_361,N_637);
or U2813 (N_2813,N_504,N_1202);
nor U2814 (N_2814,N_1311,N_1069);
or U2815 (N_2815,N_823,N_534);
xnor U2816 (N_2816,N_1129,N_472);
or U2817 (N_2817,N_255,N_1177);
nand U2818 (N_2818,N_1436,N_849);
and U2819 (N_2819,N_1482,N_947);
xnor U2820 (N_2820,N_1246,N_1323);
and U2821 (N_2821,N_439,N_919);
and U2822 (N_2822,N_772,N_1038);
or U2823 (N_2823,N_1143,N_540);
nand U2824 (N_2824,N_114,N_794);
nor U2825 (N_2825,N_171,N_439);
nor U2826 (N_2826,N_1343,N_241);
nor U2827 (N_2827,N_514,N_1070);
or U2828 (N_2828,N_641,N_1444);
and U2829 (N_2829,N_708,N_100);
nor U2830 (N_2830,N_463,N_776);
or U2831 (N_2831,N_73,N_1444);
and U2832 (N_2832,N_763,N_1477);
or U2833 (N_2833,N_497,N_223);
and U2834 (N_2834,N_716,N_1144);
xor U2835 (N_2835,N_468,N_793);
nand U2836 (N_2836,N_1473,N_1144);
and U2837 (N_2837,N_379,N_254);
nor U2838 (N_2838,N_1311,N_147);
nand U2839 (N_2839,N_35,N_382);
nor U2840 (N_2840,N_730,N_608);
or U2841 (N_2841,N_29,N_407);
and U2842 (N_2842,N_1271,N_1462);
nor U2843 (N_2843,N_517,N_894);
nand U2844 (N_2844,N_1218,N_267);
or U2845 (N_2845,N_654,N_386);
nand U2846 (N_2846,N_1185,N_857);
or U2847 (N_2847,N_1469,N_1238);
or U2848 (N_2848,N_1190,N_147);
nand U2849 (N_2849,N_1445,N_1003);
nor U2850 (N_2850,N_1242,N_838);
nor U2851 (N_2851,N_674,N_679);
and U2852 (N_2852,N_595,N_13);
nand U2853 (N_2853,N_1125,N_4);
nor U2854 (N_2854,N_649,N_22);
and U2855 (N_2855,N_1065,N_207);
and U2856 (N_2856,N_138,N_882);
nor U2857 (N_2857,N_1097,N_1117);
or U2858 (N_2858,N_634,N_1247);
nand U2859 (N_2859,N_187,N_145);
xor U2860 (N_2860,N_929,N_408);
nor U2861 (N_2861,N_57,N_293);
and U2862 (N_2862,N_1272,N_107);
and U2863 (N_2863,N_972,N_1285);
and U2864 (N_2864,N_942,N_1005);
nor U2865 (N_2865,N_798,N_187);
nand U2866 (N_2866,N_1229,N_1331);
and U2867 (N_2867,N_1333,N_561);
xor U2868 (N_2868,N_1124,N_1492);
or U2869 (N_2869,N_1033,N_1363);
nor U2870 (N_2870,N_1215,N_1387);
xor U2871 (N_2871,N_709,N_396);
xor U2872 (N_2872,N_1428,N_1134);
nor U2873 (N_2873,N_1312,N_789);
nand U2874 (N_2874,N_651,N_254);
and U2875 (N_2875,N_346,N_1116);
nand U2876 (N_2876,N_1415,N_1454);
and U2877 (N_2877,N_146,N_1167);
nand U2878 (N_2878,N_954,N_1048);
xnor U2879 (N_2879,N_486,N_390);
xor U2880 (N_2880,N_826,N_1226);
nand U2881 (N_2881,N_114,N_495);
nand U2882 (N_2882,N_1247,N_898);
nand U2883 (N_2883,N_493,N_403);
nor U2884 (N_2884,N_467,N_412);
nor U2885 (N_2885,N_0,N_1051);
or U2886 (N_2886,N_1051,N_931);
nor U2887 (N_2887,N_628,N_471);
nor U2888 (N_2888,N_874,N_24);
xnor U2889 (N_2889,N_1030,N_494);
xnor U2890 (N_2890,N_836,N_124);
and U2891 (N_2891,N_74,N_1193);
or U2892 (N_2892,N_349,N_316);
or U2893 (N_2893,N_702,N_532);
xor U2894 (N_2894,N_680,N_1185);
nor U2895 (N_2895,N_528,N_1043);
nand U2896 (N_2896,N_37,N_1439);
nor U2897 (N_2897,N_393,N_256);
nor U2898 (N_2898,N_69,N_1079);
or U2899 (N_2899,N_1012,N_1427);
xor U2900 (N_2900,N_1386,N_1413);
and U2901 (N_2901,N_402,N_1215);
nand U2902 (N_2902,N_463,N_1159);
and U2903 (N_2903,N_1302,N_1146);
or U2904 (N_2904,N_1120,N_235);
or U2905 (N_2905,N_567,N_534);
and U2906 (N_2906,N_1254,N_506);
nand U2907 (N_2907,N_904,N_817);
or U2908 (N_2908,N_32,N_880);
and U2909 (N_2909,N_562,N_887);
and U2910 (N_2910,N_372,N_1343);
or U2911 (N_2911,N_500,N_646);
and U2912 (N_2912,N_92,N_1027);
and U2913 (N_2913,N_340,N_783);
or U2914 (N_2914,N_1449,N_1367);
nand U2915 (N_2915,N_1060,N_406);
xnor U2916 (N_2916,N_741,N_602);
xnor U2917 (N_2917,N_782,N_281);
or U2918 (N_2918,N_241,N_964);
nand U2919 (N_2919,N_26,N_259);
nor U2920 (N_2920,N_1440,N_785);
and U2921 (N_2921,N_319,N_1051);
and U2922 (N_2922,N_121,N_309);
nand U2923 (N_2923,N_1087,N_302);
xor U2924 (N_2924,N_459,N_1081);
and U2925 (N_2925,N_615,N_486);
or U2926 (N_2926,N_132,N_520);
or U2927 (N_2927,N_444,N_691);
xor U2928 (N_2928,N_345,N_381);
xor U2929 (N_2929,N_23,N_172);
and U2930 (N_2930,N_355,N_224);
nand U2931 (N_2931,N_587,N_496);
and U2932 (N_2932,N_1448,N_852);
or U2933 (N_2933,N_330,N_1306);
nor U2934 (N_2934,N_304,N_638);
nand U2935 (N_2935,N_695,N_1096);
xor U2936 (N_2936,N_1165,N_1420);
or U2937 (N_2937,N_78,N_899);
and U2938 (N_2938,N_26,N_1126);
nor U2939 (N_2939,N_885,N_104);
nand U2940 (N_2940,N_791,N_132);
nor U2941 (N_2941,N_795,N_1096);
nor U2942 (N_2942,N_959,N_39);
xor U2943 (N_2943,N_1330,N_22);
nor U2944 (N_2944,N_102,N_367);
or U2945 (N_2945,N_702,N_529);
nand U2946 (N_2946,N_1418,N_1277);
or U2947 (N_2947,N_690,N_687);
xnor U2948 (N_2948,N_757,N_926);
nor U2949 (N_2949,N_778,N_799);
and U2950 (N_2950,N_615,N_1376);
nor U2951 (N_2951,N_647,N_412);
xor U2952 (N_2952,N_1050,N_1080);
or U2953 (N_2953,N_1476,N_695);
nand U2954 (N_2954,N_152,N_1023);
or U2955 (N_2955,N_1248,N_1157);
or U2956 (N_2956,N_1363,N_801);
or U2957 (N_2957,N_261,N_473);
or U2958 (N_2958,N_559,N_673);
or U2959 (N_2959,N_704,N_908);
xor U2960 (N_2960,N_536,N_39);
nand U2961 (N_2961,N_733,N_65);
nand U2962 (N_2962,N_838,N_1065);
and U2963 (N_2963,N_217,N_989);
nor U2964 (N_2964,N_490,N_1318);
nand U2965 (N_2965,N_834,N_320);
or U2966 (N_2966,N_828,N_1425);
nand U2967 (N_2967,N_521,N_1194);
xnor U2968 (N_2968,N_100,N_1031);
nand U2969 (N_2969,N_651,N_257);
and U2970 (N_2970,N_223,N_544);
xnor U2971 (N_2971,N_933,N_580);
and U2972 (N_2972,N_234,N_287);
nor U2973 (N_2973,N_1091,N_434);
nand U2974 (N_2974,N_328,N_1225);
nand U2975 (N_2975,N_529,N_304);
and U2976 (N_2976,N_1421,N_407);
or U2977 (N_2977,N_1338,N_871);
or U2978 (N_2978,N_85,N_401);
xnor U2979 (N_2979,N_169,N_633);
and U2980 (N_2980,N_978,N_1394);
nand U2981 (N_2981,N_52,N_1092);
or U2982 (N_2982,N_1163,N_335);
xor U2983 (N_2983,N_884,N_1169);
nand U2984 (N_2984,N_693,N_86);
or U2985 (N_2985,N_437,N_629);
xnor U2986 (N_2986,N_481,N_145);
nor U2987 (N_2987,N_136,N_243);
nor U2988 (N_2988,N_478,N_1100);
xnor U2989 (N_2989,N_997,N_641);
xnor U2990 (N_2990,N_1295,N_1001);
or U2991 (N_2991,N_883,N_1373);
nand U2992 (N_2992,N_232,N_554);
nand U2993 (N_2993,N_270,N_434);
and U2994 (N_2994,N_781,N_1390);
or U2995 (N_2995,N_1012,N_117);
nor U2996 (N_2996,N_1320,N_463);
and U2997 (N_2997,N_219,N_1095);
and U2998 (N_2998,N_1248,N_467);
xor U2999 (N_2999,N_497,N_807);
nor U3000 (N_3000,N_2958,N_2390);
or U3001 (N_3001,N_1911,N_1550);
or U3002 (N_3002,N_1761,N_2242);
or U3003 (N_3003,N_2712,N_2266);
nor U3004 (N_3004,N_2702,N_2497);
xnor U3005 (N_3005,N_2288,N_2001);
nor U3006 (N_3006,N_2844,N_2180);
nor U3007 (N_3007,N_2463,N_2585);
or U3008 (N_3008,N_1693,N_2281);
and U3009 (N_3009,N_2686,N_2224);
nor U3010 (N_3010,N_2655,N_1873);
and U3011 (N_3011,N_2944,N_2229);
nand U3012 (N_3012,N_2809,N_2941);
nand U3013 (N_3013,N_2684,N_1616);
xnor U3014 (N_3014,N_2709,N_2588);
and U3015 (N_3015,N_2311,N_1851);
nor U3016 (N_3016,N_1917,N_2552);
nor U3017 (N_3017,N_2237,N_2946);
nor U3018 (N_3018,N_1714,N_2459);
and U3019 (N_3019,N_2728,N_2255);
nand U3020 (N_3020,N_2559,N_2782);
nor U3021 (N_3021,N_1884,N_2524);
or U3022 (N_3022,N_1559,N_2408);
and U3023 (N_3023,N_1619,N_2598);
xnor U3024 (N_3024,N_2439,N_1674);
and U3025 (N_3025,N_1590,N_2584);
or U3026 (N_3026,N_2006,N_1500);
xnor U3027 (N_3027,N_2149,N_2577);
and U3028 (N_3028,N_2232,N_2564);
or U3029 (N_3029,N_2558,N_1875);
and U3030 (N_3030,N_2556,N_1644);
xnor U3031 (N_3031,N_2231,N_2307);
and U3032 (N_3032,N_2545,N_2005);
nand U3033 (N_3033,N_1752,N_2828);
nor U3034 (N_3034,N_2124,N_1855);
or U3035 (N_3035,N_2355,N_2392);
or U3036 (N_3036,N_2056,N_1871);
xor U3037 (N_3037,N_2450,N_2472);
and U3038 (N_3038,N_2157,N_1886);
xor U3039 (N_3039,N_1642,N_2485);
nor U3040 (N_3040,N_1692,N_1667);
or U3041 (N_3041,N_1518,N_2331);
xnor U3042 (N_3042,N_1777,N_2103);
or U3043 (N_3043,N_2050,N_2030);
xnor U3044 (N_3044,N_2747,N_2064);
nor U3045 (N_3045,N_1632,N_2053);
nor U3046 (N_3046,N_2205,N_1792);
xnor U3047 (N_3047,N_2025,N_1996);
nor U3048 (N_3048,N_2634,N_2457);
or U3049 (N_3049,N_1919,N_2183);
nor U3050 (N_3050,N_2735,N_1574);
xor U3051 (N_3051,N_1625,N_2429);
xnor U3052 (N_3052,N_2706,N_2017);
and U3053 (N_3053,N_2928,N_2913);
nor U3054 (N_3054,N_1925,N_1572);
xor U3055 (N_3055,N_2668,N_1771);
and U3056 (N_3056,N_1582,N_1717);
or U3057 (N_3057,N_2938,N_2688);
xor U3058 (N_3058,N_2192,N_1962);
and U3059 (N_3059,N_2372,N_1738);
xnor U3060 (N_3060,N_1952,N_1535);
nor U3061 (N_3061,N_2741,N_2023);
or U3062 (N_3062,N_1689,N_2298);
or U3063 (N_3063,N_2245,N_2009);
and U3064 (N_3064,N_2832,N_1718);
xnor U3065 (N_3065,N_2531,N_2133);
or U3066 (N_3066,N_2998,N_2269);
nand U3067 (N_3067,N_1736,N_2540);
nand U3068 (N_3068,N_1618,N_1720);
nand U3069 (N_3069,N_2823,N_2434);
xor U3070 (N_3070,N_2852,N_1979);
and U3071 (N_3071,N_2125,N_1860);
or U3072 (N_3072,N_2474,N_2631);
or U3073 (N_3073,N_2072,N_2216);
xor U3074 (N_3074,N_2930,N_1638);
xor U3075 (N_3075,N_2991,N_1804);
nor U3076 (N_3076,N_1940,N_2803);
xnor U3077 (N_3077,N_2203,N_1814);
or U3078 (N_3078,N_2257,N_2493);
or U3079 (N_3079,N_2770,N_2929);
xnor U3080 (N_3080,N_2275,N_1628);
or U3081 (N_3081,N_1819,N_1778);
or U3082 (N_3082,N_2855,N_2986);
xnor U3083 (N_3083,N_2538,N_2969);
and U3084 (N_3084,N_2184,N_2113);
and U3085 (N_3085,N_1621,N_2270);
or U3086 (N_3086,N_1602,N_1823);
or U3087 (N_3087,N_2158,N_1868);
or U3088 (N_3088,N_1549,N_2123);
nand U3089 (N_3089,N_2900,N_1957);
xor U3090 (N_3090,N_1891,N_2757);
nor U3091 (N_3091,N_2397,N_2352);
nand U3092 (N_3092,N_2624,N_1878);
nor U3093 (N_3093,N_1672,N_2116);
or U3094 (N_3094,N_2338,N_2340);
or U3095 (N_3095,N_2339,N_1655);
nor U3096 (N_3096,N_2402,N_1629);
and U3097 (N_3097,N_2436,N_2324);
nor U3098 (N_3098,N_2144,N_2309);
or U3099 (N_3099,N_1731,N_1630);
xor U3100 (N_3100,N_2819,N_1813);
nor U3101 (N_3101,N_2268,N_2676);
and U3102 (N_3102,N_1707,N_2953);
and U3103 (N_3103,N_1608,N_2409);
and U3104 (N_3104,N_1844,N_2640);
or U3105 (N_3105,N_2626,N_2326);
nand U3106 (N_3106,N_2563,N_2066);
nand U3107 (N_3107,N_1532,N_2202);
or U3108 (N_3108,N_2579,N_2512);
nand U3109 (N_3109,N_2126,N_2271);
or U3110 (N_3110,N_1960,N_1546);
nand U3111 (N_3111,N_2957,N_2955);
or U3112 (N_3112,N_1935,N_2199);
or U3113 (N_3113,N_2127,N_2977);
xnor U3114 (N_3114,N_2618,N_2858);
nor U3115 (N_3115,N_2565,N_1675);
or U3116 (N_3116,N_1827,N_2322);
and U3117 (N_3117,N_2951,N_2342);
or U3118 (N_3118,N_2080,N_1744);
xnor U3119 (N_3119,N_1742,N_1528);
nand U3120 (N_3120,N_1695,N_1551);
and U3121 (N_3121,N_1679,N_2699);
and U3122 (N_3122,N_1853,N_1651);
or U3123 (N_3123,N_2863,N_1972);
or U3124 (N_3124,N_1956,N_2607);
and U3125 (N_3125,N_1547,N_2049);
or U3126 (N_3126,N_1613,N_1553);
or U3127 (N_3127,N_1998,N_2593);
nor U3128 (N_3128,N_2703,N_1843);
nand U3129 (N_3129,N_1712,N_2086);
xor U3130 (N_3130,N_1848,N_1936);
nand U3131 (N_3131,N_2101,N_2600);
nor U3132 (N_3132,N_2537,N_1864);
or U3133 (N_3133,N_1527,N_1888);
xnor U3134 (N_3134,N_2636,N_2454);
nor U3135 (N_3135,N_2059,N_2451);
or U3136 (N_3136,N_1680,N_2604);
and U3137 (N_3137,N_2445,N_2170);
nor U3138 (N_3138,N_2044,N_2177);
and U3139 (N_3139,N_2910,N_2888);
xnor U3140 (N_3140,N_1627,N_2093);
and U3141 (N_3141,N_1586,N_2693);
nand U3142 (N_3142,N_2061,N_2151);
or U3143 (N_3143,N_2628,N_1561);
or U3144 (N_3144,N_2571,N_2258);
nor U3145 (N_3145,N_2767,N_2207);
and U3146 (N_3146,N_2155,N_1656);
nand U3147 (N_3147,N_2896,N_2868);
and U3148 (N_3148,N_2014,N_1834);
nor U3149 (N_3149,N_2873,N_2104);
or U3150 (N_3150,N_2567,N_2385);
nor U3151 (N_3151,N_2572,N_2260);
nand U3152 (N_3152,N_2905,N_1846);
nor U3153 (N_3153,N_2950,N_2547);
nand U3154 (N_3154,N_2619,N_2750);
or U3155 (N_3155,N_1711,N_2610);
nand U3156 (N_3156,N_1808,N_1737);
or U3157 (N_3157,N_2759,N_2821);
nor U3158 (N_3158,N_2833,N_2252);
nor U3159 (N_3159,N_1845,N_2129);
xnor U3160 (N_3160,N_2272,N_1636);
and U3161 (N_3161,N_1650,N_1906);
or U3162 (N_3162,N_2096,N_1784);
and U3163 (N_3163,N_2892,N_1698);
xnor U3164 (N_3164,N_2037,N_2801);
and U3165 (N_3165,N_1874,N_2671);
or U3166 (N_3166,N_2812,N_2313);
or U3167 (N_3167,N_1794,N_2303);
nor U3168 (N_3168,N_2779,N_2483);
nor U3169 (N_3169,N_1964,N_2961);
xor U3170 (N_3170,N_1926,N_2107);
nand U3171 (N_3171,N_2394,N_1539);
and U3172 (N_3172,N_2358,N_1918);
nand U3173 (N_3173,N_2375,N_1982);
and U3174 (N_3174,N_2570,N_1785);
and U3175 (N_3175,N_2878,N_2359);
nor U3176 (N_3176,N_1709,N_2842);
nand U3177 (N_3177,N_2638,N_1978);
or U3178 (N_3178,N_1531,N_2904);
xor U3179 (N_3179,N_2012,N_1748);
nand U3180 (N_3180,N_2089,N_1601);
nor U3181 (N_3181,N_2283,N_2669);
and U3182 (N_3182,N_2415,N_1706);
and U3183 (N_3183,N_2193,N_2327);
nor U3184 (N_3184,N_2188,N_2046);
or U3185 (N_3185,N_1668,N_1665);
nand U3186 (N_3186,N_2112,N_2948);
and U3187 (N_3187,N_1734,N_2914);
xnor U3188 (N_3188,N_1912,N_1839);
nand U3189 (N_3189,N_1842,N_1802);
xor U3190 (N_3190,N_1991,N_2943);
nand U3191 (N_3191,N_2404,N_2613);
nand U3192 (N_3192,N_2911,N_1757);
xnor U3193 (N_3193,N_2054,N_2690);
nand U3194 (N_3194,N_2460,N_2648);
and U3195 (N_3195,N_1591,N_2353);
or U3196 (N_3196,N_1806,N_2698);
or U3197 (N_3197,N_1902,N_2952);
or U3198 (N_3198,N_2576,N_2036);
and U3199 (N_3199,N_1920,N_2016);
xnor U3200 (N_3200,N_2795,N_2514);
nand U3201 (N_3201,N_1544,N_2239);
and U3202 (N_3202,N_1740,N_1677);
nand U3203 (N_3203,N_2095,N_2939);
or U3204 (N_3204,N_1781,N_1773);
or U3205 (N_3205,N_2027,N_2602);
xor U3206 (N_3206,N_2185,N_1803);
and U3207 (N_3207,N_1764,N_2186);
or U3208 (N_3208,N_1767,N_1540);
or U3209 (N_3209,N_1662,N_2763);
nand U3210 (N_3210,N_2449,N_1519);
nor U3211 (N_3211,N_2528,N_1908);
nor U3212 (N_3212,N_1597,N_2208);
xor U3213 (N_3213,N_2854,N_1741);
nor U3214 (N_3214,N_2032,N_2656);
nor U3215 (N_3215,N_2287,N_2886);
nand U3216 (N_3216,N_2561,N_2836);
or U3217 (N_3217,N_2777,N_1639);
or U3218 (N_3218,N_1829,N_1728);
nor U3219 (N_3219,N_2442,N_2612);
and U3220 (N_3220,N_2752,N_2783);
and U3221 (N_3221,N_2337,N_2805);
or U3222 (N_3222,N_2555,N_2764);
nor U3223 (N_3223,N_2091,N_1580);
xnor U3224 (N_3224,N_1726,N_2181);
nor U3225 (N_3225,N_2924,N_1904);
or U3226 (N_3226,N_2219,N_2840);
xnor U3227 (N_3227,N_2078,N_2400);
xnor U3228 (N_3228,N_2154,N_1754);
nor U3229 (N_3229,N_1716,N_2535);
xnor U3230 (N_3230,N_2716,N_2918);
or U3231 (N_3231,N_1710,N_2794);
and U3232 (N_3232,N_2508,N_2074);
or U3233 (N_3233,N_2261,N_2062);
nand U3234 (N_3234,N_2799,N_1526);
and U3235 (N_3235,N_2574,N_2749);
nand U3236 (N_3236,N_2282,N_1900);
nand U3237 (N_3237,N_2335,N_2330);
nand U3238 (N_3238,N_2040,N_1749);
nand U3239 (N_3239,N_2647,N_2020);
xnor U3240 (N_3240,N_2546,N_2554);
nand U3241 (N_3241,N_1985,N_1974);
xnor U3242 (N_3242,N_2465,N_2968);
nand U3243 (N_3243,N_2711,N_2517);
nand U3244 (N_3244,N_1805,N_1893);
nand U3245 (N_3245,N_2681,N_2484);
or U3246 (N_3246,N_2236,N_2877);
nand U3247 (N_3247,N_2190,N_2573);
xnor U3248 (N_3248,N_1861,N_1568);
or U3249 (N_3249,N_1899,N_1669);
xor U3250 (N_3250,N_1898,N_2468);
or U3251 (N_3251,N_1822,N_2256);
nor U3252 (N_3252,N_2458,N_1593);
nor U3253 (N_3253,N_1815,N_2639);
or U3254 (N_3254,N_2609,N_1626);
xnor U3255 (N_3255,N_1612,N_2603);
nand U3256 (N_3256,N_2425,N_2028);
xnor U3257 (N_3257,N_1782,N_1963);
nand U3258 (N_3258,N_1801,N_2599);
nor U3259 (N_3259,N_2704,N_1607);
nor U3260 (N_3260,N_2527,N_1934);
and U3261 (N_3261,N_1879,N_2228);
nor U3262 (N_3262,N_2601,N_1915);
xnor U3263 (N_3263,N_2143,N_2029);
and U3264 (N_3264,N_1947,N_2247);
xnor U3265 (N_3265,N_2179,N_2897);
nand U3266 (N_3266,N_2921,N_1615);
nor U3267 (N_3267,N_2872,N_2963);
or U3268 (N_3268,N_2707,N_2743);
or U3269 (N_3269,N_1774,N_1816);
nand U3270 (N_3270,N_1896,N_2592);
and U3271 (N_3271,N_2685,N_2959);
xor U3272 (N_3272,N_2097,N_2168);
nor U3273 (N_3273,N_2350,N_2153);
nand U3274 (N_3274,N_2075,N_2211);
xnor U3275 (N_3275,N_1755,N_2804);
nand U3276 (N_3276,N_2008,N_2867);
nand U3277 (N_3277,N_2428,N_2616);
nand U3278 (N_3278,N_2115,N_1913);
nor U3279 (N_3279,N_2694,N_2865);
nor U3280 (N_3280,N_1520,N_2343);
or U3281 (N_3281,N_2387,N_1570);
and U3282 (N_3282,N_2146,N_2377);
nand U3283 (N_3283,N_1595,N_2388);
or U3284 (N_3284,N_2427,N_2280);
and U3285 (N_3285,N_2680,N_1666);
nand U3286 (N_3286,N_2504,N_1820);
and U3287 (N_3287,N_2182,N_1566);
nand U3288 (N_3288,N_2695,N_2407);
nand U3289 (N_3289,N_2135,N_1876);
nor U3290 (N_3290,N_2513,N_2305);
and U3291 (N_3291,N_2866,N_2662);
nand U3292 (N_3292,N_2543,N_2167);
and U3293 (N_3293,N_1633,N_2846);
xor U3294 (N_3294,N_2487,N_2784);
xnor U3295 (N_3295,N_2725,N_1708);
nor U3296 (N_3296,N_2818,N_2336);
nand U3297 (N_3297,N_1558,N_2022);
nor U3298 (N_3298,N_1701,N_2507);
nand U3299 (N_3299,N_1975,N_1990);
or U3300 (N_3300,N_1505,N_2548);
nor U3301 (N_3301,N_2917,N_1786);
nand U3302 (N_3302,N_2849,N_2156);
and U3303 (N_3303,N_2768,N_2802);
nand U3304 (N_3304,N_1976,N_1907);
nor U3305 (N_3305,N_2591,N_1942);
xnor U3306 (N_3306,N_2843,N_1694);
nand U3307 (N_3307,N_1944,N_2002);
xnor U3308 (N_3308,N_2841,N_2940);
and U3309 (N_3309,N_2765,N_1730);
xor U3310 (N_3310,N_2810,N_2820);
xor U3311 (N_3311,N_2979,N_2720);
nand U3312 (N_3312,N_1759,N_2837);
nand U3313 (N_3313,N_1838,N_2525);
xor U3314 (N_3314,N_2455,N_2826);
and U3315 (N_3315,N_2899,N_1758);
or U3316 (N_3316,N_1654,N_1598);
nand U3317 (N_3317,N_1811,N_1939);
xor U3318 (N_3318,N_2294,N_1821);
xor U3319 (N_3319,N_2238,N_1895);
nor U3320 (N_3320,N_2912,N_1577);
nand U3321 (N_3321,N_2092,N_1931);
xnor U3322 (N_3322,N_1746,N_2401);
nand U3323 (N_3323,N_2992,N_2018);
and U3324 (N_3324,N_2210,N_2675);
and U3325 (N_3325,N_2346,N_2325);
nor U3326 (N_3326,N_2557,N_2470);
or U3327 (N_3327,N_1620,N_2937);
and U3328 (N_3328,N_2495,N_2630);
or U3329 (N_3329,N_2614,N_2296);
or U3330 (N_3330,N_2164,N_1733);
xor U3331 (N_3331,N_1930,N_2111);
nand U3332 (N_3332,N_2226,N_1583);
and U3333 (N_3333,N_2300,N_2551);
nand U3334 (N_3334,N_1852,N_2444);
nor U3335 (N_3335,N_2085,N_2486);
xor U3336 (N_3336,N_2850,N_1872);
xor U3337 (N_3337,N_2882,N_2003);
xnor U3338 (N_3338,N_2480,N_2769);
nand U3339 (N_3339,N_2978,N_1969);
nand U3340 (N_3340,N_1576,N_1807);
or U3341 (N_3341,N_1954,N_1966);
xor U3342 (N_3342,N_2319,N_1652);
or U3343 (N_3343,N_2898,N_2633);
and U3344 (N_3344,N_2994,N_2230);
or U3345 (N_3345,N_2931,N_1850);
nor U3346 (N_3346,N_2597,N_2138);
and U3347 (N_3347,N_1903,N_1983);
nand U3348 (N_3348,N_1909,N_2047);
nand U3349 (N_3349,N_2919,N_2787);
and U3350 (N_3350,N_2440,N_2437);
nor U3351 (N_3351,N_2289,N_1923);
nand U3352 (N_3352,N_2021,N_1658);
xnor U3353 (N_3353,N_1530,N_2422);
nand U3354 (N_3354,N_2152,N_2646);
and U3355 (N_3355,N_2290,N_2566);
nand U3356 (N_3356,N_1713,N_1953);
or U3357 (N_3357,N_2890,N_1703);
and U3358 (N_3358,N_2430,N_2995);
and U3359 (N_3359,N_1763,N_2972);
or U3360 (N_3360,N_2539,N_2932);
xnor U3361 (N_3361,N_2162,N_2736);
or U3362 (N_3362,N_2973,N_1682);
or U3363 (N_3363,N_2310,N_1606);
nand U3364 (N_3364,N_2887,N_2773);
nor U3365 (N_3365,N_1600,N_2011);
and U3366 (N_3366,N_1769,N_2587);
and U3367 (N_3367,N_1578,N_2317);
nand U3368 (N_3368,N_1830,N_1854);
nor U3369 (N_3369,N_1515,N_2291);
nand U3370 (N_3370,N_2222,N_2263);
nand U3371 (N_3371,N_2622,N_2893);
xor U3372 (N_3372,N_1660,N_1715);
nand U3373 (N_3373,N_2778,N_2700);
xnor U3374 (N_3374,N_2119,N_2560);
nand U3375 (N_3375,N_2448,N_1614);
xnor U3376 (N_3376,N_1649,N_2344);
or U3377 (N_3377,N_2605,N_1828);
nand U3378 (N_3378,N_2578,N_2715);
nand U3379 (N_3379,N_2443,N_1699);
and U3380 (N_3380,N_1922,N_2881);
nor U3381 (N_3381,N_1722,N_2169);
or U3382 (N_3382,N_2412,N_2039);
xnor U3383 (N_3383,N_1508,N_1880);
xor U3384 (N_3384,N_2580,N_2860);
nor U3385 (N_3385,N_1890,N_1750);
nor U3386 (N_3386,N_1504,N_1529);
nand U3387 (N_3387,N_2569,N_1797);
or U3388 (N_3388,N_2248,N_2391);
or U3389 (N_3389,N_2063,N_2051);
nor U3390 (N_3390,N_1955,N_2235);
nand U3391 (N_3391,N_2731,N_1721);
nor U3392 (N_3392,N_1604,N_2383);
nor U3393 (N_3393,N_1563,N_2374);
or U3394 (N_3394,N_2246,N_1684);
and U3395 (N_3395,N_1700,N_2632);
and U3396 (N_3396,N_1637,N_2447);
nand U3397 (N_3397,N_1768,N_2723);
or U3398 (N_3398,N_1683,N_1533);
and U3399 (N_3399,N_2477,N_2780);
nand U3400 (N_3400,N_1747,N_2729);
or U3401 (N_3401,N_2357,N_2217);
nand U3402 (N_3402,N_2532,N_2982);
nor U3403 (N_3403,N_1800,N_2173);
nand U3404 (N_3404,N_2935,N_1503);
or U3405 (N_3405,N_2673,N_2666);
and U3406 (N_3406,N_1910,N_2734);
and U3407 (N_3407,N_1847,N_2903);
nand U3408 (N_3408,N_1511,N_2934);
and U3409 (N_3409,N_2481,N_2347);
or U3410 (N_3410,N_1671,N_1832);
xnor U3411 (N_3411,N_1631,N_2923);
xnor U3412 (N_3412,N_2315,N_2534);
and U3413 (N_3413,N_1836,N_2265);
nand U3414 (N_3414,N_2751,N_2033);
and U3415 (N_3415,N_1863,N_1705);
nand U3416 (N_3416,N_1688,N_2253);
xor U3417 (N_3417,N_1663,N_2758);
nor U3418 (N_3418,N_1623,N_2035);
or U3419 (N_3419,N_2368,N_2687);
xnor U3420 (N_3420,N_1697,N_2273);
nor U3421 (N_3421,N_2332,N_1881);
or U3422 (N_3422,N_2114,N_2891);
nor U3423 (N_3423,N_2811,N_1866);
or U3424 (N_3424,N_1512,N_2172);
or U3425 (N_3425,N_2740,N_2302);
nor U3426 (N_3426,N_2090,N_1523);
xnor U3427 (N_3427,N_1916,N_2431);
xor U3428 (N_3428,N_1594,N_1640);
nor U3429 (N_3429,N_1970,N_2042);
or U3430 (N_3430,N_2013,N_2249);
or U3431 (N_3431,N_2233,N_2753);
xnor U3432 (N_3432,N_2259,N_1727);
xnor U3433 (N_3433,N_1534,N_2989);
nand U3434 (N_3434,N_2464,N_2195);
or U3435 (N_3435,N_1812,N_2478);
or U3436 (N_3436,N_2364,N_2869);
nor U3437 (N_3437,N_1980,N_1933);
nor U3438 (N_3438,N_1790,N_1973);
xor U3439 (N_3439,N_2057,N_2034);
or U3440 (N_3440,N_2435,N_2070);
or U3441 (N_3441,N_1653,N_1921);
nand U3442 (N_3442,N_2718,N_2506);
nand U3443 (N_3443,N_1552,N_2761);
nand U3444 (N_3444,N_2476,N_1555);
nand U3445 (N_3445,N_2424,N_2708);
nand U3446 (N_3446,N_2775,N_1772);
and U3447 (N_3447,N_1635,N_1524);
and U3448 (N_3448,N_2889,N_2363);
and U3449 (N_3449,N_2874,N_2822);
and U3450 (N_3450,N_2079,N_1877);
nor U3451 (N_3451,N_2664,N_1766);
or U3452 (N_3452,N_2542,N_2240);
or U3453 (N_3453,N_2590,N_2582);
or U3454 (N_3454,N_2641,N_1948);
and U3455 (N_3455,N_1798,N_2595);
and U3456 (N_3456,N_2220,N_2026);
nor U3457 (N_3457,N_1770,N_2365);
xor U3458 (N_3458,N_2212,N_2562);
or U3459 (N_3459,N_2088,N_2159);
nand U3460 (N_3460,N_1927,N_2583);
nor U3461 (N_3461,N_2150,N_1732);
nand U3462 (N_3462,N_1984,N_2254);
nor U3463 (N_3463,N_1791,N_2348);
xnor U3464 (N_3464,N_2677,N_2575);
or U3465 (N_3465,N_2654,N_1571);
nor U3466 (N_3466,N_2984,N_2069);
and U3467 (N_3467,N_1690,N_2065);
nand U3468 (N_3468,N_2625,N_2321);
xnor U3469 (N_3469,N_2629,N_2617);
and U3470 (N_3470,N_2297,N_1858);
nor U3471 (N_3471,N_1729,N_2974);
nand U3472 (N_3472,N_1617,N_2134);
or U3473 (N_3473,N_2774,N_2081);
or U3474 (N_3474,N_2936,N_2649);
and U3475 (N_3475,N_2145,N_2985);
and U3476 (N_3476,N_2526,N_2853);
nor U3477 (N_3477,N_1691,N_1554);
and U3478 (N_3478,N_2083,N_1901);
and U3479 (N_3479,N_2314,N_1575);
and U3480 (N_3480,N_2672,N_2857);
nor U3481 (N_3481,N_2067,N_2847);
nand U3482 (N_3482,N_2277,N_1719);
xnor U3483 (N_3483,N_2824,N_2206);
nor U3484 (N_3484,N_2349,N_2674);
nor U3485 (N_3485,N_2993,N_1999);
nand U3486 (N_3486,N_1596,N_2608);
and U3487 (N_3487,N_2052,N_2499);
nand U3488 (N_3488,N_2721,N_2413);
xnor U3489 (N_3489,N_2864,N_2568);
and U3490 (N_3490,N_1776,N_1857);
and U3491 (N_3491,N_1525,N_2299);
nand U3492 (N_3492,N_1743,N_2304);
or U3493 (N_3493,N_2663,N_1502);
or U3494 (N_3494,N_2370,N_2643);
nor U3495 (N_3495,N_2509,N_2323);
xnor U3496 (N_3496,N_2652,N_2713);
and U3497 (N_3497,N_2956,N_1609);
and U3498 (N_3498,N_2724,N_2108);
xnor U3499 (N_3499,N_2077,N_1579);
and U3500 (N_3500,N_1951,N_2420);
xor U3501 (N_3501,N_1646,N_2657);
nand U3502 (N_3502,N_1959,N_1795);
or U3503 (N_3503,N_1564,N_2379);
nand U3504 (N_3504,N_1992,N_2738);
or U3505 (N_3505,N_2043,N_1541);
or U3506 (N_3506,N_1756,N_2594);
and U3507 (N_3507,N_2267,N_1509);
nor U3508 (N_3508,N_1961,N_2122);
xnor U3509 (N_3509,N_2800,N_1870);
xnor U3510 (N_3510,N_2378,N_1685);
or U3511 (N_3511,N_2665,N_2227);
and U3512 (N_3512,N_2502,N_2831);
and U3513 (N_3513,N_2292,N_2243);
and U3514 (N_3514,N_2328,N_2362);
and U3515 (N_3515,N_2981,N_1687);
and U3516 (N_3516,N_1817,N_2845);
nor U3517 (N_3517,N_2885,N_1536);
or U3518 (N_3518,N_2471,N_2732);
or U3519 (N_3519,N_2019,N_2644);
and U3520 (N_3520,N_2453,N_1567);
xor U3521 (N_3521,N_2789,N_2174);
or U3522 (N_3522,N_1994,N_2200);
nor U3523 (N_3523,N_2264,N_1929);
nor U3524 (N_3524,N_2667,N_2856);
xnor U3525 (N_3525,N_2744,N_2909);
xnor U3526 (N_3526,N_2825,N_1647);
nand U3527 (N_3527,N_1585,N_1905);
nand U3528 (N_3528,N_2187,N_1605);
nand U3529 (N_3529,N_1581,N_1765);
nand U3530 (N_3530,N_2660,N_1835);
and U3531 (N_3531,N_2176,N_2611);
or U3532 (N_3532,N_2004,N_2682);
and U3533 (N_3533,N_1859,N_2398);
nand U3534 (N_3534,N_1661,N_1818);
nand U3535 (N_3535,N_2717,N_1634);
and U3536 (N_3536,N_2137,N_2679);
and U3537 (N_3537,N_2788,N_1603);
and U3538 (N_3538,N_2772,N_1696);
or U3539 (N_3539,N_2623,N_2645);
nor U3540 (N_3540,N_2908,N_1833);
or U3541 (N_3541,N_2606,N_2163);
or U3542 (N_3542,N_2405,N_2658);
nor U3543 (N_3543,N_2421,N_2945);
and U3544 (N_3544,N_1589,N_2691);
nand U3545 (N_3545,N_1981,N_2511);
and U3546 (N_3546,N_1989,N_1599);
nand U3547 (N_3547,N_1510,N_2136);
and U3548 (N_3548,N_2189,N_2970);
xor U3549 (N_3549,N_2790,N_2279);
nor U3550 (N_3550,N_2118,N_2722);
or U3551 (N_3551,N_1673,N_2786);
nor U3552 (N_3552,N_2519,N_2637);
and U3553 (N_3553,N_1648,N_2650);
xor U3554 (N_3554,N_2102,N_1670);
and U3555 (N_3555,N_2432,N_2295);
or U3556 (N_3556,N_2714,N_2414);
or U3557 (N_3557,N_2586,N_2906);
and U3558 (N_3558,N_2653,N_1796);
and U3559 (N_3559,N_2692,N_2354);
or U3560 (N_3560,N_2380,N_2902);
nor U3561 (N_3561,N_2369,N_2971);
nor U3562 (N_3562,N_2416,N_1592);
xnor U3563 (N_3563,N_2500,N_1678);
and U3564 (N_3564,N_1968,N_2234);
nand U3565 (N_3565,N_1775,N_2705);
and U3566 (N_3566,N_1501,N_2395);
and U3567 (N_3567,N_1522,N_2386);
nand U3568 (N_3568,N_2130,N_2988);
or U3569 (N_3569,N_2678,N_1751);
and U3570 (N_3570,N_2926,N_1745);
nand U3571 (N_3571,N_2661,N_2696);
nor U3572 (N_3572,N_1894,N_1941);
xor U3573 (N_3573,N_1762,N_2110);
xor U3574 (N_3574,N_2382,N_2438);
nand U3575 (N_3575,N_2423,N_1521);
or U3576 (N_3576,N_2148,N_2830);
or U3577 (N_3577,N_2947,N_1882);
nand U3578 (N_3578,N_1987,N_2894);
nand U3579 (N_3579,N_2048,N_2284);
or U3580 (N_3580,N_2949,N_2895);
xor U3581 (N_3581,N_1841,N_2927);
and U3582 (N_3582,N_1557,N_2007);
and U3583 (N_3583,N_2417,N_1793);
nand U3584 (N_3584,N_2754,N_2316);
xnor U3585 (N_3585,N_1686,N_2197);
or U3586 (N_3586,N_2082,N_2225);
or U3587 (N_3587,N_2798,N_2178);
nor U3588 (N_3588,N_1641,N_2384);
nor U3589 (N_3589,N_2360,N_1938);
and U3590 (N_3590,N_2366,N_1883);
nand U3591 (N_3591,N_1681,N_2333);
or U3592 (N_3592,N_2503,N_2518);
nand U3593 (N_3593,N_1516,N_2466);
nor U3594 (N_3594,N_1840,N_2120);
or U3595 (N_3595,N_2139,N_2479);
nand U3596 (N_3596,N_2615,N_2859);
xor U3597 (N_3597,N_2419,N_1507);
xor U3598 (N_3598,N_1914,N_2975);
or U3599 (N_3599,N_2806,N_1513);
nand U3600 (N_3600,N_1588,N_2492);
or U3601 (N_3601,N_2544,N_2683);
nand U3602 (N_3602,N_2516,N_2791);
nand U3603 (N_3603,N_2329,N_1865);
or U3604 (N_3604,N_2807,N_2276);
nand U3605 (N_3605,N_1610,N_2376);
and U3606 (N_3606,N_1949,N_2814);
or U3607 (N_3607,N_2880,N_2879);
xnor U3608 (N_3608,N_1548,N_2838);
or U3609 (N_3609,N_1997,N_2496);
nor U3610 (N_3610,N_1704,N_2907);
nor U3611 (N_3611,N_1869,N_2489);
or U3612 (N_3612,N_2055,N_1825);
and U3613 (N_3613,N_1810,N_1937);
and U3614 (N_3614,N_2301,N_2550);
or U3615 (N_3615,N_1945,N_1885);
nand U3616 (N_3616,N_2796,N_2739);
or U3617 (N_3617,N_2161,N_2726);
and U3618 (N_3618,N_2635,N_2175);
and U3619 (N_3619,N_1739,N_2121);
and U3620 (N_3620,N_2073,N_2771);
nand U3621 (N_3621,N_1537,N_2515);
nor U3622 (N_3622,N_2746,N_1624);
and U3623 (N_3623,N_2727,N_2642);
nor U3624 (N_3624,N_2627,N_2915);
and U3625 (N_3625,N_2106,N_2488);
nor U3626 (N_3626,N_2371,N_2141);
or U3627 (N_3627,N_1977,N_2475);
and U3628 (N_3628,N_2244,N_2373);
xor U3629 (N_3629,N_2140,N_2456);
and U3630 (N_3630,N_1967,N_1659);
nor U3631 (N_3631,N_2214,N_1657);
nor U3632 (N_3632,N_2965,N_2285);
or U3633 (N_3633,N_2094,N_2737);
and U3634 (N_3634,N_2274,N_2862);
nand U3635 (N_3635,N_2748,N_2797);
xor U3636 (N_3636,N_1676,N_2293);
or U3637 (N_3637,N_2839,N_2201);
xor U3638 (N_3638,N_2038,N_1760);
nor U3639 (N_3639,N_2967,N_2209);
and U3640 (N_3640,N_2813,N_2549);
or U3641 (N_3641,N_2933,N_2620);
xnor U3642 (N_3642,N_1789,N_2452);
and U3643 (N_3643,N_2581,N_2015);
and U3644 (N_3644,N_1565,N_1892);
nor U3645 (N_3645,N_2223,N_1643);
xnor U3646 (N_3646,N_2745,N_1645);
nor U3647 (N_3647,N_2999,N_2165);
and U3648 (N_3648,N_2521,N_2762);
nor U3649 (N_3649,N_2966,N_2808);
nor U3650 (N_3650,N_2491,N_2462);
and U3651 (N_3651,N_2541,N_2980);
xnor U3652 (N_3652,N_2533,N_2320);
xnor U3653 (N_3653,N_1986,N_2334);
or U3654 (N_3654,N_2925,N_2996);
nor U3655 (N_3655,N_1971,N_1569);
xnor U3656 (N_3656,N_2393,N_2976);
and U3657 (N_3657,N_2031,N_1988);
xor U3658 (N_3658,N_2817,N_2875);
nand U3659 (N_3659,N_1995,N_2060);
or U3660 (N_3660,N_2997,N_2262);
nor U3661 (N_3661,N_1611,N_2250);
nand U3662 (N_3662,N_2983,N_2071);
and U3663 (N_3663,N_2529,N_2396);
nor U3664 (N_3664,N_1556,N_2710);
nor U3665 (N_3665,N_2510,N_2530);
nor U3666 (N_3666,N_2204,N_2087);
and U3667 (N_3667,N_2954,N_2221);
xor U3668 (N_3668,N_2446,N_2884);
xor U3669 (N_3669,N_1542,N_2160);
xnor U3670 (N_3670,N_2418,N_2962);
xnor U3671 (N_3671,N_2058,N_2883);
or U3672 (N_3672,N_2689,N_2827);
xnor U3673 (N_3673,N_2191,N_2861);
or U3674 (N_3674,N_1849,N_1562);
xnor U3675 (N_3675,N_2441,N_2010);
nor U3676 (N_3676,N_2922,N_2312);
nand U3677 (N_3677,N_2848,N_2697);
nand U3678 (N_3678,N_2194,N_2171);
nor U3679 (N_3679,N_2659,N_2621);
or U3680 (N_3680,N_1924,N_2901);
and U3681 (N_3681,N_2068,N_1826);
or U3682 (N_3682,N_2520,N_2920);
and U3683 (N_3683,N_2109,N_2461);
and U3684 (N_3684,N_2670,N_1724);
or U3685 (N_3685,N_2041,N_1862);
xor U3686 (N_3686,N_2105,N_1545);
xor U3687 (N_3687,N_2367,N_1735);
or U3688 (N_3688,N_2467,N_1809);
xnor U3689 (N_3689,N_2498,N_2166);
and U3690 (N_3690,N_2776,N_2490);
and U3691 (N_3691,N_2719,N_1787);
or U3692 (N_3692,N_2815,N_2781);
nor U3693 (N_3693,N_2651,N_1837);
and U3694 (N_3694,N_1664,N_2100);
and U3695 (N_3695,N_1723,N_1799);
nor U3696 (N_3696,N_2942,N_2536);
and U3697 (N_3697,N_2589,N_2381);
nor U3698 (N_3698,N_1560,N_1946);
nor U3699 (N_3699,N_2870,N_2389);
and U3700 (N_3700,N_2341,N_1584);
nor U3701 (N_3701,N_1867,N_2084);
nand U3702 (N_3702,N_1950,N_2351);
nor U3703 (N_3703,N_2960,N_2990);
or U3704 (N_3704,N_1889,N_2755);
nor U3705 (N_3705,N_2835,N_2505);
and U3706 (N_3706,N_1779,N_2045);
and U3707 (N_3707,N_2132,N_2793);
and U3708 (N_3708,N_2596,N_1725);
and U3709 (N_3709,N_2142,N_2117);
nor U3710 (N_3710,N_2000,N_2785);
and U3711 (N_3711,N_2733,N_2318);
xor U3712 (N_3712,N_2406,N_1506);
xnor U3713 (N_3713,N_1932,N_2553);
nand U3714 (N_3714,N_1928,N_1897);
xor U3715 (N_3715,N_2756,N_1702);
and U3716 (N_3716,N_2760,N_1943);
or U3717 (N_3717,N_2128,N_1517);
or U3718 (N_3718,N_2099,N_2876);
and U3719 (N_3719,N_2473,N_2306);
or U3720 (N_3720,N_2308,N_1753);
nand U3721 (N_3721,N_1856,N_2286);
nand U3722 (N_3722,N_2730,N_2147);
xnor U3723 (N_3723,N_2399,N_1965);
and U3724 (N_3724,N_1538,N_2482);
xor U3725 (N_3725,N_2361,N_1514);
nand U3726 (N_3726,N_2251,N_2871);
nand U3727 (N_3727,N_2829,N_2241);
nand U3728 (N_3728,N_2834,N_2215);
nor U3729 (N_3729,N_2218,N_2523);
nor U3730 (N_3730,N_2356,N_1587);
and U3731 (N_3731,N_2131,N_2278);
and U3732 (N_3732,N_2076,N_2494);
or U3733 (N_3733,N_2098,N_1780);
nor U3734 (N_3734,N_1573,N_1831);
or U3735 (N_3735,N_1958,N_2501);
or U3736 (N_3736,N_2410,N_2433);
xnor U3737 (N_3737,N_2198,N_2701);
xor U3738 (N_3738,N_1543,N_2196);
or U3739 (N_3739,N_2816,N_1993);
xnor U3740 (N_3740,N_2469,N_2403);
nor U3741 (N_3741,N_2792,N_2964);
and U3742 (N_3742,N_2766,N_2851);
nand U3743 (N_3743,N_2411,N_1788);
nand U3744 (N_3744,N_2742,N_2024);
and U3745 (N_3745,N_1622,N_1887);
and U3746 (N_3746,N_2426,N_2213);
xor U3747 (N_3747,N_2987,N_2522);
nand U3748 (N_3748,N_2916,N_1783);
nand U3749 (N_3749,N_2345,N_1824);
nand U3750 (N_3750,N_1575,N_2567);
nand U3751 (N_3751,N_2209,N_2317);
or U3752 (N_3752,N_2213,N_1725);
or U3753 (N_3753,N_2353,N_1821);
xnor U3754 (N_3754,N_1846,N_2950);
or U3755 (N_3755,N_2705,N_1960);
and U3756 (N_3756,N_2142,N_2534);
nand U3757 (N_3757,N_2423,N_2731);
xnor U3758 (N_3758,N_1573,N_2325);
nand U3759 (N_3759,N_2195,N_2797);
nor U3760 (N_3760,N_2855,N_2683);
nand U3761 (N_3761,N_2768,N_2652);
and U3762 (N_3762,N_1503,N_2791);
or U3763 (N_3763,N_2918,N_1758);
or U3764 (N_3764,N_1514,N_2659);
xor U3765 (N_3765,N_2681,N_1846);
or U3766 (N_3766,N_2702,N_2802);
nand U3767 (N_3767,N_2515,N_1670);
nor U3768 (N_3768,N_1609,N_2096);
nor U3769 (N_3769,N_1584,N_2003);
and U3770 (N_3770,N_2846,N_1931);
xor U3771 (N_3771,N_2379,N_2770);
and U3772 (N_3772,N_2809,N_2813);
xor U3773 (N_3773,N_2599,N_2821);
xnor U3774 (N_3774,N_2372,N_2968);
nor U3775 (N_3775,N_2770,N_1718);
nand U3776 (N_3776,N_2322,N_2013);
or U3777 (N_3777,N_2093,N_1527);
nor U3778 (N_3778,N_2966,N_2721);
xor U3779 (N_3779,N_1815,N_2154);
xor U3780 (N_3780,N_1649,N_1690);
or U3781 (N_3781,N_2310,N_2641);
or U3782 (N_3782,N_2951,N_2932);
xor U3783 (N_3783,N_2826,N_1654);
nand U3784 (N_3784,N_2000,N_2595);
xor U3785 (N_3785,N_1626,N_2402);
and U3786 (N_3786,N_2778,N_2679);
xor U3787 (N_3787,N_2183,N_2820);
xor U3788 (N_3788,N_2953,N_2760);
nand U3789 (N_3789,N_2982,N_1579);
nand U3790 (N_3790,N_1984,N_2770);
nor U3791 (N_3791,N_2879,N_2534);
nor U3792 (N_3792,N_2440,N_2061);
and U3793 (N_3793,N_2987,N_2190);
nor U3794 (N_3794,N_1800,N_1692);
or U3795 (N_3795,N_2267,N_1636);
xor U3796 (N_3796,N_1978,N_2232);
or U3797 (N_3797,N_1647,N_1688);
or U3798 (N_3798,N_2447,N_1926);
nor U3799 (N_3799,N_2202,N_2127);
and U3800 (N_3800,N_1647,N_2325);
and U3801 (N_3801,N_2598,N_2600);
xor U3802 (N_3802,N_2862,N_2183);
nand U3803 (N_3803,N_2066,N_1771);
or U3804 (N_3804,N_2217,N_2426);
or U3805 (N_3805,N_2072,N_2840);
or U3806 (N_3806,N_1751,N_1684);
nor U3807 (N_3807,N_2439,N_2294);
xnor U3808 (N_3808,N_2000,N_2826);
nand U3809 (N_3809,N_2175,N_1628);
xor U3810 (N_3810,N_2958,N_2012);
or U3811 (N_3811,N_2517,N_2598);
and U3812 (N_3812,N_2030,N_1968);
xnor U3813 (N_3813,N_2717,N_2998);
nor U3814 (N_3814,N_2266,N_2046);
and U3815 (N_3815,N_2678,N_2388);
nor U3816 (N_3816,N_2528,N_1884);
and U3817 (N_3817,N_2595,N_2059);
xnor U3818 (N_3818,N_2896,N_2438);
and U3819 (N_3819,N_2904,N_1526);
and U3820 (N_3820,N_2230,N_2208);
and U3821 (N_3821,N_2458,N_2711);
nor U3822 (N_3822,N_2027,N_1647);
nor U3823 (N_3823,N_2371,N_2749);
or U3824 (N_3824,N_2290,N_1965);
nand U3825 (N_3825,N_2672,N_2660);
and U3826 (N_3826,N_2470,N_2112);
and U3827 (N_3827,N_1810,N_2909);
nand U3828 (N_3828,N_1903,N_1934);
nor U3829 (N_3829,N_1569,N_1860);
xnor U3830 (N_3830,N_2313,N_2160);
xnor U3831 (N_3831,N_2493,N_1548);
nand U3832 (N_3832,N_1644,N_2985);
nor U3833 (N_3833,N_2415,N_2124);
nor U3834 (N_3834,N_2511,N_1998);
nand U3835 (N_3835,N_2441,N_2291);
and U3836 (N_3836,N_1618,N_1744);
or U3837 (N_3837,N_2978,N_1973);
or U3838 (N_3838,N_2452,N_1591);
nor U3839 (N_3839,N_2751,N_2235);
or U3840 (N_3840,N_2184,N_2811);
nand U3841 (N_3841,N_1792,N_1513);
xor U3842 (N_3842,N_2853,N_1543);
or U3843 (N_3843,N_2199,N_2287);
and U3844 (N_3844,N_2475,N_1558);
nor U3845 (N_3845,N_1698,N_1754);
nor U3846 (N_3846,N_2235,N_1783);
xnor U3847 (N_3847,N_2687,N_1908);
nor U3848 (N_3848,N_2731,N_2504);
and U3849 (N_3849,N_2776,N_1880);
nand U3850 (N_3850,N_1820,N_2708);
nor U3851 (N_3851,N_2736,N_1600);
or U3852 (N_3852,N_1884,N_1833);
nand U3853 (N_3853,N_2759,N_2628);
or U3854 (N_3854,N_2481,N_2770);
nand U3855 (N_3855,N_2054,N_2557);
xor U3856 (N_3856,N_2051,N_2618);
xnor U3857 (N_3857,N_2739,N_2399);
nand U3858 (N_3858,N_2253,N_2650);
and U3859 (N_3859,N_1537,N_1701);
and U3860 (N_3860,N_2309,N_2458);
or U3861 (N_3861,N_1951,N_2994);
nand U3862 (N_3862,N_2301,N_1957);
nand U3863 (N_3863,N_2894,N_2673);
nor U3864 (N_3864,N_2426,N_2889);
and U3865 (N_3865,N_1941,N_2297);
and U3866 (N_3866,N_2887,N_1522);
nand U3867 (N_3867,N_1724,N_1911);
nor U3868 (N_3868,N_1830,N_1621);
xnor U3869 (N_3869,N_2545,N_2573);
nor U3870 (N_3870,N_1933,N_2687);
and U3871 (N_3871,N_2884,N_2725);
and U3872 (N_3872,N_1683,N_2011);
xnor U3873 (N_3873,N_2882,N_1950);
or U3874 (N_3874,N_2096,N_1526);
and U3875 (N_3875,N_2009,N_2778);
and U3876 (N_3876,N_2105,N_2229);
nor U3877 (N_3877,N_1994,N_2541);
nand U3878 (N_3878,N_1757,N_1924);
xor U3879 (N_3879,N_2885,N_1503);
or U3880 (N_3880,N_2713,N_2530);
xor U3881 (N_3881,N_2021,N_1936);
xor U3882 (N_3882,N_2034,N_2542);
and U3883 (N_3883,N_2320,N_1503);
nor U3884 (N_3884,N_2086,N_2157);
nor U3885 (N_3885,N_2288,N_2926);
nor U3886 (N_3886,N_2789,N_1744);
nor U3887 (N_3887,N_1595,N_2208);
nand U3888 (N_3888,N_2539,N_1847);
or U3889 (N_3889,N_1636,N_2901);
nor U3890 (N_3890,N_2083,N_1565);
and U3891 (N_3891,N_1621,N_2491);
xor U3892 (N_3892,N_2618,N_2293);
nand U3893 (N_3893,N_2083,N_2854);
xor U3894 (N_3894,N_2616,N_2075);
nand U3895 (N_3895,N_2833,N_1852);
and U3896 (N_3896,N_1942,N_1570);
nor U3897 (N_3897,N_2942,N_1725);
nor U3898 (N_3898,N_2557,N_2646);
or U3899 (N_3899,N_2902,N_2539);
and U3900 (N_3900,N_2394,N_1704);
nand U3901 (N_3901,N_1892,N_2727);
and U3902 (N_3902,N_2519,N_2085);
and U3903 (N_3903,N_2127,N_2041);
or U3904 (N_3904,N_1859,N_1949);
nand U3905 (N_3905,N_1937,N_2881);
or U3906 (N_3906,N_2203,N_2359);
or U3907 (N_3907,N_2529,N_2644);
nand U3908 (N_3908,N_2062,N_2384);
or U3909 (N_3909,N_2391,N_2789);
and U3910 (N_3910,N_2016,N_2919);
and U3911 (N_3911,N_1953,N_2538);
nand U3912 (N_3912,N_2369,N_1806);
nand U3913 (N_3913,N_1545,N_1888);
xor U3914 (N_3914,N_2050,N_2428);
xor U3915 (N_3915,N_2882,N_1843);
nor U3916 (N_3916,N_2634,N_1942);
nand U3917 (N_3917,N_2618,N_2291);
or U3918 (N_3918,N_1612,N_2938);
xor U3919 (N_3919,N_2561,N_2478);
or U3920 (N_3920,N_1954,N_1593);
or U3921 (N_3921,N_1966,N_2480);
nor U3922 (N_3922,N_1890,N_2630);
and U3923 (N_3923,N_1535,N_1896);
nand U3924 (N_3924,N_2129,N_2535);
or U3925 (N_3925,N_2019,N_2362);
nor U3926 (N_3926,N_2588,N_1501);
xor U3927 (N_3927,N_2297,N_2340);
and U3928 (N_3928,N_2525,N_2071);
nand U3929 (N_3929,N_2175,N_2052);
nand U3930 (N_3930,N_2898,N_2847);
xnor U3931 (N_3931,N_2725,N_2830);
and U3932 (N_3932,N_1547,N_2908);
and U3933 (N_3933,N_1693,N_2401);
or U3934 (N_3934,N_2876,N_1987);
nand U3935 (N_3935,N_1618,N_2293);
nor U3936 (N_3936,N_2805,N_2064);
xor U3937 (N_3937,N_2085,N_1591);
nor U3938 (N_3938,N_1700,N_2841);
nor U3939 (N_3939,N_2416,N_2079);
nor U3940 (N_3940,N_1901,N_2167);
and U3941 (N_3941,N_2653,N_1801);
and U3942 (N_3942,N_1567,N_2990);
xor U3943 (N_3943,N_2220,N_1645);
and U3944 (N_3944,N_2803,N_2864);
xnor U3945 (N_3945,N_2193,N_2651);
nor U3946 (N_3946,N_2989,N_2615);
and U3947 (N_3947,N_1604,N_2266);
nor U3948 (N_3948,N_1610,N_2628);
nor U3949 (N_3949,N_2580,N_1625);
and U3950 (N_3950,N_2661,N_1603);
nand U3951 (N_3951,N_2041,N_2787);
xnor U3952 (N_3952,N_2652,N_2470);
and U3953 (N_3953,N_2150,N_2894);
or U3954 (N_3954,N_2047,N_2217);
nor U3955 (N_3955,N_2667,N_1995);
nor U3956 (N_3956,N_2135,N_2166);
nand U3957 (N_3957,N_2600,N_2324);
nor U3958 (N_3958,N_2627,N_2952);
and U3959 (N_3959,N_2470,N_1708);
and U3960 (N_3960,N_1894,N_2247);
nand U3961 (N_3961,N_2296,N_2542);
xor U3962 (N_3962,N_2909,N_2678);
or U3963 (N_3963,N_2051,N_2314);
nand U3964 (N_3964,N_2316,N_1916);
xor U3965 (N_3965,N_2825,N_2186);
nor U3966 (N_3966,N_2677,N_2718);
nor U3967 (N_3967,N_1819,N_2490);
nor U3968 (N_3968,N_1786,N_2540);
nand U3969 (N_3969,N_2112,N_2236);
xnor U3970 (N_3970,N_2437,N_2980);
nor U3971 (N_3971,N_2096,N_2386);
xnor U3972 (N_3972,N_2829,N_2917);
nand U3973 (N_3973,N_2988,N_2275);
or U3974 (N_3974,N_2062,N_1668);
xnor U3975 (N_3975,N_2261,N_1930);
nand U3976 (N_3976,N_2024,N_2994);
and U3977 (N_3977,N_1665,N_2333);
nand U3978 (N_3978,N_1655,N_2573);
nand U3979 (N_3979,N_1667,N_1556);
and U3980 (N_3980,N_2315,N_1716);
nor U3981 (N_3981,N_2345,N_2459);
nor U3982 (N_3982,N_2953,N_2449);
xor U3983 (N_3983,N_2762,N_2310);
and U3984 (N_3984,N_2494,N_2709);
nand U3985 (N_3985,N_1765,N_2476);
xor U3986 (N_3986,N_2476,N_2642);
and U3987 (N_3987,N_2800,N_2594);
xor U3988 (N_3988,N_1865,N_2581);
nor U3989 (N_3989,N_2103,N_1929);
or U3990 (N_3990,N_2346,N_2851);
and U3991 (N_3991,N_1726,N_2915);
nor U3992 (N_3992,N_2654,N_2817);
nand U3993 (N_3993,N_1885,N_1635);
xor U3994 (N_3994,N_2449,N_1805);
or U3995 (N_3995,N_1971,N_2722);
and U3996 (N_3996,N_1835,N_1931);
and U3997 (N_3997,N_2931,N_1686);
or U3998 (N_3998,N_2602,N_1524);
xnor U3999 (N_3999,N_1698,N_1857);
and U4000 (N_4000,N_1675,N_1581);
xor U4001 (N_4001,N_1891,N_1649);
nand U4002 (N_4002,N_2433,N_2605);
nand U4003 (N_4003,N_2234,N_2820);
or U4004 (N_4004,N_2923,N_2914);
xnor U4005 (N_4005,N_1742,N_2953);
or U4006 (N_4006,N_1615,N_2383);
nor U4007 (N_4007,N_2587,N_2462);
or U4008 (N_4008,N_2706,N_2896);
xnor U4009 (N_4009,N_2890,N_2078);
and U4010 (N_4010,N_2862,N_2424);
or U4011 (N_4011,N_2547,N_1750);
and U4012 (N_4012,N_2336,N_2029);
nor U4013 (N_4013,N_1517,N_1651);
xnor U4014 (N_4014,N_2867,N_2028);
or U4015 (N_4015,N_2123,N_2189);
nor U4016 (N_4016,N_1560,N_2392);
and U4017 (N_4017,N_2903,N_1939);
and U4018 (N_4018,N_1543,N_2671);
xor U4019 (N_4019,N_2237,N_2794);
nand U4020 (N_4020,N_2248,N_1851);
nand U4021 (N_4021,N_1693,N_2482);
or U4022 (N_4022,N_2603,N_2703);
or U4023 (N_4023,N_2264,N_1986);
and U4024 (N_4024,N_2787,N_2684);
nand U4025 (N_4025,N_2932,N_2623);
xnor U4026 (N_4026,N_2846,N_1746);
or U4027 (N_4027,N_2531,N_1568);
and U4028 (N_4028,N_2650,N_2282);
nor U4029 (N_4029,N_1896,N_2431);
or U4030 (N_4030,N_2282,N_1821);
or U4031 (N_4031,N_2145,N_1838);
or U4032 (N_4032,N_1988,N_1621);
nor U4033 (N_4033,N_2084,N_2223);
or U4034 (N_4034,N_2700,N_1748);
or U4035 (N_4035,N_1826,N_2969);
nor U4036 (N_4036,N_2302,N_2856);
xnor U4037 (N_4037,N_2345,N_2386);
nand U4038 (N_4038,N_2185,N_2242);
nor U4039 (N_4039,N_1945,N_1974);
or U4040 (N_4040,N_2436,N_1784);
nor U4041 (N_4041,N_1835,N_2380);
nor U4042 (N_4042,N_2852,N_1975);
nor U4043 (N_4043,N_2031,N_2802);
or U4044 (N_4044,N_2835,N_2713);
and U4045 (N_4045,N_2505,N_2438);
nor U4046 (N_4046,N_2098,N_2647);
xor U4047 (N_4047,N_1572,N_1980);
nand U4048 (N_4048,N_1848,N_2301);
nor U4049 (N_4049,N_2504,N_2263);
xnor U4050 (N_4050,N_1579,N_1597);
and U4051 (N_4051,N_1581,N_1668);
xor U4052 (N_4052,N_2108,N_1937);
nor U4053 (N_4053,N_1613,N_2794);
and U4054 (N_4054,N_2668,N_1626);
and U4055 (N_4055,N_2993,N_2262);
nor U4056 (N_4056,N_2274,N_1992);
or U4057 (N_4057,N_2413,N_2952);
nor U4058 (N_4058,N_2606,N_2429);
nand U4059 (N_4059,N_1698,N_1944);
nand U4060 (N_4060,N_1808,N_1626);
or U4061 (N_4061,N_2593,N_2185);
nor U4062 (N_4062,N_2472,N_2267);
nor U4063 (N_4063,N_2452,N_2746);
and U4064 (N_4064,N_1834,N_1530);
nor U4065 (N_4065,N_2201,N_2805);
nand U4066 (N_4066,N_1561,N_2151);
or U4067 (N_4067,N_1957,N_2102);
xnor U4068 (N_4068,N_1973,N_1901);
xnor U4069 (N_4069,N_1584,N_2441);
or U4070 (N_4070,N_2891,N_2424);
or U4071 (N_4071,N_2470,N_2376);
and U4072 (N_4072,N_2080,N_1900);
nand U4073 (N_4073,N_2122,N_2907);
xnor U4074 (N_4074,N_2637,N_1957);
nor U4075 (N_4075,N_2317,N_1966);
nand U4076 (N_4076,N_2895,N_2163);
xor U4077 (N_4077,N_2097,N_2352);
and U4078 (N_4078,N_2810,N_2027);
nand U4079 (N_4079,N_2005,N_2029);
and U4080 (N_4080,N_1673,N_2046);
and U4081 (N_4081,N_1782,N_2537);
nor U4082 (N_4082,N_1762,N_2717);
or U4083 (N_4083,N_2134,N_2275);
xor U4084 (N_4084,N_1832,N_2391);
and U4085 (N_4085,N_2975,N_2941);
nor U4086 (N_4086,N_2669,N_2989);
and U4087 (N_4087,N_1985,N_2037);
nor U4088 (N_4088,N_2908,N_2058);
nor U4089 (N_4089,N_2476,N_2721);
nor U4090 (N_4090,N_2049,N_2904);
nor U4091 (N_4091,N_2048,N_1707);
or U4092 (N_4092,N_2455,N_2038);
and U4093 (N_4093,N_1989,N_2534);
and U4094 (N_4094,N_2686,N_2801);
xor U4095 (N_4095,N_1749,N_2165);
xnor U4096 (N_4096,N_2192,N_2479);
and U4097 (N_4097,N_1609,N_1512);
xor U4098 (N_4098,N_2826,N_2047);
nand U4099 (N_4099,N_1685,N_1882);
and U4100 (N_4100,N_1686,N_1506);
nor U4101 (N_4101,N_1701,N_2015);
or U4102 (N_4102,N_2582,N_2067);
nand U4103 (N_4103,N_2602,N_1648);
nand U4104 (N_4104,N_1650,N_1530);
nor U4105 (N_4105,N_2198,N_2675);
and U4106 (N_4106,N_2395,N_2733);
xnor U4107 (N_4107,N_2450,N_1856);
nor U4108 (N_4108,N_2577,N_2021);
and U4109 (N_4109,N_2233,N_1736);
or U4110 (N_4110,N_1839,N_2099);
xor U4111 (N_4111,N_2630,N_2401);
nor U4112 (N_4112,N_2013,N_1745);
xor U4113 (N_4113,N_1919,N_2521);
and U4114 (N_4114,N_2913,N_1712);
nor U4115 (N_4115,N_2273,N_2325);
xor U4116 (N_4116,N_2784,N_2810);
nand U4117 (N_4117,N_2207,N_2219);
nand U4118 (N_4118,N_1726,N_1600);
or U4119 (N_4119,N_1771,N_2592);
nor U4120 (N_4120,N_2295,N_2006);
xor U4121 (N_4121,N_2499,N_1696);
nor U4122 (N_4122,N_2416,N_2838);
nand U4123 (N_4123,N_2605,N_1882);
xor U4124 (N_4124,N_2770,N_2714);
or U4125 (N_4125,N_2934,N_2519);
or U4126 (N_4126,N_2618,N_2328);
nor U4127 (N_4127,N_2390,N_2575);
or U4128 (N_4128,N_2148,N_1797);
nand U4129 (N_4129,N_2255,N_2108);
xor U4130 (N_4130,N_2434,N_2279);
and U4131 (N_4131,N_1657,N_2673);
nand U4132 (N_4132,N_2296,N_2809);
and U4133 (N_4133,N_2185,N_1786);
xor U4134 (N_4134,N_2186,N_2328);
nor U4135 (N_4135,N_1805,N_2087);
nor U4136 (N_4136,N_2645,N_1855);
and U4137 (N_4137,N_2345,N_2771);
nor U4138 (N_4138,N_2369,N_2476);
nor U4139 (N_4139,N_2206,N_2721);
or U4140 (N_4140,N_2111,N_1705);
xor U4141 (N_4141,N_1815,N_2103);
nor U4142 (N_4142,N_2249,N_1645);
or U4143 (N_4143,N_2229,N_2598);
or U4144 (N_4144,N_1516,N_2202);
xnor U4145 (N_4145,N_1875,N_2793);
nand U4146 (N_4146,N_1516,N_1518);
nor U4147 (N_4147,N_1931,N_2273);
nor U4148 (N_4148,N_2659,N_2867);
and U4149 (N_4149,N_2004,N_2597);
xor U4150 (N_4150,N_2680,N_2127);
and U4151 (N_4151,N_2943,N_1531);
or U4152 (N_4152,N_2246,N_1809);
or U4153 (N_4153,N_2469,N_2568);
nor U4154 (N_4154,N_1591,N_2686);
and U4155 (N_4155,N_2449,N_1648);
nand U4156 (N_4156,N_2949,N_1811);
xnor U4157 (N_4157,N_2998,N_2577);
nand U4158 (N_4158,N_1914,N_2350);
xnor U4159 (N_4159,N_1818,N_2791);
and U4160 (N_4160,N_2199,N_2280);
nor U4161 (N_4161,N_2345,N_2614);
xnor U4162 (N_4162,N_1676,N_2527);
nor U4163 (N_4163,N_2019,N_2015);
nand U4164 (N_4164,N_2652,N_2034);
nand U4165 (N_4165,N_1883,N_2195);
nor U4166 (N_4166,N_2613,N_1751);
xnor U4167 (N_4167,N_2136,N_2056);
xnor U4168 (N_4168,N_1635,N_2322);
nand U4169 (N_4169,N_1792,N_1681);
xnor U4170 (N_4170,N_1686,N_2709);
or U4171 (N_4171,N_1633,N_2709);
nand U4172 (N_4172,N_2364,N_1805);
nor U4173 (N_4173,N_1510,N_2795);
or U4174 (N_4174,N_2477,N_2033);
nand U4175 (N_4175,N_2306,N_2148);
nor U4176 (N_4176,N_1748,N_2201);
and U4177 (N_4177,N_2358,N_1705);
xnor U4178 (N_4178,N_1947,N_2172);
nor U4179 (N_4179,N_2073,N_2962);
and U4180 (N_4180,N_2613,N_2220);
nand U4181 (N_4181,N_2494,N_2623);
nand U4182 (N_4182,N_1574,N_1780);
xor U4183 (N_4183,N_1970,N_2222);
nand U4184 (N_4184,N_2580,N_2576);
or U4185 (N_4185,N_2021,N_1692);
xor U4186 (N_4186,N_2593,N_2845);
and U4187 (N_4187,N_2638,N_2374);
or U4188 (N_4188,N_2456,N_2707);
nand U4189 (N_4189,N_2447,N_2270);
nand U4190 (N_4190,N_2191,N_2528);
nor U4191 (N_4191,N_2826,N_2983);
xnor U4192 (N_4192,N_1594,N_2654);
nand U4193 (N_4193,N_2919,N_1850);
xor U4194 (N_4194,N_2479,N_2787);
or U4195 (N_4195,N_1824,N_2117);
nor U4196 (N_4196,N_1982,N_2111);
nand U4197 (N_4197,N_2443,N_2708);
and U4198 (N_4198,N_2334,N_2242);
xnor U4199 (N_4199,N_1536,N_2434);
nand U4200 (N_4200,N_2756,N_1981);
nand U4201 (N_4201,N_2931,N_2721);
nand U4202 (N_4202,N_1501,N_2289);
nand U4203 (N_4203,N_2655,N_2475);
xnor U4204 (N_4204,N_1768,N_1755);
or U4205 (N_4205,N_2242,N_2603);
xnor U4206 (N_4206,N_2225,N_1645);
and U4207 (N_4207,N_2337,N_2978);
xnor U4208 (N_4208,N_1698,N_2563);
xor U4209 (N_4209,N_2671,N_2298);
and U4210 (N_4210,N_2703,N_2960);
xnor U4211 (N_4211,N_2496,N_2257);
and U4212 (N_4212,N_2739,N_2140);
nor U4213 (N_4213,N_1527,N_2921);
nand U4214 (N_4214,N_2084,N_2506);
nor U4215 (N_4215,N_2383,N_2003);
nor U4216 (N_4216,N_2219,N_2173);
or U4217 (N_4217,N_1608,N_2349);
nand U4218 (N_4218,N_2078,N_2314);
or U4219 (N_4219,N_1907,N_2176);
nand U4220 (N_4220,N_2808,N_2076);
or U4221 (N_4221,N_2522,N_2258);
nor U4222 (N_4222,N_2784,N_2428);
and U4223 (N_4223,N_2545,N_2290);
or U4224 (N_4224,N_1769,N_1699);
nor U4225 (N_4225,N_1740,N_2685);
and U4226 (N_4226,N_2952,N_2526);
xnor U4227 (N_4227,N_1850,N_2633);
nand U4228 (N_4228,N_1963,N_1612);
or U4229 (N_4229,N_2384,N_2130);
and U4230 (N_4230,N_1838,N_2588);
and U4231 (N_4231,N_2463,N_1831);
or U4232 (N_4232,N_2590,N_1980);
nor U4233 (N_4233,N_2546,N_1610);
or U4234 (N_4234,N_2445,N_1619);
nand U4235 (N_4235,N_2368,N_2863);
nor U4236 (N_4236,N_1624,N_2691);
nand U4237 (N_4237,N_2398,N_2793);
nor U4238 (N_4238,N_2122,N_2310);
nand U4239 (N_4239,N_2488,N_1617);
or U4240 (N_4240,N_2133,N_2001);
xnor U4241 (N_4241,N_2380,N_1568);
nand U4242 (N_4242,N_2631,N_2412);
nand U4243 (N_4243,N_2466,N_2850);
or U4244 (N_4244,N_2061,N_1667);
or U4245 (N_4245,N_2409,N_2786);
or U4246 (N_4246,N_2017,N_1812);
nand U4247 (N_4247,N_1594,N_2088);
xnor U4248 (N_4248,N_2004,N_1877);
and U4249 (N_4249,N_2062,N_2736);
or U4250 (N_4250,N_2982,N_2594);
nor U4251 (N_4251,N_2662,N_2251);
nor U4252 (N_4252,N_1552,N_1955);
nor U4253 (N_4253,N_1795,N_2421);
nor U4254 (N_4254,N_1717,N_1544);
nand U4255 (N_4255,N_2704,N_1791);
xnor U4256 (N_4256,N_2069,N_1516);
or U4257 (N_4257,N_2382,N_1925);
xnor U4258 (N_4258,N_2450,N_2352);
and U4259 (N_4259,N_1901,N_2791);
or U4260 (N_4260,N_1908,N_2772);
nand U4261 (N_4261,N_2437,N_2963);
xor U4262 (N_4262,N_1536,N_2694);
xor U4263 (N_4263,N_2947,N_1573);
xor U4264 (N_4264,N_1866,N_1643);
nand U4265 (N_4265,N_2193,N_2243);
xor U4266 (N_4266,N_2335,N_1645);
xnor U4267 (N_4267,N_2253,N_1809);
nor U4268 (N_4268,N_2517,N_1744);
nor U4269 (N_4269,N_2702,N_2636);
and U4270 (N_4270,N_2379,N_2990);
nand U4271 (N_4271,N_2353,N_1839);
nand U4272 (N_4272,N_2150,N_1824);
xnor U4273 (N_4273,N_1922,N_2140);
nor U4274 (N_4274,N_1516,N_1875);
nor U4275 (N_4275,N_2965,N_2127);
or U4276 (N_4276,N_2968,N_2678);
nor U4277 (N_4277,N_1682,N_2153);
xnor U4278 (N_4278,N_2965,N_2680);
nor U4279 (N_4279,N_2866,N_2977);
xnor U4280 (N_4280,N_2276,N_2397);
or U4281 (N_4281,N_2580,N_1887);
nand U4282 (N_4282,N_2563,N_2139);
nand U4283 (N_4283,N_1976,N_1751);
or U4284 (N_4284,N_1731,N_2910);
xor U4285 (N_4285,N_2177,N_2713);
and U4286 (N_4286,N_1571,N_2629);
nor U4287 (N_4287,N_1751,N_2306);
xor U4288 (N_4288,N_2627,N_1694);
and U4289 (N_4289,N_2352,N_2548);
nor U4290 (N_4290,N_1530,N_2282);
xnor U4291 (N_4291,N_2017,N_2984);
nand U4292 (N_4292,N_2382,N_1973);
or U4293 (N_4293,N_2104,N_2188);
nand U4294 (N_4294,N_2216,N_1506);
nand U4295 (N_4295,N_2035,N_2579);
nor U4296 (N_4296,N_2822,N_2129);
and U4297 (N_4297,N_2211,N_2190);
nor U4298 (N_4298,N_2552,N_2430);
xnor U4299 (N_4299,N_1569,N_1870);
nand U4300 (N_4300,N_2076,N_2799);
nand U4301 (N_4301,N_2871,N_2066);
nor U4302 (N_4302,N_2140,N_2127);
or U4303 (N_4303,N_1940,N_2584);
nand U4304 (N_4304,N_2555,N_2147);
and U4305 (N_4305,N_1641,N_2281);
and U4306 (N_4306,N_2710,N_2532);
xnor U4307 (N_4307,N_2440,N_2313);
or U4308 (N_4308,N_2483,N_2572);
or U4309 (N_4309,N_2245,N_2974);
xnor U4310 (N_4310,N_1667,N_2350);
and U4311 (N_4311,N_1719,N_1782);
nand U4312 (N_4312,N_1705,N_2988);
nor U4313 (N_4313,N_2251,N_2431);
and U4314 (N_4314,N_2957,N_2984);
nand U4315 (N_4315,N_2001,N_2451);
and U4316 (N_4316,N_2714,N_2838);
and U4317 (N_4317,N_1872,N_2822);
or U4318 (N_4318,N_1551,N_2428);
or U4319 (N_4319,N_2881,N_1530);
nor U4320 (N_4320,N_2024,N_2288);
xor U4321 (N_4321,N_2396,N_1762);
nor U4322 (N_4322,N_2169,N_1537);
and U4323 (N_4323,N_1828,N_1769);
or U4324 (N_4324,N_1656,N_1505);
nor U4325 (N_4325,N_2859,N_2855);
or U4326 (N_4326,N_2106,N_2245);
and U4327 (N_4327,N_1642,N_1718);
or U4328 (N_4328,N_2853,N_2983);
nor U4329 (N_4329,N_2723,N_2144);
xnor U4330 (N_4330,N_2842,N_1875);
or U4331 (N_4331,N_1797,N_1528);
nor U4332 (N_4332,N_1729,N_1798);
nor U4333 (N_4333,N_2974,N_2450);
and U4334 (N_4334,N_2791,N_2667);
nor U4335 (N_4335,N_2885,N_2628);
nand U4336 (N_4336,N_2714,N_2254);
nor U4337 (N_4337,N_2695,N_2490);
and U4338 (N_4338,N_2293,N_2091);
nand U4339 (N_4339,N_2927,N_2464);
or U4340 (N_4340,N_2376,N_2327);
or U4341 (N_4341,N_2507,N_1961);
nor U4342 (N_4342,N_2709,N_2464);
and U4343 (N_4343,N_1527,N_2437);
xnor U4344 (N_4344,N_2877,N_2524);
and U4345 (N_4345,N_2963,N_2930);
nor U4346 (N_4346,N_2657,N_2670);
or U4347 (N_4347,N_2215,N_1764);
xor U4348 (N_4348,N_1505,N_2243);
nor U4349 (N_4349,N_2426,N_1798);
xor U4350 (N_4350,N_2387,N_2964);
nand U4351 (N_4351,N_2340,N_2787);
xor U4352 (N_4352,N_2485,N_2421);
xor U4353 (N_4353,N_2505,N_2408);
nor U4354 (N_4354,N_2530,N_2395);
nor U4355 (N_4355,N_2095,N_2260);
nand U4356 (N_4356,N_2456,N_2711);
or U4357 (N_4357,N_1710,N_2742);
or U4358 (N_4358,N_2320,N_2331);
xor U4359 (N_4359,N_2335,N_2355);
and U4360 (N_4360,N_2722,N_1794);
nor U4361 (N_4361,N_2401,N_1767);
xor U4362 (N_4362,N_1697,N_1553);
xnor U4363 (N_4363,N_2418,N_1528);
nor U4364 (N_4364,N_2303,N_2655);
nand U4365 (N_4365,N_1924,N_2223);
nand U4366 (N_4366,N_2802,N_1770);
nand U4367 (N_4367,N_2067,N_2721);
nor U4368 (N_4368,N_2261,N_2843);
and U4369 (N_4369,N_2233,N_2653);
xor U4370 (N_4370,N_2876,N_1905);
and U4371 (N_4371,N_2304,N_1929);
and U4372 (N_4372,N_2833,N_2165);
or U4373 (N_4373,N_1619,N_1838);
or U4374 (N_4374,N_1809,N_2072);
or U4375 (N_4375,N_1802,N_2447);
or U4376 (N_4376,N_2069,N_2540);
nor U4377 (N_4377,N_1671,N_1600);
xor U4378 (N_4378,N_1510,N_1723);
and U4379 (N_4379,N_1668,N_2597);
xnor U4380 (N_4380,N_2415,N_2110);
or U4381 (N_4381,N_2479,N_1987);
nor U4382 (N_4382,N_2247,N_2483);
nor U4383 (N_4383,N_2680,N_1597);
nand U4384 (N_4384,N_2693,N_1802);
xnor U4385 (N_4385,N_2766,N_2070);
nor U4386 (N_4386,N_2054,N_1550);
nor U4387 (N_4387,N_1715,N_2620);
and U4388 (N_4388,N_1693,N_2738);
xnor U4389 (N_4389,N_2964,N_2827);
xor U4390 (N_4390,N_2601,N_2920);
nand U4391 (N_4391,N_2768,N_2891);
and U4392 (N_4392,N_2980,N_1760);
and U4393 (N_4393,N_2684,N_2672);
nand U4394 (N_4394,N_1935,N_2053);
nor U4395 (N_4395,N_1832,N_2198);
nand U4396 (N_4396,N_2657,N_1597);
and U4397 (N_4397,N_2028,N_2638);
and U4398 (N_4398,N_2641,N_1776);
xor U4399 (N_4399,N_2972,N_2553);
xnor U4400 (N_4400,N_1672,N_1876);
xor U4401 (N_4401,N_1837,N_1517);
nor U4402 (N_4402,N_2593,N_1682);
or U4403 (N_4403,N_2634,N_1627);
nand U4404 (N_4404,N_2930,N_2658);
xor U4405 (N_4405,N_2829,N_2361);
nand U4406 (N_4406,N_1832,N_2218);
and U4407 (N_4407,N_2180,N_2613);
nand U4408 (N_4408,N_2890,N_2456);
xnor U4409 (N_4409,N_1658,N_1988);
xor U4410 (N_4410,N_2334,N_1778);
nor U4411 (N_4411,N_1542,N_2304);
xor U4412 (N_4412,N_2556,N_2373);
xnor U4413 (N_4413,N_2132,N_2238);
nor U4414 (N_4414,N_1879,N_2404);
nor U4415 (N_4415,N_2800,N_2324);
nand U4416 (N_4416,N_1869,N_2901);
or U4417 (N_4417,N_1779,N_1564);
xor U4418 (N_4418,N_1912,N_2945);
or U4419 (N_4419,N_2318,N_2145);
nand U4420 (N_4420,N_1967,N_2385);
nor U4421 (N_4421,N_2030,N_1604);
xor U4422 (N_4422,N_2948,N_2257);
xnor U4423 (N_4423,N_2254,N_1914);
and U4424 (N_4424,N_2594,N_2556);
nand U4425 (N_4425,N_1943,N_2514);
nor U4426 (N_4426,N_2077,N_2414);
nand U4427 (N_4427,N_1815,N_2986);
and U4428 (N_4428,N_1862,N_1943);
and U4429 (N_4429,N_1636,N_1846);
xnor U4430 (N_4430,N_1679,N_2575);
or U4431 (N_4431,N_1992,N_1681);
xor U4432 (N_4432,N_2448,N_2527);
nand U4433 (N_4433,N_2412,N_1511);
nand U4434 (N_4434,N_1697,N_2549);
or U4435 (N_4435,N_2918,N_2056);
xnor U4436 (N_4436,N_2812,N_1533);
and U4437 (N_4437,N_2138,N_2185);
and U4438 (N_4438,N_2630,N_2559);
and U4439 (N_4439,N_2169,N_1721);
or U4440 (N_4440,N_1672,N_2592);
or U4441 (N_4441,N_2769,N_2665);
or U4442 (N_4442,N_1543,N_2858);
or U4443 (N_4443,N_2912,N_2479);
nand U4444 (N_4444,N_2291,N_2123);
or U4445 (N_4445,N_2048,N_2373);
or U4446 (N_4446,N_2336,N_2267);
or U4447 (N_4447,N_2057,N_2548);
nor U4448 (N_4448,N_1889,N_1854);
or U4449 (N_4449,N_2638,N_1807);
and U4450 (N_4450,N_2068,N_2871);
or U4451 (N_4451,N_2344,N_1565);
nor U4452 (N_4452,N_1643,N_1993);
nor U4453 (N_4453,N_1700,N_2612);
and U4454 (N_4454,N_2310,N_2550);
and U4455 (N_4455,N_2730,N_1825);
xnor U4456 (N_4456,N_2538,N_2136);
nor U4457 (N_4457,N_2189,N_2520);
and U4458 (N_4458,N_1973,N_2264);
nor U4459 (N_4459,N_2969,N_1619);
nor U4460 (N_4460,N_2441,N_2423);
nand U4461 (N_4461,N_2981,N_1868);
nor U4462 (N_4462,N_2807,N_2398);
or U4463 (N_4463,N_2043,N_1865);
nor U4464 (N_4464,N_2657,N_1814);
and U4465 (N_4465,N_2927,N_2186);
nand U4466 (N_4466,N_2833,N_2301);
nand U4467 (N_4467,N_2025,N_1527);
nand U4468 (N_4468,N_2383,N_1556);
and U4469 (N_4469,N_2207,N_2469);
nand U4470 (N_4470,N_2132,N_1748);
and U4471 (N_4471,N_2082,N_1714);
nor U4472 (N_4472,N_2135,N_2971);
xor U4473 (N_4473,N_2246,N_1871);
xnor U4474 (N_4474,N_2166,N_2245);
xnor U4475 (N_4475,N_2487,N_2564);
nor U4476 (N_4476,N_2419,N_2508);
or U4477 (N_4477,N_2904,N_2378);
xnor U4478 (N_4478,N_2110,N_1712);
nand U4479 (N_4479,N_2583,N_1926);
and U4480 (N_4480,N_2713,N_1875);
or U4481 (N_4481,N_2223,N_2818);
nand U4482 (N_4482,N_2498,N_2762);
xor U4483 (N_4483,N_2433,N_1856);
and U4484 (N_4484,N_2233,N_2370);
nand U4485 (N_4485,N_2696,N_2561);
or U4486 (N_4486,N_2599,N_1713);
nor U4487 (N_4487,N_2431,N_2642);
or U4488 (N_4488,N_2623,N_2937);
xor U4489 (N_4489,N_1959,N_2644);
nor U4490 (N_4490,N_1612,N_2014);
nor U4491 (N_4491,N_2361,N_2634);
nand U4492 (N_4492,N_2177,N_2183);
nand U4493 (N_4493,N_2339,N_1843);
and U4494 (N_4494,N_2042,N_1893);
nand U4495 (N_4495,N_2443,N_1579);
nand U4496 (N_4496,N_1819,N_2719);
or U4497 (N_4497,N_1959,N_2974);
xor U4498 (N_4498,N_1966,N_1766);
xor U4499 (N_4499,N_1981,N_2289);
nand U4500 (N_4500,N_3632,N_4436);
and U4501 (N_4501,N_4057,N_3471);
or U4502 (N_4502,N_3678,N_3092);
and U4503 (N_4503,N_3435,N_3715);
or U4504 (N_4504,N_3111,N_4273);
and U4505 (N_4505,N_3407,N_3008);
nand U4506 (N_4506,N_3874,N_4482);
nor U4507 (N_4507,N_3935,N_3699);
nor U4508 (N_4508,N_4055,N_4022);
nand U4509 (N_4509,N_3677,N_4212);
nand U4510 (N_4510,N_3709,N_3021);
and U4511 (N_4511,N_4362,N_3266);
nand U4512 (N_4512,N_3304,N_4002);
nor U4513 (N_4513,N_3548,N_3576);
and U4514 (N_4514,N_3805,N_3164);
nand U4515 (N_4515,N_4082,N_3762);
nor U4516 (N_4516,N_3364,N_4007);
and U4517 (N_4517,N_4173,N_4324);
nand U4518 (N_4518,N_3898,N_3983);
xnor U4519 (N_4519,N_4448,N_3116);
and U4520 (N_4520,N_3769,N_3726);
or U4521 (N_4521,N_3568,N_3071);
nand U4522 (N_4522,N_3032,N_3154);
and U4523 (N_4523,N_3968,N_3792);
xnor U4524 (N_4524,N_4117,N_3251);
nor U4525 (N_4525,N_3499,N_3084);
and U4526 (N_4526,N_3401,N_3245);
and U4527 (N_4527,N_4187,N_3205);
and U4528 (N_4528,N_3518,N_3775);
nand U4529 (N_4529,N_4365,N_4064);
nand U4530 (N_4530,N_3979,N_4041);
xnor U4531 (N_4531,N_3423,N_3190);
nand U4532 (N_4532,N_3146,N_3460);
or U4533 (N_4533,N_3652,N_4167);
nand U4534 (N_4534,N_3836,N_3505);
nor U4535 (N_4535,N_3105,N_4428);
xor U4536 (N_4536,N_3734,N_3155);
nor U4537 (N_4537,N_3786,N_3733);
or U4538 (N_4538,N_3274,N_3090);
and U4539 (N_4539,N_4455,N_3227);
xnor U4540 (N_4540,N_4164,N_3130);
nand U4541 (N_4541,N_3224,N_3450);
xnor U4542 (N_4542,N_4244,N_3177);
nor U4543 (N_4543,N_4315,N_3627);
xor U4544 (N_4544,N_4264,N_3840);
nand U4545 (N_4545,N_4462,N_3741);
nand U4546 (N_4546,N_4447,N_3540);
nor U4547 (N_4547,N_3419,N_3270);
nor U4548 (N_4548,N_3911,N_4274);
nand U4549 (N_4549,N_3322,N_4368);
and U4550 (N_4550,N_4354,N_3700);
and U4551 (N_4551,N_4397,N_4377);
nand U4552 (N_4552,N_3140,N_4165);
nand U4553 (N_4553,N_4336,N_3943);
nand U4554 (N_4554,N_3358,N_4032);
xnor U4555 (N_4555,N_4018,N_3153);
nor U4556 (N_4556,N_3987,N_3914);
nor U4557 (N_4557,N_3318,N_4459);
or U4558 (N_4558,N_3226,N_4139);
nor U4559 (N_4559,N_3168,N_3504);
xor U4560 (N_4560,N_3239,N_3844);
nand U4561 (N_4561,N_4169,N_3664);
or U4562 (N_4562,N_3004,N_4160);
and U4563 (N_4563,N_3575,N_4246);
nand U4564 (N_4564,N_3309,N_3927);
and U4565 (N_4565,N_3708,N_3737);
xnor U4566 (N_4566,N_3779,N_4060);
and U4567 (N_4567,N_3108,N_3661);
nand U4568 (N_4568,N_3824,N_3254);
nor U4569 (N_4569,N_3740,N_3767);
or U4570 (N_4570,N_3656,N_3856);
xor U4571 (N_4571,N_3372,N_3657);
and U4572 (N_4572,N_3170,N_3222);
or U4573 (N_4573,N_3075,N_4218);
nand U4574 (N_4574,N_3392,N_3379);
or U4575 (N_4575,N_3683,N_3049);
or U4576 (N_4576,N_3875,N_4297);
or U4577 (N_4577,N_4090,N_4402);
and U4578 (N_4578,N_4488,N_4376);
xor U4579 (N_4579,N_3953,N_3204);
and U4580 (N_4580,N_3705,N_3511);
nand U4581 (N_4581,N_3044,N_3563);
nand U4582 (N_4582,N_3917,N_4069);
and U4583 (N_4583,N_4296,N_3897);
and U4584 (N_4584,N_3022,N_4314);
xnor U4585 (N_4585,N_3999,N_4446);
or U4586 (N_4586,N_3790,N_4312);
nand U4587 (N_4587,N_3633,N_3973);
or U4588 (N_4588,N_3565,N_3408);
nor U4589 (N_4589,N_3234,N_4471);
nand U4590 (N_4590,N_3711,N_4494);
nor U4591 (N_4591,N_3113,N_4284);
and U4592 (N_4592,N_3115,N_4190);
or U4593 (N_4593,N_3112,N_3502);
nor U4594 (N_4594,N_4370,N_3820);
or U4595 (N_4595,N_3959,N_3232);
nor U4596 (N_4596,N_3131,N_3742);
nor U4597 (N_4597,N_3217,N_3040);
nor U4598 (N_4598,N_3888,N_3469);
xor U4599 (N_4599,N_4414,N_3919);
xor U4600 (N_4600,N_3553,N_4299);
and U4601 (N_4601,N_3595,N_3949);
and U4602 (N_4602,N_4341,N_4182);
xnor U4603 (N_4603,N_3373,N_3206);
and U4604 (N_4604,N_4205,N_4305);
nand U4605 (N_4605,N_3102,N_4150);
or U4606 (N_4606,N_3926,N_3852);
and U4607 (N_4607,N_3387,N_3745);
nand U4608 (N_4608,N_3298,N_4313);
or U4609 (N_4609,N_3476,N_3203);
xnor U4610 (N_4610,N_3730,N_4036);
and U4611 (N_4611,N_4476,N_4356);
xor U4612 (N_4612,N_3583,N_4398);
nor U4613 (N_4613,N_4159,N_3359);
nand U4614 (N_4614,N_3864,N_3581);
nand U4615 (N_4615,N_4326,N_3931);
and U4616 (N_4616,N_3380,N_3489);
nor U4617 (N_4617,N_3910,N_3908);
nand U4618 (N_4618,N_3724,N_3213);
or U4619 (N_4619,N_3671,N_3334);
or U4620 (N_4620,N_3448,N_3037);
or U4621 (N_4621,N_3057,N_3808);
or U4622 (N_4622,N_3451,N_4088);
nand U4623 (N_4623,N_3339,N_3967);
and U4624 (N_4624,N_4390,N_4434);
nor U4625 (N_4625,N_3244,N_3788);
and U4626 (N_4626,N_3971,N_4175);
and U4627 (N_4627,N_3867,N_3582);
or U4628 (N_4628,N_3912,N_3252);
and U4629 (N_4629,N_4110,N_3552);
or U4630 (N_4630,N_3473,N_3682);
nand U4631 (N_4631,N_3366,N_4113);
xor U4632 (N_4632,N_3296,N_3142);
nor U4633 (N_4633,N_3596,N_4497);
nand U4634 (N_4634,N_3370,N_3617);
xnor U4635 (N_4635,N_3857,N_3795);
and U4636 (N_4636,N_4387,N_3027);
xor U4637 (N_4637,N_3615,N_3028);
xor U4638 (N_4638,N_3849,N_3486);
or U4639 (N_4639,N_4358,N_3600);
or U4640 (N_4640,N_3727,N_3761);
nand U4641 (N_4641,N_3332,N_4413);
nand U4642 (N_4642,N_4388,N_3295);
and U4643 (N_4643,N_4158,N_3965);
nand U4644 (N_4644,N_3637,N_3909);
nand U4645 (N_4645,N_4236,N_3942);
nor U4646 (N_4646,N_3011,N_3586);
or U4647 (N_4647,N_3316,N_4003);
and U4648 (N_4648,N_4043,N_3340);
or U4649 (N_4649,N_3995,N_3496);
and U4650 (N_4650,N_3345,N_3353);
or U4651 (N_4651,N_3194,N_3530);
nor U4652 (N_4652,N_3058,N_4039);
and U4653 (N_4653,N_4066,N_4340);
xnor U4654 (N_4654,N_4103,N_3900);
and U4655 (N_4655,N_3346,N_4411);
xor U4656 (N_4656,N_4058,N_4225);
nor U4657 (N_4657,N_3438,N_3033);
nor U4658 (N_4658,N_4149,N_4347);
xnor U4659 (N_4659,N_3845,N_3242);
nor U4660 (N_4660,N_4319,N_3030);
or U4661 (N_4661,N_3992,N_3892);
or U4662 (N_4662,N_3443,N_4063);
nor U4663 (N_4663,N_3760,N_3421);
and U4664 (N_4664,N_3713,N_3798);
nand U4665 (N_4665,N_3587,N_3466);
nand U4666 (N_4666,N_4485,N_3822);
and U4667 (N_4667,N_3570,N_3406);
nor U4668 (N_4668,N_3123,N_3034);
xnor U4669 (N_4669,N_3237,N_4374);
nand U4670 (N_4670,N_4238,N_3261);
nand U4671 (N_4671,N_4230,N_3644);
nor U4672 (N_4672,N_3389,N_3097);
and U4673 (N_4673,N_4210,N_4479);
nand U4674 (N_4674,N_3147,N_3431);
nand U4675 (N_4675,N_4138,N_4412);
nand U4676 (N_4676,N_3026,N_4227);
xnor U4677 (N_4677,N_3143,N_3765);
and U4678 (N_4678,N_3870,N_3378);
nor U4679 (N_4679,N_4237,N_4251);
nand U4680 (N_4680,N_3879,N_3646);
nand U4681 (N_4681,N_4067,N_3161);
and U4682 (N_4682,N_3225,N_3126);
and U4683 (N_4683,N_4292,N_4287);
xnor U4684 (N_4684,N_3286,N_3262);
nor U4685 (N_4685,N_3197,N_4247);
and U4686 (N_4686,N_3209,N_3179);
xnor U4687 (N_4687,N_3236,N_3602);
or U4688 (N_4688,N_3738,N_3667);
nor U4689 (N_4689,N_4048,N_3104);
or U4690 (N_4690,N_3488,N_4013);
or U4691 (N_4691,N_3002,N_4140);
xnor U4692 (N_4692,N_3273,N_4091);
xor U4693 (N_4693,N_4381,N_4062);
and U4694 (N_4694,N_4100,N_3235);
xor U4695 (N_4695,N_4391,N_3208);
or U4696 (N_4696,N_4081,N_3827);
xnor U4697 (N_4697,N_3982,N_4196);
xor U4698 (N_4698,N_3106,N_3806);
nor U4699 (N_4699,N_4176,N_4047);
nand U4700 (N_4700,N_3085,N_4440);
nand U4701 (N_4701,N_3706,N_4404);
or U4702 (N_4702,N_3970,N_3484);
or U4703 (N_4703,N_3220,N_3704);
xnor U4704 (N_4704,N_4318,N_3079);
nor U4705 (N_4705,N_3182,N_3783);
and U4706 (N_4706,N_3279,N_3925);
xor U4707 (N_4707,N_3804,N_3409);
nand U4708 (N_4708,N_4243,N_4144);
and U4709 (N_4709,N_3754,N_3117);
xnor U4710 (N_4710,N_3559,N_3189);
nand U4711 (N_4711,N_3305,N_3752);
and U4712 (N_4712,N_3394,N_3173);
or U4713 (N_4713,N_3422,N_3088);
or U4714 (N_4714,N_3437,N_4033);
nor U4715 (N_4715,N_4372,N_4277);
and U4716 (N_4716,N_3230,N_3495);
xnor U4717 (N_4717,N_3690,N_3152);
nand U4718 (N_4718,N_4442,N_3386);
and U4719 (N_4719,N_4121,N_4141);
or U4720 (N_4720,N_3894,N_3297);
and U4721 (N_4721,N_3271,N_3756);
nor U4722 (N_4722,N_4009,N_3947);
or U4723 (N_4723,N_3969,N_3782);
and U4724 (N_4724,N_3639,N_3785);
or U4725 (N_4725,N_3649,N_4118);
nand U4726 (N_4726,N_3461,N_3416);
nor U4727 (N_4727,N_3962,N_3744);
nand U4728 (N_4728,N_4094,N_4310);
nor U4729 (N_4729,N_4204,N_4153);
nand U4730 (N_4730,N_4078,N_3736);
nor U4731 (N_4731,N_4385,N_3180);
nor U4732 (N_4732,N_3751,N_3127);
or U4733 (N_4733,N_3636,N_3755);
nor U4734 (N_4734,N_4099,N_3047);
and U4735 (N_4735,N_3939,N_3513);
xor U4736 (N_4736,N_3776,N_4104);
or U4737 (N_4737,N_4122,N_4054);
or U4738 (N_4738,N_3937,N_3120);
nor U4739 (N_4739,N_3485,N_3464);
or U4740 (N_4740,N_3186,N_3089);
nand U4741 (N_4741,N_3948,N_3418);
nor U4742 (N_4742,N_3641,N_3086);
nor U4743 (N_4743,N_4386,N_3398);
xor U4744 (N_4744,N_3569,N_4481);
xnor U4745 (N_4745,N_3412,N_4294);
xnor U4746 (N_4746,N_3136,N_3915);
or U4747 (N_4747,N_4478,N_4148);
and U4748 (N_4748,N_4421,N_3543);
or U4749 (N_4749,N_4460,N_4235);
xor U4750 (N_4750,N_4426,N_3958);
and U4751 (N_4751,N_3800,N_3594);
xor U4752 (N_4752,N_3689,N_3932);
nor U4753 (N_4753,N_3536,N_3929);
and U4754 (N_4754,N_3584,N_3562);
xor U4755 (N_4755,N_3045,N_4178);
nor U4756 (N_4756,N_4226,N_3415);
xnor U4757 (N_4757,N_4267,N_3384);
xor U4758 (N_4758,N_3528,N_4030);
nor U4759 (N_4759,N_4405,N_4389);
nor U4760 (N_4760,N_3520,N_3338);
nor U4761 (N_4761,N_3149,N_3608);
or U4762 (N_4762,N_3402,N_3121);
and U4763 (N_4763,N_3355,N_3367);
nand U4764 (N_4764,N_3281,N_3472);
and U4765 (N_4765,N_4407,N_4275);
xor U4766 (N_4766,N_4320,N_4450);
xnor U4767 (N_4767,N_3467,N_3966);
and U4768 (N_4768,N_4156,N_4283);
and U4769 (N_4769,N_4219,N_3414);
xor U4770 (N_4770,N_4008,N_4157);
nand U4771 (N_4771,N_4458,N_4337);
xnor U4772 (N_4772,N_4427,N_4371);
and U4773 (N_4773,N_3626,N_3853);
xor U4774 (N_4774,N_3855,N_3643);
xor U4775 (N_4775,N_3672,N_3538);
or U4776 (N_4776,N_3803,N_3228);
xor U4777 (N_4777,N_3167,N_4461);
nand U4778 (N_4778,N_3591,N_3006);
or U4779 (N_4779,N_3201,N_3183);
and U4780 (N_4780,N_4269,N_4217);
xnor U4781 (N_4781,N_3132,N_3846);
or U4782 (N_4782,N_3895,N_3918);
nand U4783 (N_4783,N_3527,N_3439);
xnor U4784 (N_4784,N_3383,N_3986);
xor U4785 (N_4785,N_3861,N_4346);
xor U4786 (N_4786,N_3818,N_3043);
nor U4787 (N_4787,N_3145,N_3426);
xor U4788 (N_4788,N_4163,N_3374);
or U4789 (N_4789,N_3272,N_4061);
or U4790 (N_4790,N_4351,N_3507);
or U4791 (N_4791,N_3067,N_3328);
or U4792 (N_4792,N_3498,N_3425);
nand U4793 (N_4793,N_3631,N_3427);
nand U4794 (N_4794,N_4107,N_4480);
or U4795 (N_4795,N_4124,N_3860);
nor U4796 (N_4796,N_3863,N_3732);
and U4797 (N_4797,N_3753,N_4498);
and U4798 (N_4798,N_3100,N_3441);
xnor U4799 (N_4799,N_4015,N_4456);
nor U4800 (N_4800,N_3436,N_3212);
nand U4801 (N_4801,N_3887,N_4191);
and U4802 (N_4802,N_3793,N_3821);
and U4803 (N_4803,N_3980,N_4306);
nand U4804 (N_4804,N_3635,N_4215);
nand U4805 (N_4805,N_3319,N_4367);
or U4806 (N_4806,N_4396,N_3487);
nand U4807 (N_4807,N_3739,N_3302);
nor U4808 (N_4808,N_3590,N_3869);
and U4809 (N_4809,N_3264,N_3393);
xor U4810 (N_4810,N_4499,N_3198);
and U4811 (N_4811,N_4345,N_3588);
or U4812 (N_4812,N_3957,N_4184);
or U4813 (N_4813,N_3256,N_3797);
and U4814 (N_4814,N_3572,N_3963);
or U4815 (N_4815,N_4457,N_3331);
nor U4816 (N_4816,N_3687,N_4114);
nor U4817 (N_4817,N_3300,N_3924);
and U4818 (N_4818,N_4258,N_3665);
nor U4819 (N_4819,N_3482,N_4171);
xnor U4820 (N_4820,N_3828,N_3534);
nand U4821 (N_4821,N_3357,N_4352);
nor U4822 (N_4822,N_3556,N_3901);
xor U4823 (N_4823,N_3816,N_4323);
nand U4824 (N_4824,N_4119,N_4344);
nor U4825 (N_4825,N_4425,N_3452);
or U4826 (N_4826,N_4403,N_3138);
and U4827 (N_4827,N_4130,N_3533);
xnor U4828 (N_4828,N_3063,N_4253);
nor U4829 (N_4829,N_3549,N_3329);
and U4830 (N_4830,N_3989,N_3660);
nor U4831 (N_4831,N_4111,N_3865);
nand U4832 (N_4832,N_3059,N_3899);
nand U4833 (N_4833,N_3280,N_4252);
or U4834 (N_4834,N_3442,N_3095);
or U4835 (N_4835,N_3344,N_3223);
nand U4836 (N_4836,N_3811,N_3009);
or U4837 (N_4837,N_4255,N_4166);
nand U4838 (N_4838,N_3289,N_4311);
or U4839 (N_4839,N_3248,N_4183);
xor U4840 (N_4840,N_3873,N_3087);
nand U4841 (N_4841,N_3702,N_3477);
nand U4842 (N_4842,N_3317,N_3200);
nand U4843 (N_4843,N_3679,N_3337);
nand U4844 (N_4844,N_4132,N_3056);
nand U4845 (N_4845,N_3542,N_4484);
xor U4846 (N_4846,N_3510,N_3363);
and U4847 (N_4847,N_3000,N_4301);
and U4848 (N_4848,N_4295,N_3694);
or U4849 (N_4849,N_3369,N_3159);
and U4850 (N_4850,N_4281,N_3265);
nand U4851 (N_4851,N_3053,N_4392);
and U4852 (N_4852,N_3391,N_3868);
and U4853 (N_4853,N_3650,N_3202);
xor U4854 (N_4854,N_4070,N_4490);
and U4855 (N_4855,N_4146,N_3382);
or U4856 (N_4856,N_3065,N_3381);
and U4857 (N_4857,N_3069,N_4137);
nor U4858 (N_4858,N_4168,N_3526);
or U4859 (N_4859,N_3162,N_3195);
nor U4860 (N_4860,N_3509,N_3796);
nand U4861 (N_4861,N_3663,N_4179);
or U4862 (N_4862,N_4031,N_4256);
or U4863 (N_4863,N_3050,N_3604);
nor U4864 (N_4864,N_4293,N_4430);
and U4865 (N_4865,N_4317,N_3137);
nand U4866 (N_4866,N_4334,N_3889);
nor U4867 (N_4867,N_3955,N_3923);
or U4868 (N_4868,N_3259,N_4116);
nand U4869 (N_4869,N_3350,N_3314);
xnor U4870 (N_4870,N_4201,N_3692);
xor U4871 (N_4871,N_4473,N_3385);
and U4872 (N_4872,N_3268,N_3221);
xnor U4873 (N_4873,N_4271,N_3284);
nand U4874 (N_4874,N_4406,N_4180);
or U4875 (N_4875,N_3686,N_3158);
nand U4876 (N_4876,N_3698,N_3936);
and U4877 (N_4877,N_4228,N_3787);
and U4878 (N_4878,N_3012,N_3749);
xnor U4879 (N_4879,N_3455,N_4192);
xor U4880 (N_4880,N_3449,N_3199);
xor U4881 (N_4881,N_4475,N_4465);
xnor U4882 (N_4882,N_3192,N_3163);
nor U4883 (N_4883,N_4399,N_3566);
xor U4884 (N_4884,N_4342,N_3481);
xor U4885 (N_4885,N_3913,N_3301);
nor U4886 (N_4886,N_3746,N_4254);
nor U4887 (N_4887,N_3638,N_3515);
nor U4888 (N_4888,N_4350,N_4439);
nand U4889 (N_4889,N_3397,N_3883);
nand U4890 (N_4890,N_3522,N_4097);
xor U4891 (N_4891,N_3144,N_3772);
xnor U4892 (N_4892,N_4162,N_4185);
and U4893 (N_4893,N_3763,N_3076);
nand U4894 (N_4894,N_3759,N_4423);
or U4895 (N_4895,N_3557,N_3750);
or U4896 (N_4896,N_4223,N_3312);
xor U4897 (N_4897,N_3125,N_4016);
or U4898 (N_4898,N_3061,N_4195);
or U4899 (N_4899,N_3766,N_4327);
nand U4900 (N_4900,N_3880,N_4154);
xor U4901 (N_4901,N_3514,N_3214);
nand U4902 (N_4902,N_3257,N_3185);
xnor U4903 (N_4903,N_3833,N_3778);
nor U4904 (N_4904,N_3434,N_3952);
or U4905 (N_4905,N_4093,N_3547);
nor U4906 (N_4906,N_3343,N_3103);
nor U4907 (N_4907,N_4136,N_4194);
nand U4908 (N_4908,N_3109,N_3964);
xnor U4909 (N_4909,N_3048,N_3042);
or U4910 (N_4910,N_3977,N_3404);
or U4911 (N_4911,N_3082,N_3747);
xnor U4912 (N_4912,N_3255,N_3457);
nand U4913 (N_4913,N_3697,N_3710);
or U4914 (N_4914,N_3099,N_3324);
xor U4915 (N_4915,N_3368,N_4135);
xor U4916 (N_4916,N_3721,N_3589);
xor U4917 (N_4917,N_4089,N_3893);
or U4918 (N_4918,N_4056,N_3376);
and U4919 (N_4919,N_3078,N_4290);
or U4920 (N_4920,N_3122,N_4231);
nand U4921 (N_4921,N_3292,N_3794);
or U4922 (N_4922,N_4155,N_3628);
xor U4923 (N_4923,N_3015,N_3607);
or U4924 (N_4924,N_4240,N_3998);
xor U4925 (N_4925,N_4181,N_3523);
or U4926 (N_4926,N_3770,N_3166);
and U4927 (N_4927,N_4186,N_3890);
nor U4928 (N_4928,N_4260,N_3128);
nor U4929 (N_4929,N_3110,N_3541);
nand U4930 (N_4930,N_4077,N_3585);
nor U4931 (N_4931,N_3462,N_3187);
nand U4932 (N_4932,N_3577,N_3001);
and U4933 (N_4933,N_3196,N_4383);
xnor U4934 (N_4934,N_3405,N_3352);
nand U4935 (N_4935,N_3249,N_3695);
or U4936 (N_4936,N_3722,N_4131);
or U4937 (N_4937,N_3905,N_3862);
and U4938 (N_4938,N_3693,N_4328);
nand U4939 (N_4939,N_3444,N_3360);
or U4940 (N_4940,N_3290,N_3723);
or U4941 (N_4941,N_3491,N_4453);
nand U4942 (N_4942,N_4489,N_3555);
nand U4943 (N_4943,N_4416,N_4075);
nor U4944 (N_4944,N_3567,N_4035);
and U4945 (N_4945,N_4360,N_3459);
and U4946 (N_4946,N_3073,N_3519);
or U4947 (N_4947,N_3480,N_4338);
nor U4948 (N_4948,N_4085,N_3453);
or U4949 (N_4949,N_4105,N_3062);
xor U4950 (N_4950,N_3240,N_4375);
nand U4951 (N_4951,N_3940,N_3377);
nand U4952 (N_4952,N_3014,N_3974);
nor U4953 (N_4953,N_4241,N_4084);
nand U4954 (N_4954,N_3493,N_3801);
nor U4955 (N_4955,N_3269,N_3717);
and U4956 (N_4956,N_3950,N_3321);
nand U4957 (N_4957,N_4045,N_4496);
xor U4958 (N_4958,N_4393,N_4395);
or U4959 (N_4959,N_4006,N_3630);
or U4960 (N_4960,N_3277,N_3624);
xnor U4961 (N_4961,N_4034,N_3263);
or U4962 (N_4962,N_3283,N_4373);
xor U4963 (N_4963,N_3029,N_3815);
nor U4964 (N_4964,N_3260,N_4408);
nor U4965 (N_4965,N_3817,N_3193);
and U4966 (N_4966,N_3716,N_4282);
nor U4967 (N_4967,N_3207,N_3599);
or U4968 (N_4968,N_4133,N_4435);
and U4969 (N_4969,N_3619,N_3018);
nor U4970 (N_4970,N_4014,N_3320);
nor U4971 (N_4971,N_4308,N_4203);
or U4972 (N_4972,N_3229,N_4415);
or U4973 (N_4973,N_4040,N_4112);
or U4974 (N_4974,N_3070,N_4172);
nand U4975 (N_4975,N_4072,N_3521);
nor U4976 (N_4976,N_3010,N_3680);
nand U4977 (N_4977,N_4335,N_3780);
nand U4978 (N_4978,N_3035,N_4359);
nor U4979 (N_4979,N_3839,N_3219);
or U4980 (N_4980,N_3410,N_3458);
and U4981 (N_4981,N_4445,N_3446);
nor U4982 (N_4982,N_3610,N_4272);
nand U4983 (N_4983,N_4245,N_4189);
and U4984 (N_4984,N_4316,N_3851);
and U4985 (N_4985,N_3039,N_3961);
nand U4986 (N_4986,N_4134,N_3774);
or U4987 (N_4987,N_3544,N_4353);
nand U4988 (N_4988,N_3238,N_3859);
and U4989 (N_4989,N_3233,N_3250);
or U4990 (N_4990,N_3315,N_3701);
and U4991 (N_4991,N_3703,N_4023);
xor U4992 (N_4992,N_3928,N_4333);
nor U4993 (N_4993,N_4369,N_4142);
and U4994 (N_4994,N_4248,N_4004);
or U4995 (N_4995,N_3535,N_3838);
nor U4996 (N_4996,N_3258,N_3347);
xnor U4997 (N_4997,N_4424,N_3605);
nor U4998 (N_4998,N_4242,N_4042);
xor U4999 (N_4999,N_3294,N_3634);
or U5000 (N_5000,N_3313,N_3642);
nor U5001 (N_5001,N_3848,N_3842);
and U5002 (N_5002,N_3311,N_3956);
and U5003 (N_5003,N_4092,N_3068);
and U5004 (N_5004,N_4270,N_3083);
and U5005 (N_5005,N_3539,N_3016);
nor U5006 (N_5006,N_3483,N_3282);
or U5007 (N_5007,N_3981,N_3941);
nand U5008 (N_5008,N_4329,N_4145);
and U5009 (N_5009,N_3181,N_3188);
nor U5010 (N_5010,N_4307,N_4470);
xor U5011 (N_5011,N_4309,N_3896);
nor U5012 (N_5012,N_3764,N_3516);
nor U5013 (N_5013,N_4029,N_4417);
or U5014 (N_5014,N_3654,N_3148);
nor U5015 (N_5015,N_3133,N_3662);
nor U5016 (N_5016,N_3420,N_3371);
nor U5017 (N_5017,N_3670,N_3151);
xor U5018 (N_5018,N_3843,N_4261);
nand U5019 (N_5019,N_3653,N_3066);
nor U5020 (N_5020,N_4364,N_3945);
and U5021 (N_5021,N_3922,N_3323);
nor U5022 (N_5022,N_4280,N_3501);
nor U5023 (N_5023,N_3921,N_4108);
nor U5024 (N_5024,N_3609,N_3799);
or U5025 (N_5025,N_3812,N_4493);
or U5026 (N_5026,N_4012,N_4037);
nor U5027 (N_5027,N_3688,N_3506);
xor U5028 (N_5028,N_3571,N_3184);
or U5029 (N_5029,N_3094,N_3276);
nor U5030 (N_5030,N_3241,N_4207);
nand U5031 (N_5031,N_3330,N_3960);
xor U5032 (N_5032,N_3287,N_3091);
nor U5033 (N_5033,N_3390,N_3813);
nor U5034 (N_5034,N_4431,N_3972);
and U5035 (N_5035,N_3479,N_3906);
nor U5036 (N_5036,N_3303,N_4288);
nand U5037 (N_5037,N_4302,N_4220);
or U5038 (N_5038,N_3601,N_4332);
nand U5039 (N_5039,N_3574,N_4209);
xor U5040 (N_5040,N_3327,N_4222);
or U5041 (N_5041,N_3191,N_4129);
or U5042 (N_5042,N_3648,N_4161);
and U5043 (N_5043,N_3041,N_3278);
and U5044 (N_5044,N_4106,N_3573);
nor U5045 (N_5045,N_4420,N_4083);
xnor U5046 (N_5046,N_3210,N_3691);
xor U5047 (N_5047,N_3375,N_3165);
nand U5048 (N_5048,N_4343,N_3561);
nand U5049 (N_5049,N_3529,N_3003);
nand U5050 (N_5050,N_4152,N_3651);
nand U5051 (N_5051,N_3944,N_4474);
and U5052 (N_5052,N_4233,N_4019);
nor U5053 (N_5053,N_3807,N_3023);
nand U5054 (N_5054,N_4409,N_3342);
or U5055 (N_5055,N_3475,N_3550);
and U5056 (N_5056,N_4068,N_3712);
or U5057 (N_5057,N_3156,N_4059);
nand U5058 (N_5058,N_4079,N_4262);
and U5059 (N_5059,N_3614,N_3508);
xnor U5060 (N_5060,N_4049,N_4279);
nor U5061 (N_5061,N_4467,N_4027);
and U5062 (N_5062,N_3990,N_4266);
or U5063 (N_5063,N_3465,N_3396);
nand U5064 (N_5064,N_4410,N_3681);
or U5065 (N_5065,N_4357,N_3175);
nand U5066 (N_5066,N_3141,N_3307);
xor U5067 (N_5067,N_4257,N_3684);
xnor U5068 (N_5068,N_3592,N_3835);
nor U5069 (N_5069,N_3275,N_3597);
nor U5070 (N_5070,N_3611,N_4291);
or U5071 (N_5071,N_3038,N_3036);
nand U5072 (N_5072,N_4147,N_4126);
or U5073 (N_5073,N_3432,N_4101);
nor U5074 (N_5074,N_3847,N_3024);
and U5075 (N_5075,N_3525,N_3077);
xnor U5076 (N_5076,N_3777,N_3267);
xnor U5077 (N_5077,N_3554,N_3169);
nor U5078 (N_5078,N_4065,N_4234);
xnor U5079 (N_5079,N_3333,N_4339);
or U5080 (N_5080,N_3413,N_3055);
or U5081 (N_5081,N_3872,N_3019);
nor U5082 (N_5082,N_3666,N_3129);
or U5083 (N_5083,N_4200,N_4486);
and U5084 (N_5084,N_3545,N_3171);
xnor U5085 (N_5085,N_4109,N_3674);
and U5086 (N_5086,N_4197,N_3858);
xnor U5087 (N_5087,N_3878,N_3388);
and U5088 (N_5088,N_3781,N_3714);
xor U5089 (N_5089,N_3668,N_3841);
nand U5090 (N_5090,N_4394,N_3551);
nor U5091 (N_5091,N_3579,N_4123);
nor U5092 (N_5092,N_3005,N_3119);
xor U5093 (N_5093,N_4239,N_3335);
xnor U5094 (N_5094,N_4363,N_3768);
nand U5095 (N_5095,N_3866,N_3007);
or U5096 (N_5096,N_3231,N_3834);
nand U5097 (N_5097,N_3988,N_4444);
or U5098 (N_5098,N_3362,N_3080);
or U5099 (N_5099,N_3243,N_3017);
or U5100 (N_5100,N_4379,N_4286);
nor U5101 (N_5101,N_3985,N_3629);
nor U5102 (N_5102,N_3341,N_3429);
xor U5103 (N_5103,N_4438,N_4285);
or U5104 (N_5104,N_4366,N_4250);
nand U5105 (N_5105,N_3773,N_3882);
nor U5106 (N_5106,N_3951,N_3096);
nor U5107 (N_5107,N_3178,N_4259);
nand U5108 (N_5108,N_4361,N_4384);
xor U5109 (N_5109,N_4177,N_4355);
nor U5110 (N_5110,N_4125,N_4001);
or U5111 (N_5111,N_4115,N_4466);
xnor U5112 (N_5112,N_3946,N_3211);
nor U5113 (N_5113,N_4024,N_3884);
and U5114 (N_5114,N_4095,N_3216);
and U5115 (N_5115,N_4469,N_4224);
nand U5116 (N_5116,N_4213,N_4198);
xor U5117 (N_5117,N_3365,N_3052);
and U5118 (N_5118,N_3454,N_3532);
or U5119 (N_5119,N_4174,N_4098);
nor U5120 (N_5120,N_4216,N_3215);
xnor U5121 (N_5121,N_4401,N_4429);
xnor U5122 (N_5122,N_3993,N_3403);
xor U5123 (N_5123,N_3399,N_3658);
xor U5124 (N_5124,N_3468,N_4276);
or U5125 (N_5125,N_3902,N_3696);
or U5126 (N_5126,N_4073,N_3578);
and U5127 (N_5127,N_3160,N_3791);
xnor U5128 (N_5128,N_4265,N_3417);
nand U5129 (N_5129,N_3020,N_4076);
nand U5130 (N_5130,N_4441,N_3625);
xnor U5131 (N_5131,N_3810,N_4278);
nor U5132 (N_5132,N_3445,N_3885);
xor U5133 (N_5133,N_3060,N_4468);
nand U5134 (N_5134,N_4452,N_4380);
or U5135 (N_5135,N_3433,N_3253);
and U5136 (N_5136,N_4495,N_3118);
or U5137 (N_5137,N_4263,N_4071);
nor U5138 (N_5138,N_3524,N_3046);
and U5139 (N_5139,N_3673,N_3517);
xor U5140 (N_5140,N_3871,N_4463);
and U5141 (N_5141,N_3819,N_4143);
xor U5142 (N_5142,N_4268,N_3051);
or U5143 (N_5143,N_4087,N_3247);
or U5144 (N_5144,N_3440,N_3411);
and U5145 (N_5145,N_4021,N_3996);
nand U5146 (N_5146,N_3622,N_4378);
xnor U5147 (N_5147,N_4322,N_3291);
xnor U5148 (N_5148,N_3991,N_4020);
xor U5149 (N_5149,N_4330,N_4051);
and U5150 (N_5150,N_4303,N_3456);
nand U5151 (N_5151,N_3400,N_4289);
and U5152 (N_5152,N_4483,N_4211);
xor U5153 (N_5153,N_4028,N_3101);
nor U5154 (N_5154,N_3361,N_4321);
xnor U5155 (N_5155,N_4052,N_3494);
and U5156 (N_5156,N_4053,N_3503);
xor U5157 (N_5157,N_3531,N_3428);
xor U5158 (N_5158,N_3877,N_3336);
nor U5159 (N_5159,N_3837,N_4044);
nor U5160 (N_5160,N_3830,N_3172);
nor U5161 (N_5161,N_3424,N_3325);
nand U5162 (N_5162,N_4382,N_3725);
nor U5163 (N_5163,N_3771,N_3310);
or U5164 (N_5164,N_3669,N_4433);
nor U5165 (N_5165,N_3537,N_4331);
xnor U5166 (N_5166,N_4202,N_3802);
and U5167 (N_5167,N_3500,N_4491);
nand U5168 (N_5168,N_3354,N_3623);
xnor U5169 (N_5169,N_3685,N_4304);
nand U5170 (N_5170,N_4492,N_3814);
nand U5171 (N_5171,N_3072,N_3150);
or U5172 (N_5172,N_3826,N_3490);
or U5173 (N_5173,N_3593,N_3299);
xnor U5174 (N_5174,N_3308,N_3157);
or U5175 (N_5175,N_3640,N_4437);
and U5176 (N_5176,N_3613,N_3886);
nand U5177 (N_5177,N_4127,N_4472);
nand U5178 (N_5178,N_3881,N_3655);
xnor U5179 (N_5179,N_3728,N_3348);
or U5180 (N_5180,N_3603,N_3984);
or U5181 (N_5181,N_4193,N_3933);
nand U5182 (N_5182,N_3606,N_3025);
nand U5183 (N_5183,N_4249,N_3139);
xnor U5184 (N_5184,N_3114,N_3463);
xor U5185 (N_5185,N_3731,N_4229);
and U5186 (N_5186,N_4017,N_3064);
nand U5187 (N_5187,N_3735,N_4038);
and U5188 (N_5188,N_4199,N_4086);
nand U5189 (N_5189,N_4300,N_4325);
or U5190 (N_5190,N_3659,N_3174);
nor U5191 (N_5191,N_4000,N_4170);
and U5192 (N_5192,N_4348,N_3430);
xor U5193 (N_5193,N_3829,N_3447);
and U5194 (N_5194,N_4221,N_3620);
xnor U5195 (N_5195,N_3618,N_4050);
nand U5196 (N_5196,N_3031,N_3621);
or U5197 (N_5197,N_4074,N_3124);
nor U5198 (N_5198,N_3546,N_3903);
nor U5199 (N_5199,N_3757,N_3832);
and U5200 (N_5200,N_3564,N_3647);
nand U5201 (N_5201,N_4449,N_4026);
nand U5202 (N_5202,N_4005,N_4487);
or U5203 (N_5203,N_3560,N_4451);
nor U5204 (N_5204,N_3976,N_3598);
nor U5205 (N_5205,N_3997,N_3395);
nand U5206 (N_5206,N_4454,N_3326);
and U5207 (N_5207,N_3707,N_3134);
nor U5208 (N_5208,N_4080,N_4046);
or U5209 (N_5209,N_3854,N_4443);
xnor U5210 (N_5210,N_4102,N_4010);
nand U5211 (N_5211,N_3719,N_3013);
nand U5212 (N_5212,N_3978,N_4418);
and U5213 (N_5213,N_4214,N_3789);
or U5214 (N_5214,N_3784,N_3825);
and U5215 (N_5215,N_3758,N_3975);
or U5216 (N_5216,N_3074,N_3938);
and U5217 (N_5217,N_3176,N_3093);
nor U5218 (N_5218,N_3492,N_3930);
nor U5219 (N_5219,N_3720,N_3098);
nand U5220 (N_5220,N_4206,N_3994);
xor U5221 (N_5221,N_3285,N_3718);
xor U5222 (N_5222,N_4151,N_3907);
or U5223 (N_5223,N_3876,N_3616);
nor U5224 (N_5224,N_3729,N_3497);
nand U5225 (N_5225,N_3580,N_3512);
xnor U5226 (N_5226,N_4422,N_3645);
and U5227 (N_5227,N_3349,N_4025);
nand U5228 (N_5228,N_3351,N_3293);
and U5229 (N_5229,N_4011,N_3850);
nor U5230 (N_5230,N_4232,N_4349);
xor U5231 (N_5231,N_3107,N_3218);
and U5232 (N_5232,N_4188,N_4128);
nor U5233 (N_5233,N_3288,N_3823);
or U5234 (N_5234,N_3920,N_3916);
or U5235 (N_5235,N_3081,N_4432);
and U5236 (N_5236,N_4419,N_3054);
and U5237 (N_5237,N_4464,N_3748);
or U5238 (N_5238,N_3743,N_3306);
nor U5239 (N_5239,N_3558,N_3934);
nor U5240 (N_5240,N_4208,N_3676);
or U5241 (N_5241,N_3675,N_3246);
and U5242 (N_5242,N_4096,N_4298);
and U5243 (N_5243,N_3478,N_3356);
and U5244 (N_5244,N_3954,N_4120);
and U5245 (N_5245,N_3904,N_4477);
nor U5246 (N_5246,N_4400,N_3831);
nand U5247 (N_5247,N_3470,N_3135);
or U5248 (N_5248,N_3891,N_3474);
nand U5249 (N_5249,N_3809,N_3612);
nor U5250 (N_5250,N_4167,N_4321);
xor U5251 (N_5251,N_3203,N_3181);
nand U5252 (N_5252,N_3023,N_4381);
and U5253 (N_5253,N_3257,N_3651);
nand U5254 (N_5254,N_3234,N_3492);
nor U5255 (N_5255,N_4125,N_3304);
xor U5256 (N_5256,N_4416,N_4180);
nand U5257 (N_5257,N_3345,N_4480);
and U5258 (N_5258,N_3102,N_3475);
xnor U5259 (N_5259,N_4315,N_3268);
and U5260 (N_5260,N_4335,N_3487);
or U5261 (N_5261,N_4203,N_4277);
nand U5262 (N_5262,N_3842,N_4174);
nor U5263 (N_5263,N_3769,N_4233);
or U5264 (N_5264,N_3297,N_3319);
xnor U5265 (N_5265,N_3634,N_4169);
xor U5266 (N_5266,N_3125,N_3089);
or U5267 (N_5267,N_4422,N_3591);
and U5268 (N_5268,N_3188,N_3819);
xnor U5269 (N_5269,N_3729,N_3895);
nor U5270 (N_5270,N_3208,N_4173);
nor U5271 (N_5271,N_3407,N_4097);
nor U5272 (N_5272,N_3191,N_3929);
xnor U5273 (N_5273,N_3345,N_3598);
nand U5274 (N_5274,N_3778,N_3957);
nand U5275 (N_5275,N_3220,N_3651);
or U5276 (N_5276,N_3878,N_3351);
nand U5277 (N_5277,N_3648,N_3647);
or U5278 (N_5278,N_3732,N_3036);
or U5279 (N_5279,N_4306,N_3374);
nand U5280 (N_5280,N_3279,N_4036);
or U5281 (N_5281,N_4405,N_3191);
xor U5282 (N_5282,N_3425,N_3111);
xor U5283 (N_5283,N_4028,N_4378);
nand U5284 (N_5284,N_3490,N_4265);
nor U5285 (N_5285,N_3831,N_4304);
nor U5286 (N_5286,N_4386,N_3957);
xnor U5287 (N_5287,N_3528,N_3017);
nor U5288 (N_5288,N_3538,N_3769);
xor U5289 (N_5289,N_3475,N_3364);
or U5290 (N_5290,N_3692,N_4262);
nand U5291 (N_5291,N_3284,N_3035);
nand U5292 (N_5292,N_3544,N_3026);
or U5293 (N_5293,N_4404,N_3946);
xor U5294 (N_5294,N_4110,N_4078);
xor U5295 (N_5295,N_3315,N_4386);
nand U5296 (N_5296,N_4025,N_3065);
and U5297 (N_5297,N_3653,N_3080);
and U5298 (N_5298,N_3564,N_4313);
nor U5299 (N_5299,N_3695,N_3769);
or U5300 (N_5300,N_4361,N_3100);
nand U5301 (N_5301,N_3992,N_4168);
nand U5302 (N_5302,N_4033,N_4074);
nor U5303 (N_5303,N_3141,N_4078);
or U5304 (N_5304,N_4423,N_3802);
and U5305 (N_5305,N_3896,N_3257);
and U5306 (N_5306,N_3347,N_4467);
or U5307 (N_5307,N_3693,N_4108);
and U5308 (N_5308,N_3483,N_3466);
nand U5309 (N_5309,N_3426,N_3031);
nand U5310 (N_5310,N_3833,N_3011);
nor U5311 (N_5311,N_4091,N_3458);
or U5312 (N_5312,N_3819,N_3554);
nand U5313 (N_5313,N_3801,N_3221);
or U5314 (N_5314,N_4114,N_3876);
xor U5315 (N_5315,N_3256,N_3517);
nor U5316 (N_5316,N_4475,N_4490);
or U5317 (N_5317,N_4044,N_3198);
xor U5318 (N_5318,N_3765,N_3932);
nor U5319 (N_5319,N_4491,N_3821);
nand U5320 (N_5320,N_3224,N_3147);
nor U5321 (N_5321,N_4088,N_3945);
xor U5322 (N_5322,N_3957,N_4468);
xor U5323 (N_5323,N_4112,N_4271);
xor U5324 (N_5324,N_4365,N_3556);
xnor U5325 (N_5325,N_3026,N_3983);
xor U5326 (N_5326,N_3759,N_3583);
nand U5327 (N_5327,N_3649,N_3001);
or U5328 (N_5328,N_3632,N_4266);
nor U5329 (N_5329,N_3012,N_3092);
or U5330 (N_5330,N_4364,N_3328);
xnor U5331 (N_5331,N_4232,N_4477);
xor U5332 (N_5332,N_3875,N_3483);
xor U5333 (N_5333,N_4381,N_3188);
nor U5334 (N_5334,N_3206,N_3314);
or U5335 (N_5335,N_3576,N_3306);
nor U5336 (N_5336,N_4383,N_3676);
nor U5337 (N_5337,N_3290,N_3966);
nor U5338 (N_5338,N_3145,N_3435);
nand U5339 (N_5339,N_3279,N_4180);
and U5340 (N_5340,N_4447,N_3649);
nand U5341 (N_5341,N_3468,N_3204);
nor U5342 (N_5342,N_4206,N_3440);
and U5343 (N_5343,N_3462,N_3080);
nor U5344 (N_5344,N_3217,N_4114);
nor U5345 (N_5345,N_3733,N_3856);
or U5346 (N_5346,N_3676,N_3058);
xor U5347 (N_5347,N_3156,N_3114);
nand U5348 (N_5348,N_3495,N_4393);
and U5349 (N_5349,N_3369,N_4181);
nor U5350 (N_5350,N_4349,N_4409);
nand U5351 (N_5351,N_4237,N_3752);
and U5352 (N_5352,N_3541,N_3821);
nand U5353 (N_5353,N_4303,N_3926);
nor U5354 (N_5354,N_3956,N_4304);
nor U5355 (N_5355,N_3964,N_3316);
nor U5356 (N_5356,N_3770,N_3022);
xnor U5357 (N_5357,N_3603,N_3977);
xnor U5358 (N_5358,N_4167,N_3365);
or U5359 (N_5359,N_3192,N_3853);
and U5360 (N_5360,N_3418,N_3261);
xor U5361 (N_5361,N_4167,N_3070);
nand U5362 (N_5362,N_3651,N_3729);
xnor U5363 (N_5363,N_3709,N_3529);
nor U5364 (N_5364,N_3189,N_3166);
or U5365 (N_5365,N_3001,N_3436);
or U5366 (N_5366,N_3358,N_4168);
xor U5367 (N_5367,N_3574,N_3152);
nand U5368 (N_5368,N_3144,N_3834);
xor U5369 (N_5369,N_4310,N_4130);
nor U5370 (N_5370,N_3803,N_3163);
and U5371 (N_5371,N_4473,N_3490);
nor U5372 (N_5372,N_3082,N_3198);
nand U5373 (N_5373,N_4136,N_3946);
nor U5374 (N_5374,N_4410,N_3572);
nand U5375 (N_5375,N_4357,N_4193);
or U5376 (N_5376,N_3916,N_4162);
nand U5377 (N_5377,N_3251,N_4432);
or U5378 (N_5378,N_4194,N_3840);
or U5379 (N_5379,N_3976,N_4153);
and U5380 (N_5380,N_3200,N_4341);
xnor U5381 (N_5381,N_4145,N_3917);
nand U5382 (N_5382,N_4027,N_3660);
xnor U5383 (N_5383,N_3737,N_4282);
nand U5384 (N_5384,N_4107,N_3862);
nor U5385 (N_5385,N_3140,N_4372);
xor U5386 (N_5386,N_3847,N_4278);
nand U5387 (N_5387,N_4306,N_3952);
or U5388 (N_5388,N_4021,N_3162);
nand U5389 (N_5389,N_3863,N_4465);
xor U5390 (N_5390,N_3358,N_3644);
and U5391 (N_5391,N_3015,N_4187);
nand U5392 (N_5392,N_3322,N_4387);
nor U5393 (N_5393,N_3859,N_4416);
nor U5394 (N_5394,N_4185,N_3268);
nor U5395 (N_5395,N_3862,N_3998);
nand U5396 (N_5396,N_4331,N_4058);
xnor U5397 (N_5397,N_3049,N_4111);
nor U5398 (N_5398,N_3185,N_4436);
nand U5399 (N_5399,N_4289,N_3714);
or U5400 (N_5400,N_3537,N_3454);
nor U5401 (N_5401,N_3201,N_3487);
and U5402 (N_5402,N_3442,N_4216);
xor U5403 (N_5403,N_3958,N_4360);
or U5404 (N_5404,N_3263,N_4262);
nand U5405 (N_5405,N_3764,N_3234);
or U5406 (N_5406,N_3006,N_3050);
nand U5407 (N_5407,N_3135,N_3172);
xor U5408 (N_5408,N_3171,N_3633);
or U5409 (N_5409,N_3662,N_3887);
nor U5410 (N_5410,N_4004,N_3960);
xor U5411 (N_5411,N_3832,N_4189);
or U5412 (N_5412,N_4109,N_4392);
nand U5413 (N_5413,N_3730,N_4254);
or U5414 (N_5414,N_3344,N_3872);
or U5415 (N_5415,N_3786,N_3493);
xnor U5416 (N_5416,N_3398,N_3857);
nand U5417 (N_5417,N_3582,N_3971);
and U5418 (N_5418,N_4437,N_3469);
xnor U5419 (N_5419,N_3993,N_4009);
xor U5420 (N_5420,N_4455,N_3403);
or U5421 (N_5421,N_3689,N_3114);
or U5422 (N_5422,N_3945,N_4203);
and U5423 (N_5423,N_3131,N_4175);
and U5424 (N_5424,N_4062,N_3371);
nand U5425 (N_5425,N_3079,N_3866);
or U5426 (N_5426,N_3433,N_4130);
or U5427 (N_5427,N_4463,N_3047);
nor U5428 (N_5428,N_4156,N_3700);
nand U5429 (N_5429,N_3495,N_3546);
nor U5430 (N_5430,N_4470,N_3936);
xnor U5431 (N_5431,N_3145,N_3368);
or U5432 (N_5432,N_3432,N_3494);
nor U5433 (N_5433,N_3633,N_3610);
or U5434 (N_5434,N_3963,N_3926);
xnor U5435 (N_5435,N_4437,N_4054);
nor U5436 (N_5436,N_3353,N_3625);
or U5437 (N_5437,N_3509,N_3722);
nand U5438 (N_5438,N_4460,N_4112);
or U5439 (N_5439,N_4470,N_4297);
nand U5440 (N_5440,N_4075,N_4338);
or U5441 (N_5441,N_4173,N_3964);
nor U5442 (N_5442,N_3598,N_3998);
nor U5443 (N_5443,N_3603,N_4342);
or U5444 (N_5444,N_4290,N_3043);
and U5445 (N_5445,N_3890,N_3937);
xor U5446 (N_5446,N_3083,N_4175);
and U5447 (N_5447,N_3564,N_4085);
nor U5448 (N_5448,N_4460,N_3472);
and U5449 (N_5449,N_4081,N_3220);
nand U5450 (N_5450,N_4300,N_4454);
xor U5451 (N_5451,N_3192,N_3311);
xor U5452 (N_5452,N_4135,N_4355);
nand U5453 (N_5453,N_3500,N_3295);
or U5454 (N_5454,N_3120,N_4121);
nor U5455 (N_5455,N_3870,N_3995);
nand U5456 (N_5456,N_3815,N_3059);
or U5457 (N_5457,N_4435,N_3462);
and U5458 (N_5458,N_4238,N_4098);
xnor U5459 (N_5459,N_4262,N_3896);
and U5460 (N_5460,N_3446,N_3539);
and U5461 (N_5461,N_3502,N_3219);
or U5462 (N_5462,N_3157,N_3272);
or U5463 (N_5463,N_3232,N_4374);
nor U5464 (N_5464,N_4419,N_3712);
and U5465 (N_5465,N_3579,N_3205);
nand U5466 (N_5466,N_3205,N_3595);
and U5467 (N_5467,N_3194,N_3848);
or U5468 (N_5468,N_3867,N_3759);
nand U5469 (N_5469,N_4220,N_3385);
or U5470 (N_5470,N_3805,N_3813);
and U5471 (N_5471,N_4414,N_3086);
nand U5472 (N_5472,N_3994,N_3316);
nand U5473 (N_5473,N_4112,N_3477);
and U5474 (N_5474,N_3896,N_4406);
xor U5475 (N_5475,N_3845,N_4239);
or U5476 (N_5476,N_3161,N_3404);
or U5477 (N_5477,N_3174,N_4355);
nor U5478 (N_5478,N_3227,N_3696);
and U5479 (N_5479,N_4032,N_4118);
xor U5480 (N_5480,N_3082,N_3248);
and U5481 (N_5481,N_4404,N_3392);
nor U5482 (N_5482,N_3470,N_4360);
nor U5483 (N_5483,N_3579,N_3033);
nor U5484 (N_5484,N_4165,N_4123);
xnor U5485 (N_5485,N_3280,N_4130);
nand U5486 (N_5486,N_4364,N_3236);
or U5487 (N_5487,N_4073,N_3246);
or U5488 (N_5488,N_3043,N_3447);
nand U5489 (N_5489,N_3845,N_4249);
or U5490 (N_5490,N_4468,N_3748);
xor U5491 (N_5491,N_3524,N_3860);
and U5492 (N_5492,N_4058,N_4281);
or U5493 (N_5493,N_4385,N_3185);
and U5494 (N_5494,N_3512,N_3419);
xnor U5495 (N_5495,N_3115,N_3346);
nor U5496 (N_5496,N_4200,N_3034);
nand U5497 (N_5497,N_3568,N_3621);
and U5498 (N_5498,N_3652,N_4168);
and U5499 (N_5499,N_3906,N_3648);
nand U5500 (N_5500,N_4452,N_4279);
and U5501 (N_5501,N_3689,N_3752);
nand U5502 (N_5502,N_3479,N_4433);
nor U5503 (N_5503,N_4395,N_4018);
nor U5504 (N_5504,N_3414,N_4460);
and U5505 (N_5505,N_3297,N_3962);
nand U5506 (N_5506,N_3615,N_3549);
and U5507 (N_5507,N_4104,N_3273);
xnor U5508 (N_5508,N_4060,N_3122);
nor U5509 (N_5509,N_3267,N_3450);
and U5510 (N_5510,N_4200,N_4178);
xnor U5511 (N_5511,N_3231,N_3181);
or U5512 (N_5512,N_3953,N_4137);
nor U5513 (N_5513,N_3604,N_3765);
nand U5514 (N_5514,N_3734,N_3826);
and U5515 (N_5515,N_4134,N_3192);
nor U5516 (N_5516,N_3443,N_3128);
xnor U5517 (N_5517,N_3102,N_3266);
nor U5518 (N_5518,N_3749,N_3373);
or U5519 (N_5519,N_3429,N_3241);
and U5520 (N_5520,N_3186,N_4367);
nor U5521 (N_5521,N_4426,N_4058);
and U5522 (N_5522,N_4394,N_4482);
xor U5523 (N_5523,N_3744,N_3492);
or U5524 (N_5524,N_3936,N_3244);
xnor U5525 (N_5525,N_3695,N_3059);
or U5526 (N_5526,N_3733,N_4283);
or U5527 (N_5527,N_3677,N_3087);
nor U5528 (N_5528,N_4093,N_3493);
nor U5529 (N_5529,N_3401,N_4429);
and U5530 (N_5530,N_3696,N_4405);
nor U5531 (N_5531,N_4316,N_4082);
nand U5532 (N_5532,N_3216,N_3244);
xnor U5533 (N_5533,N_3168,N_4419);
xnor U5534 (N_5534,N_4451,N_4079);
xnor U5535 (N_5535,N_4279,N_4108);
or U5536 (N_5536,N_4182,N_3043);
nand U5537 (N_5537,N_3413,N_4233);
and U5538 (N_5538,N_3230,N_4030);
nor U5539 (N_5539,N_3422,N_3572);
nand U5540 (N_5540,N_4375,N_4419);
and U5541 (N_5541,N_3007,N_3944);
xnor U5542 (N_5542,N_4032,N_4165);
nand U5543 (N_5543,N_4158,N_3118);
or U5544 (N_5544,N_3431,N_3201);
nor U5545 (N_5545,N_3201,N_3669);
or U5546 (N_5546,N_4068,N_3002);
nand U5547 (N_5547,N_3090,N_4019);
xor U5548 (N_5548,N_3720,N_3630);
xnor U5549 (N_5549,N_3359,N_3382);
and U5550 (N_5550,N_3899,N_4090);
nand U5551 (N_5551,N_4226,N_3327);
or U5552 (N_5552,N_3710,N_3121);
or U5553 (N_5553,N_3235,N_4093);
or U5554 (N_5554,N_3032,N_3363);
nor U5555 (N_5555,N_3614,N_3018);
nor U5556 (N_5556,N_4221,N_4137);
and U5557 (N_5557,N_4001,N_4144);
xnor U5558 (N_5558,N_3548,N_3512);
nand U5559 (N_5559,N_3209,N_3359);
xor U5560 (N_5560,N_3468,N_3038);
nand U5561 (N_5561,N_4316,N_3402);
nand U5562 (N_5562,N_3225,N_3641);
and U5563 (N_5563,N_3955,N_4219);
xor U5564 (N_5564,N_4115,N_4395);
or U5565 (N_5565,N_4066,N_3047);
xor U5566 (N_5566,N_4394,N_3904);
and U5567 (N_5567,N_3967,N_3485);
nor U5568 (N_5568,N_3845,N_3644);
xor U5569 (N_5569,N_3440,N_4073);
nand U5570 (N_5570,N_3377,N_3037);
or U5571 (N_5571,N_4374,N_3625);
nor U5572 (N_5572,N_3184,N_3460);
or U5573 (N_5573,N_4431,N_3705);
and U5574 (N_5574,N_3078,N_3187);
xnor U5575 (N_5575,N_3387,N_3208);
and U5576 (N_5576,N_4172,N_4284);
xnor U5577 (N_5577,N_3689,N_3121);
xor U5578 (N_5578,N_3933,N_3877);
nand U5579 (N_5579,N_3102,N_3373);
or U5580 (N_5580,N_3399,N_4426);
or U5581 (N_5581,N_3344,N_3968);
nand U5582 (N_5582,N_3982,N_3124);
nor U5583 (N_5583,N_3032,N_3062);
nor U5584 (N_5584,N_3410,N_3277);
nor U5585 (N_5585,N_3769,N_3706);
or U5586 (N_5586,N_4256,N_3074);
nor U5587 (N_5587,N_3683,N_3333);
and U5588 (N_5588,N_3977,N_3469);
xor U5589 (N_5589,N_4241,N_3832);
or U5590 (N_5590,N_3397,N_3470);
or U5591 (N_5591,N_4018,N_3874);
xor U5592 (N_5592,N_4245,N_3290);
or U5593 (N_5593,N_3692,N_3684);
nand U5594 (N_5594,N_4138,N_3105);
and U5595 (N_5595,N_4413,N_3273);
xnor U5596 (N_5596,N_3744,N_3044);
or U5597 (N_5597,N_3418,N_4172);
xor U5598 (N_5598,N_3945,N_4321);
or U5599 (N_5599,N_3728,N_3876);
or U5600 (N_5600,N_3740,N_3511);
nor U5601 (N_5601,N_4331,N_4439);
nand U5602 (N_5602,N_3458,N_3990);
xnor U5603 (N_5603,N_4331,N_3174);
or U5604 (N_5604,N_3274,N_3701);
and U5605 (N_5605,N_4265,N_4341);
xor U5606 (N_5606,N_4499,N_3414);
and U5607 (N_5607,N_3162,N_4291);
nand U5608 (N_5608,N_3266,N_3508);
nand U5609 (N_5609,N_3873,N_3357);
nand U5610 (N_5610,N_3639,N_4496);
nand U5611 (N_5611,N_4439,N_4297);
nor U5612 (N_5612,N_4337,N_4320);
and U5613 (N_5613,N_4008,N_3976);
and U5614 (N_5614,N_3483,N_4258);
nand U5615 (N_5615,N_3306,N_3870);
or U5616 (N_5616,N_3208,N_3797);
xnor U5617 (N_5617,N_3681,N_4057);
nand U5618 (N_5618,N_4240,N_3096);
and U5619 (N_5619,N_3936,N_4463);
xnor U5620 (N_5620,N_3682,N_4479);
nor U5621 (N_5621,N_4192,N_3475);
nor U5622 (N_5622,N_3769,N_3447);
nand U5623 (N_5623,N_3727,N_3476);
nand U5624 (N_5624,N_3427,N_4244);
and U5625 (N_5625,N_3728,N_3614);
xnor U5626 (N_5626,N_4078,N_3905);
nor U5627 (N_5627,N_4020,N_3107);
and U5628 (N_5628,N_3334,N_3115);
nor U5629 (N_5629,N_3084,N_4023);
nor U5630 (N_5630,N_3353,N_4420);
or U5631 (N_5631,N_3401,N_4209);
and U5632 (N_5632,N_4079,N_4288);
or U5633 (N_5633,N_4088,N_3952);
nor U5634 (N_5634,N_3733,N_3947);
nor U5635 (N_5635,N_3415,N_3348);
xor U5636 (N_5636,N_4256,N_4130);
nand U5637 (N_5637,N_3158,N_3951);
nand U5638 (N_5638,N_3000,N_3116);
or U5639 (N_5639,N_3147,N_4427);
xnor U5640 (N_5640,N_3355,N_3516);
nand U5641 (N_5641,N_3595,N_4385);
nand U5642 (N_5642,N_3065,N_3417);
or U5643 (N_5643,N_3412,N_3141);
nand U5644 (N_5644,N_3523,N_4000);
and U5645 (N_5645,N_4380,N_4386);
or U5646 (N_5646,N_3713,N_3751);
nand U5647 (N_5647,N_3682,N_4106);
xnor U5648 (N_5648,N_3032,N_3796);
and U5649 (N_5649,N_3055,N_3501);
nor U5650 (N_5650,N_4151,N_3713);
xor U5651 (N_5651,N_3268,N_3266);
nor U5652 (N_5652,N_3365,N_3569);
xnor U5653 (N_5653,N_4180,N_4328);
and U5654 (N_5654,N_3538,N_3758);
or U5655 (N_5655,N_3781,N_3138);
nand U5656 (N_5656,N_3386,N_4362);
nand U5657 (N_5657,N_4371,N_3645);
nor U5658 (N_5658,N_4334,N_3822);
nand U5659 (N_5659,N_3911,N_4185);
xor U5660 (N_5660,N_4461,N_3063);
nor U5661 (N_5661,N_3574,N_3621);
nand U5662 (N_5662,N_4397,N_3889);
and U5663 (N_5663,N_3948,N_3660);
or U5664 (N_5664,N_3773,N_3025);
and U5665 (N_5665,N_4379,N_4367);
and U5666 (N_5666,N_3781,N_4111);
xnor U5667 (N_5667,N_4441,N_3474);
nand U5668 (N_5668,N_3295,N_3064);
nor U5669 (N_5669,N_4238,N_3612);
nand U5670 (N_5670,N_3049,N_4268);
or U5671 (N_5671,N_3285,N_4256);
nand U5672 (N_5672,N_4409,N_3690);
xnor U5673 (N_5673,N_3674,N_3173);
or U5674 (N_5674,N_3256,N_4191);
or U5675 (N_5675,N_4258,N_3595);
nand U5676 (N_5676,N_4100,N_3006);
nand U5677 (N_5677,N_4254,N_4111);
or U5678 (N_5678,N_4021,N_3163);
and U5679 (N_5679,N_3500,N_3808);
or U5680 (N_5680,N_4451,N_3513);
nor U5681 (N_5681,N_4223,N_4272);
xnor U5682 (N_5682,N_4235,N_3710);
xor U5683 (N_5683,N_3127,N_4251);
or U5684 (N_5684,N_4441,N_3821);
or U5685 (N_5685,N_4301,N_3556);
xor U5686 (N_5686,N_3371,N_4146);
nor U5687 (N_5687,N_4171,N_3635);
nor U5688 (N_5688,N_4332,N_4027);
or U5689 (N_5689,N_4398,N_3334);
nand U5690 (N_5690,N_3430,N_4121);
xnor U5691 (N_5691,N_3701,N_3876);
and U5692 (N_5692,N_4267,N_3196);
xor U5693 (N_5693,N_4234,N_4477);
nand U5694 (N_5694,N_4219,N_3431);
xnor U5695 (N_5695,N_4216,N_3829);
nand U5696 (N_5696,N_3620,N_3200);
xnor U5697 (N_5697,N_3779,N_3529);
or U5698 (N_5698,N_3584,N_4479);
nand U5699 (N_5699,N_4288,N_3957);
or U5700 (N_5700,N_3700,N_4499);
or U5701 (N_5701,N_4214,N_3319);
nand U5702 (N_5702,N_3142,N_3035);
nand U5703 (N_5703,N_3399,N_4104);
or U5704 (N_5704,N_3353,N_3658);
or U5705 (N_5705,N_3442,N_4009);
nor U5706 (N_5706,N_4489,N_3439);
xnor U5707 (N_5707,N_3189,N_3213);
or U5708 (N_5708,N_3065,N_3805);
and U5709 (N_5709,N_4256,N_3681);
or U5710 (N_5710,N_4144,N_4358);
xor U5711 (N_5711,N_4104,N_3052);
nand U5712 (N_5712,N_4203,N_3410);
nand U5713 (N_5713,N_3496,N_3962);
nor U5714 (N_5714,N_4251,N_3853);
nand U5715 (N_5715,N_4280,N_4462);
xnor U5716 (N_5716,N_4395,N_4218);
xor U5717 (N_5717,N_3913,N_4446);
or U5718 (N_5718,N_3045,N_4367);
and U5719 (N_5719,N_3713,N_3601);
and U5720 (N_5720,N_4286,N_4080);
nor U5721 (N_5721,N_3968,N_3432);
or U5722 (N_5722,N_3054,N_4193);
nor U5723 (N_5723,N_3195,N_3134);
xor U5724 (N_5724,N_3372,N_3270);
or U5725 (N_5725,N_3780,N_4192);
or U5726 (N_5726,N_3276,N_4328);
nor U5727 (N_5727,N_3996,N_4264);
or U5728 (N_5728,N_4335,N_3404);
or U5729 (N_5729,N_3093,N_3834);
nand U5730 (N_5730,N_3823,N_4132);
and U5731 (N_5731,N_3065,N_4347);
nor U5732 (N_5732,N_4087,N_3828);
xnor U5733 (N_5733,N_4156,N_4206);
xnor U5734 (N_5734,N_3666,N_4054);
and U5735 (N_5735,N_3544,N_4125);
xnor U5736 (N_5736,N_3337,N_4468);
xor U5737 (N_5737,N_3134,N_4283);
xor U5738 (N_5738,N_3342,N_3735);
nand U5739 (N_5739,N_3435,N_3673);
and U5740 (N_5740,N_3951,N_4024);
nand U5741 (N_5741,N_3017,N_4431);
nor U5742 (N_5742,N_3416,N_3088);
nand U5743 (N_5743,N_3874,N_3442);
and U5744 (N_5744,N_3056,N_3572);
and U5745 (N_5745,N_3020,N_4107);
and U5746 (N_5746,N_3677,N_3315);
or U5747 (N_5747,N_3357,N_3438);
and U5748 (N_5748,N_3266,N_3110);
or U5749 (N_5749,N_3354,N_3144);
or U5750 (N_5750,N_3356,N_3549);
nand U5751 (N_5751,N_3966,N_3360);
xor U5752 (N_5752,N_3584,N_3526);
and U5753 (N_5753,N_3320,N_4325);
nand U5754 (N_5754,N_3336,N_3193);
and U5755 (N_5755,N_3850,N_4089);
xnor U5756 (N_5756,N_3117,N_3024);
xnor U5757 (N_5757,N_3377,N_4375);
and U5758 (N_5758,N_3410,N_4008);
xor U5759 (N_5759,N_3409,N_3459);
xor U5760 (N_5760,N_3546,N_4480);
nand U5761 (N_5761,N_3817,N_4296);
nand U5762 (N_5762,N_3831,N_3066);
or U5763 (N_5763,N_4449,N_3351);
xnor U5764 (N_5764,N_3843,N_4076);
nand U5765 (N_5765,N_3106,N_4471);
nand U5766 (N_5766,N_3139,N_4114);
and U5767 (N_5767,N_3216,N_4104);
nor U5768 (N_5768,N_4195,N_4449);
or U5769 (N_5769,N_3615,N_3253);
or U5770 (N_5770,N_3319,N_4231);
or U5771 (N_5771,N_4333,N_4204);
xnor U5772 (N_5772,N_4065,N_4317);
xor U5773 (N_5773,N_3821,N_3815);
nand U5774 (N_5774,N_3849,N_3499);
nor U5775 (N_5775,N_3301,N_4337);
and U5776 (N_5776,N_3714,N_3856);
nand U5777 (N_5777,N_3409,N_3536);
or U5778 (N_5778,N_3617,N_3948);
or U5779 (N_5779,N_3252,N_3316);
nor U5780 (N_5780,N_3244,N_3967);
nand U5781 (N_5781,N_4378,N_3231);
nor U5782 (N_5782,N_3550,N_3349);
nor U5783 (N_5783,N_4225,N_3581);
nand U5784 (N_5784,N_4249,N_3972);
and U5785 (N_5785,N_3890,N_3208);
and U5786 (N_5786,N_3294,N_3671);
nor U5787 (N_5787,N_4442,N_3460);
or U5788 (N_5788,N_3276,N_3389);
nand U5789 (N_5789,N_3645,N_3089);
or U5790 (N_5790,N_3086,N_3576);
nor U5791 (N_5791,N_3438,N_3286);
xor U5792 (N_5792,N_3715,N_3530);
nor U5793 (N_5793,N_3250,N_4481);
xnor U5794 (N_5794,N_3874,N_3646);
or U5795 (N_5795,N_3611,N_3418);
nor U5796 (N_5796,N_4249,N_3330);
or U5797 (N_5797,N_3045,N_4087);
nand U5798 (N_5798,N_4132,N_3104);
xnor U5799 (N_5799,N_3753,N_4006);
or U5800 (N_5800,N_3598,N_3296);
nand U5801 (N_5801,N_3304,N_3291);
or U5802 (N_5802,N_3931,N_3510);
nand U5803 (N_5803,N_4107,N_3256);
xnor U5804 (N_5804,N_3424,N_3896);
xnor U5805 (N_5805,N_3206,N_3018);
xor U5806 (N_5806,N_3635,N_3427);
or U5807 (N_5807,N_3063,N_3639);
nand U5808 (N_5808,N_3436,N_3172);
nor U5809 (N_5809,N_3377,N_3133);
nand U5810 (N_5810,N_3614,N_3540);
nand U5811 (N_5811,N_4181,N_3359);
nand U5812 (N_5812,N_4496,N_3443);
xor U5813 (N_5813,N_4417,N_3078);
and U5814 (N_5814,N_3195,N_4357);
nand U5815 (N_5815,N_3413,N_3475);
xnor U5816 (N_5816,N_4447,N_3351);
xnor U5817 (N_5817,N_4105,N_3491);
nand U5818 (N_5818,N_3827,N_3121);
nand U5819 (N_5819,N_4484,N_4083);
xnor U5820 (N_5820,N_4491,N_3562);
nand U5821 (N_5821,N_3900,N_3563);
and U5822 (N_5822,N_3732,N_3265);
and U5823 (N_5823,N_3843,N_3771);
nand U5824 (N_5824,N_3176,N_4018);
or U5825 (N_5825,N_4470,N_3522);
nand U5826 (N_5826,N_3957,N_3379);
nor U5827 (N_5827,N_3315,N_3880);
and U5828 (N_5828,N_3599,N_4075);
or U5829 (N_5829,N_3460,N_3387);
nand U5830 (N_5830,N_3328,N_3500);
and U5831 (N_5831,N_3616,N_4455);
or U5832 (N_5832,N_3893,N_3530);
and U5833 (N_5833,N_4004,N_3464);
and U5834 (N_5834,N_3083,N_4160);
or U5835 (N_5835,N_3515,N_3160);
nand U5836 (N_5836,N_4100,N_4126);
and U5837 (N_5837,N_3872,N_3921);
nor U5838 (N_5838,N_3912,N_3210);
nand U5839 (N_5839,N_3046,N_4186);
nor U5840 (N_5840,N_3096,N_3847);
and U5841 (N_5841,N_3893,N_3129);
and U5842 (N_5842,N_3381,N_3858);
and U5843 (N_5843,N_3929,N_3033);
or U5844 (N_5844,N_3868,N_3072);
and U5845 (N_5845,N_4212,N_3852);
and U5846 (N_5846,N_3493,N_3313);
and U5847 (N_5847,N_3662,N_3296);
and U5848 (N_5848,N_3572,N_4067);
nor U5849 (N_5849,N_3434,N_3329);
and U5850 (N_5850,N_3643,N_3574);
and U5851 (N_5851,N_3414,N_4396);
or U5852 (N_5852,N_3513,N_4326);
or U5853 (N_5853,N_4442,N_4218);
nand U5854 (N_5854,N_3576,N_3912);
xor U5855 (N_5855,N_4112,N_3694);
and U5856 (N_5856,N_3624,N_3436);
xnor U5857 (N_5857,N_3909,N_3096);
nor U5858 (N_5858,N_3663,N_3477);
nor U5859 (N_5859,N_3098,N_3978);
and U5860 (N_5860,N_3396,N_3171);
or U5861 (N_5861,N_3956,N_4424);
nand U5862 (N_5862,N_3424,N_3376);
nand U5863 (N_5863,N_4355,N_3517);
or U5864 (N_5864,N_3246,N_3661);
or U5865 (N_5865,N_3498,N_4378);
and U5866 (N_5866,N_4095,N_3596);
and U5867 (N_5867,N_3045,N_4496);
nor U5868 (N_5868,N_3196,N_3027);
xnor U5869 (N_5869,N_4309,N_3616);
nor U5870 (N_5870,N_4059,N_4202);
nor U5871 (N_5871,N_3164,N_3699);
and U5872 (N_5872,N_4367,N_3661);
or U5873 (N_5873,N_3601,N_4308);
nand U5874 (N_5874,N_3637,N_3173);
nor U5875 (N_5875,N_3129,N_3924);
xnor U5876 (N_5876,N_4094,N_3025);
nor U5877 (N_5877,N_3673,N_4227);
nand U5878 (N_5878,N_4445,N_4195);
and U5879 (N_5879,N_3283,N_4485);
nand U5880 (N_5880,N_3352,N_3091);
or U5881 (N_5881,N_4042,N_3882);
nor U5882 (N_5882,N_3963,N_3466);
xnor U5883 (N_5883,N_3999,N_4198);
nand U5884 (N_5884,N_4035,N_4429);
xnor U5885 (N_5885,N_3507,N_4043);
xor U5886 (N_5886,N_3041,N_3965);
nand U5887 (N_5887,N_4126,N_4041);
nor U5888 (N_5888,N_3605,N_4309);
and U5889 (N_5889,N_4248,N_3084);
xnor U5890 (N_5890,N_3103,N_3898);
nand U5891 (N_5891,N_4194,N_3129);
xor U5892 (N_5892,N_3354,N_3281);
nand U5893 (N_5893,N_4119,N_3778);
or U5894 (N_5894,N_4092,N_3696);
or U5895 (N_5895,N_3800,N_3743);
or U5896 (N_5896,N_3105,N_4481);
xor U5897 (N_5897,N_3024,N_3153);
nor U5898 (N_5898,N_3662,N_4206);
and U5899 (N_5899,N_3463,N_3814);
xnor U5900 (N_5900,N_3298,N_4015);
and U5901 (N_5901,N_4362,N_3596);
and U5902 (N_5902,N_3306,N_3463);
xor U5903 (N_5903,N_3686,N_3599);
and U5904 (N_5904,N_3989,N_4440);
or U5905 (N_5905,N_3239,N_4065);
xor U5906 (N_5906,N_3475,N_4473);
xor U5907 (N_5907,N_3057,N_3414);
and U5908 (N_5908,N_4246,N_3464);
nand U5909 (N_5909,N_4144,N_3341);
or U5910 (N_5910,N_4078,N_3873);
nand U5911 (N_5911,N_3674,N_3815);
xnor U5912 (N_5912,N_3499,N_3863);
and U5913 (N_5913,N_3720,N_3254);
and U5914 (N_5914,N_3627,N_3457);
and U5915 (N_5915,N_3647,N_3047);
or U5916 (N_5916,N_3623,N_4432);
or U5917 (N_5917,N_3953,N_3913);
nand U5918 (N_5918,N_4351,N_4034);
nand U5919 (N_5919,N_4324,N_3437);
xor U5920 (N_5920,N_3464,N_3145);
or U5921 (N_5921,N_4158,N_3082);
and U5922 (N_5922,N_3328,N_3501);
xnor U5923 (N_5923,N_3290,N_4237);
and U5924 (N_5924,N_4232,N_3624);
nand U5925 (N_5925,N_4126,N_3936);
nand U5926 (N_5926,N_3293,N_3825);
or U5927 (N_5927,N_4066,N_3581);
and U5928 (N_5928,N_3719,N_3671);
or U5929 (N_5929,N_3005,N_3543);
nor U5930 (N_5930,N_3923,N_4196);
or U5931 (N_5931,N_3500,N_4135);
nor U5932 (N_5932,N_4497,N_3807);
and U5933 (N_5933,N_3245,N_3611);
nor U5934 (N_5934,N_3676,N_4116);
or U5935 (N_5935,N_3217,N_3719);
xnor U5936 (N_5936,N_3639,N_4234);
xnor U5937 (N_5937,N_3308,N_3418);
or U5938 (N_5938,N_4355,N_4229);
xor U5939 (N_5939,N_4468,N_3606);
xor U5940 (N_5940,N_4035,N_3029);
and U5941 (N_5941,N_4145,N_3798);
and U5942 (N_5942,N_3527,N_3846);
nor U5943 (N_5943,N_3453,N_4357);
and U5944 (N_5944,N_4107,N_4141);
xnor U5945 (N_5945,N_3072,N_3608);
and U5946 (N_5946,N_4129,N_3500);
xnor U5947 (N_5947,N_4323,N_3099);
nor U5948 (N_5948,N_4115,N_4022);
and U5949 (N_5949,N_3293,N_4326);
xor U5950 (N_5950,N_4303,N_3171);
nand U5951 (N_5951,N_3189,N_4190);
and U5952 (N_5952,N_4220,N_4109);
and U5953 (N_5953,N_4274,N_4183);
xnor U5954 (N_5954,N_3923,N_4407);
xor U5955 (N_5955,N_3549,N_4061);
and U5956 (N_5956,N_3515,N_3258);
or U5957 (N_5957,N_4060,N_4318);
xnor U5958 (N_5958,N_4084,N_4157);
or U5959 (N_5959,N_3467,N_3369);
nor U5960 (N_5960,N_4207,N_3754);
and U5961 (N_5961,N_4089,N_3119);
nor U5962 (N_5962,N_4332,N_3087);
xor U5963 (N_5963,N_3344,N_4221);
nor U5964 (N_5964,N_3859,N_4318);
or U5965 (N_5965,N_3407,N_3119);
or U5966 (N_5966,N_4107,N_4185);
nor U5967 (N_5967,N_3512,N_3176);
or U5968 (N_5968,N_4367,N_4052);
or U5969 (N_5969,N_3042,N_3238);
nand U5970 (N_5970,N_3634,N_3847);
nand U5971 (N_5971,N_3242,N_4423);
nand U5972 (N_5972,N_4496,N_3219);
nor U5973 (N_5973,N_3396,N_4240);
nand U5974 (N_5974,N_4272,N_4135);
nor U5975 (N_5975,N_4237,N_4164);
nor U5976 (N_5976,N_4223,N_3454);
nor U5977 (N_5977,N_3053,N_4073);
nand U5978 (N_5978,N_4202,N_3951);
nor U5979 (N_5979,N_3916,N_3774);
nor U5980 (N_5980,N_3965,N_3668);
or U5981 (N_5981,N_4152,N_3550);
xor U5982 (N_5982,N_3568,N_3091);
xor U5983 (N_5983,N_3473,N_3189);
or U5984 (N_5984,N_3194,N_4454);
or U5985 (N_5985,N_3136,N_4324);
nand U5986 (N_5986,N_3261,N_3663);
nor U5987 (N_5987,N_4416,N_4102);
xor U5988 (N_5988,N_3057,N_4194);
nand U5989 (N_5989,N_3073,N_3579);
or U5990 (N_5990,N_3492,N_3398);
and U5991 (N_5991,N_4083,N_3223);
nor U5992 (N_5992,N_4491,N_3439);
nand U5993 (N_5993,N_3264,N_4137);
xnor U5994 (N_5994,N_3608,N_4191);
or U5995 (N_5995,N_3979,N_4069);
and U5996 (N_5996,N_3711,N_3397);
nor U5997 (N_5997,N_3672,N_3890);
and U5998 (N_5998,N_3184,N_3690);
nand U5999 (N_5999,N_4415,N_3571);
xor U6000 (N_6000,N_4687,N_5896);
or U6001 (N_6001,N_5524,N_4757);
and U6002 (N_6002,N_5888,N_4630);
nand U6003 (N_6003,N_5572,N_4994);
nand U6004 (N_6004,N_4552,N_5265);
or U6005 (N_6005,N_5249,N_5085);
or U6006 (N_6006,N_5640,N_4566);
and U6007 (N_6007,N_4990,N_5660);
nor U6008 (N_6008,N_4707,N_5676);
xor U6009 (N_6009,N_5732,N_5961);
or U6010 (N_6010,N_4570,N_5080);
and U6011 (N_6011,N_5028,N_5232);
nand U6012 (N_6012,N_4634,N_5526);
nand U6013 (N_6013,N_5536,N_5221);
and U6014 (N_6014,N_5932,N_4938);
xor U6015 (N_6015,N_5656,N_5495);
nor U6016 (N_6016,N_5725,N_4815);
nand U6017 (N_6017,N_5943,N_4802);
xnor U6018 (N_6018,N_5513,N_4653);
nand U6019 (N_6019,N_5955,N_4655);
nor U6020 (N_6020,N_5785,N_4624);
or U6021 (N_6021,N_4638,N_4889);
nor U6022 (N_6022,N_4706,N_5662);
or U6023 (N_6023,N_4539,N_5523);
xnor U6024 (N_6024,N_5542,N_4523);
nand U6025 (N_6025,N_5702,N_5328);
and U6026 (N_6026,N_4750,N_4525);
nor U6027 (N_6027,N_5677,N_5100);
nor U6028 (N_6028,N_5819,N_5670);
or U6029 (N_6029,N_4897,N_5113);
or U6030 (N_6030,N_5557,N_4536);
and U6031 (N_6031,N_5000,N_5515);
xnor U6032 (N_6032,N_4722,N_5522);
xnor U6033 (N_6033,N_5307,N_5021);
and U6034 (N_6034,N_5652,N_5477);
xor U6035 (N_6035,N_4509,N_4919);
xnor U6036 (N_6036,N_5146,N_4907);
and U6037 (N_6037,N_5108,N_5438);
nor U6038 (N_6038,N_4720,N_5479);
nor U6039 (N_6039,N_4542,N_4654);
and U6040 (N_6040,N_5290,N_4648);
nor U6041 (N_6041,N_4515,N_5376);
or U6042 (N_6042,N_5134,N_5775);
nand U6043 (N_6043,N_5626,N_5433);
or U6044 (N_6044,N_5855,N_5255);
nor U6045 (N_6045,N_4874,N_5997);
or U6046 (N_6046,N_4927,N_5747);
xnor U6047 (N_6047,N_5447,N_5288);
or U6048 (N_6048,N_5074,N_5608);
nor U6049 (N_6049,N_4752,N_5800);
nor U6050 (N_6050,N_4824,N_5944);
or U6051 (N_6051,N_4605,N_5794);
nand U6052 (N_6052,N_5805,N_4916);
or U6053 (N_6053,N_4558,N_5658);
xor U6054 (N_6054,N_5500,N_5415);
nor U6055 (N_6055,N_5029,N_5234);
nand U6056 (N_6056,N_5107,N_5575);
and U6057 (N_6057,N_5865,N_4691);
nand U6058 (N_6058,N_5262,N_4579);
and U6059 (N_6059,N_4773,N_5068);
or U6060 (N_6060,N_5580,N_5009);
xor U6061 (N_6061,N_5215,N_5365);
nand U6062 (N_6062,N_4697,N_5701);
or U6063 (N_6063,N_5091,N_4950);
or U6064 (N_6064,N_4686,N_5514);
xor U6065 (N_6065,N_5468,N_5231);
or U6066 (N_6066,N_4556,N_5030);
and U6067 (N_6067,N_5271,N_4991);
or U6068 (N_6068,N_5366,N_5304);
nor U6069 (N_6069,N_4729,N_5518);
or U6070 (N_6070,N_5168,N_5082);
and U6071 (N_6071,N_4788,N_5097);
nor U6072 (N_6072,N_5179,N_4678);
or U6073 (N_6073,N_4786,N_5527);
nor U6074 (N_6074,N_5666,N_4977);
xor U6075 (N_6075,N_4577,N_5213);
xnor U6076 (N_6076,N_5472,N_5566);
or U6077 (N_6077,N_4547,N_4585);
nor U6078 (N_6078,N_5564,N_5382);
nor U6079 (N_6079,N_5037,N_5594);
or U6080 (N_6080,N_4898,N_5745);
xor U6081 (N_6081,N_4856,N_4762);
and U6082 (N_6082,N_5857,N_5095);
and U6083 (N_6083,N_5501,N_5109);
and U6084 (N_6084,N_4533,N_4761);
nor U6085 (N_6085,N_5154,N_5996);
and U6086 (N_6086,N_5435,N_4896);
xor U6087 (N_6087,N_5467,N_4621);
or U6088 (N_6088,N_5749,N_4971);
and U6089 (N_6089,N_4951,N_4915);
nor U6090 (N_6090,N_4668,N_5295);
xor U6091 (N_6091,N_5671,N_4727);
and U6092 (N_6092,N_5899,N_5807);
or U6093 (N_6093,N_5511,N_5458);
or U6094 (N_6094,N_5986,N_5088);
and U6095 (N_6095,N_5563,N_5610);
xnor U6096 (N_6096,N_5486,N_5678);
nor U6097 (N_6097,N_4740,N_5416);
nand U6098 (N_6098,N_5494,N_5320);
nand U6099 (N_6099,N_4666,N_4918);
nand U6100 (N_6100,N_4625,N_5145);
nand U6101 (N_6101,N_5436,N_5434);
nor U6102 (N_6102,N_5769,N_5343);
nand U6103 (N_6103,N_4689,N_5727);
or U6104 (N_6104,N_5103,N_5070);
or U6105 (N_6105,N_5872,N_5457);
nor U6106 (N_6106,N_5776,N_5164);
nor U6107 (N_6107,N_4510,N_5904);
and U6108 (N_6108,N_4700,N_4812);
nand U6109 (N_6109,N_4578,N_5668);
nor U6110 (N_6110,N_5974,N_5998);
nor U6111 (N_6111,N_4755,N_5182);
nand U6112 (N_6112,N_4917,N_5561);
nand U6113 (N_6113,N_4775,N_5260);
xnor U6114 (N_6114,N_4586,N_5814);
nor U6115 (N_6115,N_5019,N_5310);
and U6116 (N_6116,N_5317,N_4572);
and U6117 (N_6117,N_4945,N_4767);
or U6118 (N_6118,N_4692,N_5667);
nor U6119 (N_6119,N_4592,N_5528);
nor U6120 (N_6120,N_5659,N_5636);
nand U6121 (N_6121,N_5560,N_4575);
nand U6122 (N_6122,N_4795,N_4986);
or U6123 (N_6123,N_5717,N_5399);
and U6124 (N_6124,N_4695,N_5426);
and U6125 (N_6125,N_4804,N_5918);
xor U6126 (N_6126,N_4837,N_5346);
nand U6127 (N_6127,N_5350,N_5084);
xnor U6128 (N_6128,N_5933,N_5485);
nor U6129 (N_6129,N_5245,N_4679);
and U6130 (N_6130,N_4979,N_5173);
or U6131 (N_6131,N_4742,N_4635);
and U6132 (N_6132,N_4800,N_5614);
or U6133 (N_6133,N_5598,N_5469);
and U6134 (N_6134,N_4664,N_4739);
nor U6135 (N_6135,N_4535,N_4846);
nor U6136 (N_6136,N_5367,N_4589);
and U6137 (N_6137,N_5694,N_4975);
and U6138 (N_6138,N_5691,N_5430);
and U6139 (N_6139,N_5568,N_5770);
or U6140 (N_6140,N_4870,N_5272);
nor U6141 (N_6141,N_5554,N_4816);
or U6142 (N_6142,N_5424,N_4628);
and U6143 (N_6143,N_5064,N_5230);
xnor U6144 (N_6144,N_5228,N_4763);
nand U6145 (N_6145,N_4796,N_5651);
and U6146 (N_6146,N_5870,N_4829);
or U6147 (N_6147,N_5291,N_5593);
xor U6148 (N_6148,N_4892,N_5060);
nor U6149 (N_6149,N_5199,N_5178);
and U6150 (N_6150,N_5360,N_4885);
and U6151 (N_6151,N_4964,N_4963);
and U6152 (N_6152,N_5650,N_5908);
or U6153 (N_6153,N_4574,N_5952);
xor U6154 (N_6154,N_4561,N_5045);
and U6155 (N_6155,N_4873,N_4580);
and U6156 (N_6156,N_4583,N_5102);
or U6157 (N_6157,N_5076,N_4908);
nand U6158 (N_6158,N_5374,N_4582);
nor U6159 (N_6159,N_5638,N_4617);
nand U6160 (N_6160,N_5259,N_5569);
nand U6161 (N_6161,N_4526,N_5675);
nor U6162 (N_6162,N_5244,N_5451);
xor U6163 (N_6163,N_5333,N_5497);
and U6164 (N_6164,N_5251,N_5789);
and U6165 (N_6165,N_4598,N_5622);
or U6166 (N_6166,N_4719,N_5128);
and U6167 (N_6167,N_5861,N_5099);
and U6168 (N_6168,N_5864,N_5700);
and U6169 (N_6169,N_5852,N_5959);
and U6170 (N_6170,N_5512,N_5979);
xnor U6171 (N_6171,N_5792,N_4808);
or U6172 (N_6172,N_5395,N_5689);
or U6173 (N_6173,N_4973,N_4982);
and U6174 (N_6174,N_5254,N_5981);
nor U6175 (N_6175,N_5001,N_4925);
nor U6176 (N_6176,N_5879,N_5545);
xor U6177 (N_6177,N_5552,N_4886);
xnor U6178 (N_6178,N_5321,N_5628);
and U6179 (N_6179,N_5408,N_4685);
nand U6180 (N_6180,N_5589,N_5993);
xnor U6181 (N_6181,N_5302,N_5850);
nor U6182 (N_6182,N_5577,N_5474);
nor U6183 (N_6183,N_4759,N_5696);
nand U6184 (N_6184,N_4772,N_5236);
or U6185 (N_6185,N_4677,N_5003);
or U6186 (N_6186,N_5724,N_4869);
nor U6187 (N_6187,N_5410,N_4545);
or U6188 (N_6188,N_5369,N_5753);
or U6189 (N_6189,N_4968,N_5046);
xnor U6190 (N_6190,N_5115,N_5038);
nor U6191 (N_6191,N_5830,N_5983);
or U6192 (N_6192,N_5277,N_5726);
xor U6193 (N_6193,N_4576,N_5218);
nand U6194 (N_6194,N_4616,N_5853);
nand U6195 (N_6195,N_5773,N_4731);
xnor U6196 (N_6196,N_4553,N_5894);
and U6197 (N_6197,N_5263,N_4735);
or U6198 (N_6198,N_5345,N_5750);
nor U6199 (N_6199,N_4513,N_5687);
or U6200 (N_6200,N_4820,N_5197);
xnor U6201 (N_6201,N_5686,N_4953);
and U6202 (N_6202,N_4828,N_5849);
and U6203 (N_6203,N_5371,N_5840);
or U6204 (N_6204,N_5499,N_5869);
nor U6205 (N_6205,N_5062,N_4832);
and U6206 (N_6206,N_5484,N_4665);
and U6207 (N_6207,N_5239,N_5897);
and U6208 (N_6208,N_5657,N_4976);
xor U6209 (N_6209,N_5616,N_4882);
xor U6210 (N_6210,N_4987,N_5842);
or U6211 (N_6211,N_4784,N_5205);
nor U6212 (N_6212,N_5402,N_5643);
nor U6213 (N_6213,N_5962,N_5264);
nand U6214 (N_6214,N_5252,N_4924);
and U6215 (N_6215,N_5803,N_4659);
xor U6216 (N_6216,N_4657,N_5148);
nand U6217 (N_6217,N_5363,N_5565);
nand U6218 (N_6218,N_5692,N_5682);
nand U6219 (N_6219,N_5034,N_5836);
nand U6220 (N_6220,N_4878,N_5621);
and U6221 (N_6221,N_5703,N_5344);
nor U6222 (N_6222,N_4920,N_5892);
nand U6223 (N_6223,N_5556,N_4534);
or U6224 (N_6224,N_4839,N_5300);
xnor U6225 (N_6225,N_5308,N_5229);
nand U6226 (N_6226,N_5324,N_5942);
nand U6227 (N_6227,N_5914,N_5601);
nand U6228 (N_6228,N_5570,N_5496);
nor U6229 (N_6229,N_5920,N_4753);
or U6230 (N_6230,N_5939,N_5127);
nand U6231 (N_6231,N_5118,N_5665);
or U6232 (N_6232,N_5152,N_5664);
and U6233 (N_6233,N_4627,N_4922);
nand U6234 (N_6234,N_4849,N_4588);
xor U6235 (N_6235,N_5466,N_4875);
and U6236 (N_6236,N_5715,N_5210);
nor U6237 (N_6237,N_5829,N_5209);
xnor U6238 (N_6238,N_5279,N_5149);
nor U6239 (N_6239,N_4939,N_4955);
and U6240 (N_6240,N_5446,N_4777);
nand U6241 (N_6241,N_5900,N_5768);
nand U6242 (N_6242,N_5699,N_4745);
or U6243 (N_6243,N_4946,N_5609);
nor U6244 (N_6244,N_4765,N_5673);
nor U6245 (N_6245,N_5804,N_5809);
nand U6246 (N_6246,N_4614,N_4854);
or U6247 (N_6247,N_5404,N_4704);
or U6248 (N_6248,N_5298,N_5889);
nor U6249 (N_6249,N_4969,N_4607);
nand U6250 (N_6250,N_5340,N_4768);
and U6251 (N_6251,N_5826,N_4805);
nand U6252 (N_6252,N_5355,N_4684);
xnor U6253 (N_6253,N_4997,N_5916);
xor U6254 (N_6254,N_5086,N_5688);
or U6255 (N_6255,N_5016,N_5846);
xnor U6256 (N_6256,N_5719,N_4587);
or U6257 (N_6257,N_4967,N_5132);
or U6258 (N_6258,N_5112,N_5860);
nand U6259 (N_6259,N_4629,N_5007);
nor U6260 (N_6260,N_4673,N_5931);
or U6261 (N_6261,N_5690,N_5206);
or U6262 (N_6262,N_4505,N_5631);
or U6263 (N_6263,N_5772,N_4749);
or U6264 (N_6264,N_4632,N_5220);
or U6265 (N_6265,N_5192,N_5641);
and U6266 (N_6266,N_5353,N_5764);
and U6267 (N_6267,N_4728,N_5645);
xor U6268 (N_6268,N_5875,N_5247);
nor U6269 (N_6269,N_4845,N_5758);
nand U6270 (N_6270,N_5823,N_5352);
nor U6271 (N_6271,N_5031,N_5937);
and U6272 (N_6272,N_5450,N_5827);
nor U6273 (N_6273,N_5123,N_5165);
xor U6274 (N_6274,N_5493,N_5788);
nor U6275 (N_6275,N_5393,N_4543);
nor U6276 (N_6276,N_5716,N_4880);
nor U6277 (N_6277,N_4817,N_5384);
xnor U6278 (N_6278,N_4980,N_5967);
nor U6279 (N_6279,N_4903,N_4709);
nor U6280 (N_6280,N_5743,N_5073);
xnor U6281 (N_6281,N_4890,N_5443);
and U6282 (N_6282,N_4738,N_5377);
and U6283 (N_6283,N_5323,N_4966);
and U6284 (N_6284,N_5059,N_5005);
or U6285 (N_6285,N_4952,N_5379);
and U6286 (N_6286,N_5613,N_5521);
or U6287 (N_6287,N_4511,N_4876);
nor U6288 (N_6288,N_5627,N_5481);
xor U6289 (N_6289,N_4974,N_5297);
or U6290 (N_6290,N_5736,N_5212);
xnor U6291 (N_6291,N_4642,N_5175);
and U6292 (N_6292,N_5011,N_4996);
or U6293 (N_6293,N_5306,N_4544);
and U6294 (N_6294,N_5120,N_4581);
or U6295 (N_6295,N_5487,N_5780);
xor U6296 (N_6296,N_5498,N_5417);
and U6297 (N_6297,N_5588,N_5624);
nand U6298 (N_6298,N_5358,N_4887);
nor U6299 (N_6299,N_4895,N_5448);
xor U6300 (N_6300,N_5698,N_5002);
and U6301 (N_6301,N_5280,N_5964);
nor U6302 (N_6302,N_5817,N_5760);
nand U6303 (N_6303,N_5305,N_5562);
nor U6304 (N_6304,N_5378,N_5876);
nor U6305 (N_6305,N_5380,N_4758);
nor U6306 (N_6306,N_5111,N_5948);
nand U6307 (N_6307,N_4502,N_4944);
nand U6308 (N_6308,N_4913,N_4520);
and U6309 (N_6309,N_5880,N_4822);
nand U6310 (N_6310,N_5611,N_5543);
xnor U6311 (N_6311,N_5439,N_4711);
nand U6312 (N_6312,N_4848,N_5982);
nand U6313 (N_6313,N_4743,N_5226);
or U6314 (N_6314,N_4597,N_4584);
nor U6315 (N_6315,N_4965,N_5414);
and U6316 (N_6316,N_5381,N_4970);
nor U6317 (N_6317,N_5824,N_5821);
xor U6318 (N_6318,N_4670,N_5537);
xnor U6319 (N_6319,N_5603,N_5143);
xnor U6320 (N_6320,N_5705,N_5394);
or U6321 (N_6321,N_5104,N_4741);
or U6322 (N_6322,N_5928,N_5261);
xnor U6323 (N_6323,N_5845,N_5375);
nor U6324 (N_6324,N_5273,N_5584);
or U6325 (N_6325,N_5695,N_4599);
or U6326 (N_6326,N_5035,N_5223);
and U6327 (N_6327,N_5093,N_5738);
and U6328 (N_6328,N_5746,N_5359);
nor U6329 (N_6329,N_4516,N_4782);
xnor U6330 (N_6330,N_5924,N_5480);
or U6331 (N_6331,N_5189,N_5759);
xnor U6332 (N_6332,N_5604,N_4732);
nor U6333 (N_6333,N_4703,N_5440);
or U6334 (N_6334,N_5462,N_4864);
nand U6335 (N_6335,N_5079,N_5503);
or U6336 (N_6336,N_5482,N_5058);
nand U6337 (N_6337,N_5599,N_5765);
xnor U6338 (N_6338,N_5219,N_5409);
or U6339 (N_6339,N_5276,N_5141);
and U6340 (N_6340,N_5548,N_4960);
or U6341 (N_6341,N_5217,N_5704);
xor U6342 (N_6342,N_5941,N_5190);
xor U6343 (N_6343,N_5634,N_4676);
and U6344 (N_6344,N_5832,N_5573);
xnor U6345 (N_6345,N_4891,N_5015);
nand U6346 (N_6346,N_4540,N_5200);
nand U6347 (N_6347,N_5831,N_4603);
nor U6348 (N_6348,N_5157,N_5714);
nand U6349 (N_6349,N_4571,N_5327);
xnor U6350 (N_6350,N_4904,N_4754);
xor U6351 (N_6351,N_5401,N_5054);
and U6352 (N_6352,N_4797,N_5301);
nor U6353 (N_6353,N_5017,N_5799);
or U6354 (N_6354,N_5114,N_5354);
xnor U6355 (N_6355,N_5762,N_5072);
xor U6356 (N_6356,N_4636,N_5946);
or U6357 (N_6357,N_4914,N_4830);
and U6358 (N_6358,N_4569,N_4923);
xnor U6359 (N_6359,N_5936,N_4613);
xor U6360 (N_6360,N_4730,N_4995);
xnor U6361 (N_6361,N_5216,N_5225);
xor U6362 (N_6362,N_4734,N_5110);
nand U6363 (N_6363,N_5950,N_4529);
nor U6364 (N_6364,N_5470,N_5293);
nand U6365 (N_6365,N_5984,N_4984);
xnor U6366 (N_6366,N_5158,N_5018);
nor U6367 (N_6367,N_5923,N_5096);
nand U6368 (N_6368,N_5203,N_5407);
nor U6369 (N_6369,N_5287,N_4658);
nand U6370 (N_6370,N_5661,N_5449);
nand U6371 (N_6371,N_5286,N_5131);
and U6372 (N_6372,N_5196,N_5619);
nand U6373 (N_6373,N_5090,N_4921);
nor U6374 (N_6374,N_5331,N_5442);
xnor U6375 (N_6375,N_4751,N_4524);
and U6376 (N_6376,N_4959,N_4690);
and U6377 (N_6377,N_5796,N_4942);
nor U6378 (N_6378,N_5629,N_5253);
nor U6379 (N_6379,N_5866,N_5957);
nor U6380 (N_6380,N_5510,N_5319);
nand U6381 (N_6381,N_4948,N_5309);
nor U6382 (N_6382,N_5910,N_5071);
and U6383 (N_6383,N_4855,N_5383);
xor U6384 (N_6384,N_4541,N_5362);
nand U6385 (N_6385,N_4562,N_5140);
or U6386 (N_6386,N_5930,N_5534);
nand U6387 (N_6387,N_4860,N_5684);
nor U6388 (N_6388,N_4881,N_4811);
or U6389 (N_6389,N_5151,N_5050);
and U6390 (N_6390,N_5387,N_5585);
nor U6391 (N_6391,N_5742,N_5533);
and U6392 (N_6392,N_5597,N_5135);
nand U6393 (N_6393,N_5198,N_4660);
nor U6394 (N_6394,N_5739,N_5248);
and U6395 (N_6395,N_4593,N_5063);
nor U6396 (N_6396,N_5010,N_5623);
and U6397 (N_6397,N_4550,N_4500);
xor U6398 (N_6398,N_4650,N_4956);
or U6399 (N_6399,N_5405,N_5706);
nand U6400 (N_6400,N_4834,N_5989);
xnor U6401 (N_6401,N_5756,N_4705);
nor U6402 (N_6402,N_4647,N_4862);
and U6403 (N_6403,N_5774,N_5771);
xor U6404 (N_6404,N_4929,N_4568);
nor U6405 (N_6405,N_5184,N_5122);
nor U6406 (N_6406,N_5825,N_5389);
nor U6407 (N_6407,N_5283,N_4610);
nor U6408 (N_6408,N_5427,N_5318);
and U6409 (N_6409,N_5988,N_5160);
nor U6410 (N_6410,N_4675,N_4954);
nand U6411 (N_6411,N_5325,N_5605);
nand U6412 (N_6412,N_5454,N_5057);
xor U6413 (N_6413,N_4626,N_4501);
nand U6414 (N_6414,N_4620,N_4936);
or U6415 (N_6415,N_5195,N_5553);
nand U6416 (N_6416,N_5047,N_5453);
nand U6417 (N_6417,N_5579,N_5246);
or U6418 (N_6418,N_5403,N_5761);
nor U6419 (N_6419,N_4644,N_4601);
or U6420 (N_6420,N_5654,N_5284);
or U6421 (N_6421,N_5207,N_4883);
nor U6422 (N_6422,N_4615,N_4604);
xnor U6423 (N_6423,N_5476,N_4667);
or U6424 (N_6424,N_5183,N_4827);
nand U6425 (N_6425,N_5722,N_5538);
and U6426 (N_6426,N_5927,N_5567);
or U6427 (N_6427,N_5180,N_5364);
and U6428 (N_6428,N_5459,N_4872);
nor U6429 (N_6429,N_5004,N_4910);
and U6430 (N_6430,N_4721,N_5546);
xor U6431 (N_6431,N_5400,N_5419);
nand U6432 (N_6432,N_4645,N_4859);
nor U6433 (N_6433,N_5491,N_5890);
nor U6434 (N_6434,N_5332,N_5951);
or U6435 (N_6435,N_4714,N_5994);
and U6436 (N_6436,N_5445,N_5990);
and U6437 (N_6437,N_5532,N_5844);
nand U6438 (N_6438,N_5066,N_5867);
xnor U6439 (N_6439,N_5956,N_4527);
or U6440 (N_6440,N_5390,N_5874);
and U6441 (N_6441,N_5294,N_5036);
or U6442 (N_6442,N_5922,N_5171);
xnor U6443 (N_6443,N_5653,N_4712);
xor U6444 (N_6444,N_4672,N_5478);
xnor U6445 (N_6445,N_5707,N_5793);
nand U6446 (N_6446,N_4789,N_5540);
nand U6447 (N_6447,N_4631,N_4850);
nand U6448 (N_6448,N_5816,N_4560);
nand U6449 (N_6449,N_5966,N_5349);
nor U6450 (N_6450,N_4770,N_5361);
nand U6451 (N_6451,N_5155,N_5884);
xor U6452 (N_6452,N_5517,N_4640);
xnor U6453 (N_6453,N_5547,N_5710);
or U6454 (N_6454,N_4698,N_4867);
xnor U6455 (N_6455,N_5336,N_5602);
nand U6456 (N_6456,N_4937,N_5708);
nor U6457 (N_6457,N_5337,N_4844);
and U6458 (N_6458,N_5863,N_5181);
and U6459 (N_6459,N_5473,N_5663);
xnor U6460 (N_6460,N_4787,N_4746);
nor U6461 (N_6461,N_5783,N_5136);
and U6462 (N_6462,N_5737,N_5834);
nand U6463 (N_6463,N_4514,N_4551);
xnor U6464 (N_6464,N_5881,N_4681);
nand U6465 (N_6465,N_5963,N_5329);
and U6466 (N_6466,N_5452,N_5620);
nand U6467 (N_6467,N_5420,N_5335);
and U6468 (N_6468,N_4791,N_5960);
nand U6469 (N_6469,N_5999,N_5680);
or U6470 (N_6470,N_5648,N_4671);
or U6471 (N_6471,N_5392,N_5672);
xnor U6472 (N_6472,N_4663,N_4798);
or U6473 (N_6473,N_5023,N_5437);
nand U6474 (N_6474,N_5559,N_5887);
nand U6475 (N_6475,N_5921,N_4662);
xor U6476 (N_6476,N_5975,N_5583);
nand U6477 (N_6477,N_5505,N_4957);
xnor U6478 (N_6478,N_4785,N_5388);
xor U6479 (N_6479,N_4972,N_4733);
nor U6480 (N_6480,N_4508,N_4884);
nor U6481 (N_6481,N_5893,N_5578);
or U6482 (N_6482,N_5529,N_4652);
or U6483 (N_6483,N_5766,N_4764);
nor U6484 (N_6484,N_5778,N_5065);
nand U6485 (N_6485,N_4776,N_5041);
or U6486 (N_6486,N_5242,N_4926);
nand U6487 (N_6487,N_5506,N_4522);
xnor U6488 (N_6488,N_4682,N_5551);
nand U6489 (N_6489,N_5617,N_4517);
or U6490 (N_6490,N_4622,N_5782);
nand U6491 (N_6491,N_5460,N_5275);
or U6492 (N_6492,N_5976,N_5531);
nand U6493 (N_6493,N_5649,N_5509);
nand U6494 (N_6494,N_5733,N_5056);
and U6495 (N_6495,N_5592,N_4899);
nand U6496 (N_6496,N_5822,N_5233);
nor U6497 (N_6497,N_5754,N_5740);
nand U6498 (N_6498,N_5185,N_5464);
and U6499 (N_6499,N_5644,N_5815);
or U6500 (N_6500,N_4894,N_5397);
and U6501 (N_6501,N_5075,N_5891);
nand U6502 (N_6502,N_4530,N_4669);
xnor U6503 (N_6503,N_5587,N_5257);
nor U6504 (N_6504,N_5237,N_4934);
nor U6505 (N_6505,N_4737,N_5615);
nor U6506 (N_6506,N_5126,N_4813);
and U6507 (N_6507,N_5877,N_5954);
nor U6508 (N_6508,N_4774,N_5808);
or U6509 (N_6509,N_5373,N_5646);
or U6510 (N_6510,N_5625,N_4866);
xor U6511 (N_6511,N_5838,N_4983);
nand U6512 (N_6512,N_5847,N_4993);
and U6513 (N_6513,N_5167,N_5348);
nor U6514 (N_6514,N_5049,N_5590);
xnor U6515 (N_6515,N_5087,N_5431);
or U6516 (N_6516,N_5813,N_5618);
nor U6517 (N_6517,N_5681,N_4641);
nand U6518 (N_6518,N_5256,N_5441);
nor U6519 (N_6519,N_5292,N_4949);
nand U6520 (N_6520,N_5632,N_5856);
xnor U6521 (N_6521,N_5882,N_5790);
and U6522 (N_6522,N_5006,N_5061);
or U6523 (N_6523,N_5530,N_5266);
nand U6524 (N_6524,N_5633,N_4555);
nor U6525 (N_6525,N_4747,N_5269);
xor U6526 (N_6526,N_5465,N_5227);
nor U6527 (N_6527,N_4595,N_4546);
nand U6528 (N_6528,N_5784,N_4879);
and U6529 (N_6529,N_4748,N_5069);
nand U6530 (N_6530,N_5843,N_5600);
xnor U6531 (N_6531,N_5092,N_4590);
nand U6532 (N_6532,N_5461,N_4718);
nand U6533 (N_6533,N_4888,N_5683);
xor U6534 (N_6534,N_5422,N_4809);
and U6535 (N_6535,N_5925,N_4861);
xnor U6536 (N_6536,N_5008,N_5905);
or U6537 (N_6537,N_4736,N_4868);
nor U6538 (N_6538,N_5385,N_5341);
and U6539 (N_6539,N_5903,N_5787);
nor U6540 (N_6540,N_4688,N_4702);
xor U6541 (N_6541,N_5033,N_4619);
nand U6542 (N_6542,N_4573,N_5238);
and U6543 (N_6543,N_4793,N_5083);
xor U6544 (N_6544,N_5098,N_5044);
nor U6545 (N_6545,N_4760,N_5915);
and U6546 (N_6546,N_5406,N_5987);
nand U6547 (N_6547,N_4708,N_5444);
xnor U6548 (N_6548,N_4988,N_5767);
or U6549 (N_6549,N_5596,N_4778);
and U6550 (N_6550,N_5456,N_5917);
and U6551 (N_6551,N_5368,N_5637);
or U6552 (N_6552,N_4715,N_5516);
or U6553 (N_6553,N_5992,N_4978);
or U6554 (N_6554,N_5906,N_5243);
nor U6555 (N_6555,N_4528,N_5878);
and U6556 (N_6556,N_5119,N_5851);
nand U6557 (N_6557,N_4699,N_4701);
or U6558 (N_6558,N_4506,N_5347);
nand U6559 (N_6559,N_5818,N_5868);
nand U6560 (N_6560,N_5755,N_4600);
nor U6561 (N_6561,N_4853,N_5968);
or U6562 (N_6562,N_4548,N_4962);
nor U6563 (N_6563,N_5334,N_4680);
nand U6564 (N_6564,N_4559,N_5525);
or U6565 (N_6565,N_4639,N_5170);
and U6566 (N_6566,N_5728,N_4637);
and U6567 (N_6567,N_5586,N_4847);
nor U6568 (N_6568,N_4928,N_5806);
nand U6569 (N_6569,N_5786,N_5176);
and U6570 (N_6570,N_5267,N_5455);
and U6571 (N_6571,N_5935,N_4783);
nor U6572 (N_6572,N_5202,N_5978);
xnor U6573 (N_6573,N_5078,N_5177);
or U6574 (N_6574,N_5194,N_5980);
xnor U6575 (N_6575,N_4843,N_5492);
nand U6576 (N_6576,N_5907,N_5958);
or U6577 (N_6577,N_5147,N_4674);
xor U6578 (N_6578,N_5411,N_4756);
or U6579 (N_6579,N_5315,N_5549);
nor U6580 (N_6580,N_4661,N_5655);
nand U6581 (N_6581,N_5977,N_5913);
xnor U6582 (N_6582,N_4794,N_5535);
or U6583 (N_6583,N_5396,N_5268);
and U6584 (N_6584,N_4623,N_4909);
or U6585 (N_6585,N_5156,N_4532);
xnor U6586 (N_6586,N_5945,N_5067);
or U6587 (N_6587,N_4901,N_5712);
and U6588 (N_6588,N_4807,N_5326);
or U6589 (N_6589,N_5043,N_5105);
xnor U6590 (N_6590,N_4932,N_5121);
and U6591 (N_6591,N_5571,N_5820);
xnor U6592 (N_6592,N_5250,N_5051);
and U6593 (N_6593,N_5303,N_5296);
nor U6594 (N_6594,N_5129,N_4609);
or U6595 (N_6595,N_5972,N_5463);
xor U6596 (N_6596,N_5025,N_5055);
and U6597 (N_6597,N_4877,N_4594);
nand U6598 (N_6598,N_5912,N_4643);
or U6599 (N_6599,N_4723,N_4981);
nor U6600 (N_6600,N_5039,N_5886);
or U6601 (N_6601,N_5953,N_5833);
nand U6602 (N_6602,N_5607,N_5204);
xnor U6603 (N_6603,N_4602,N_5895);
and U6604 (N_6604,N_4596,N_5201);
or U6605 (N_6605,N_4565,N_5985);
nor U6606 (N_6606,N_4857,N_4821);
xnor U6607 (N_6607,N_5859,N_5282);
nor U6608 (N_6608,N_5871,N_5541);
nand U6609 (N_6609,N_4717,N_4531);
nor U6610 (N_6610,N_5314,N_5172);
xor U6611 (N_6611,N_5801,N_5763);
nand U6612 (N_6612,N_5647,N_5971);
nand U6613 (N_6613,N_5812,N_5270);
or U6614 (N_6614,N_4693,N_5169);
or U6615 (N_6615,N_4649,N_5581);
xor U6616 (N_6616,N_4771,N_5398);
nor U6617 (N_6617,N_5188,N_5947);
or U6618 (N_6618,N_5471,N_5995);
or U6619 (N_6619,N_5751,N_4825);
and U6620 (N_6620,N_4900,N_5429);
nand U6621 (N_6621,N_4810,N_5012);
nand U6622 (N_6622,N_5873,N_5370);
nor U6623 (N_6623,N_5391,N_5311);
xor U6624 (N_6624,N_5014,N_5539);
and U6625 (N_6625,N_5883,N_4538);
or U6626 (N_6626,N_5520,N_4801);
nor U6627 (N_6627,N_5837,N_4656);
and U6628 (N_6628,N_5752,N_5330);
nor U6629 (N_6629,N_5781,N_5117);
nand U6630 (N_6630,N_5744,N_4557);
nand U6631 (N_6631,N_4618,N_5679);
or U6632 (N_6632,N_4611,N_4779);
and U6633 (N_6633,N_5144,N_5848);
nor U6634 (N_6634,N_5133,N_5779);
and U6635 (N_6635,N_4567,N_5211);
or U6636 (N_6636,N_5423,N_5558);
and U6637 (N_6637,N_5235,N_5965);
and U6638 (N_6638,N_5901,N_4999);
nor U6639 (N_6639,N_5413,N_4818);
and U6640 (N_6640,N_4564,N_5929);
or U6641 (N_6641,N_5791,N_4512);
nand U6642 (N_6642,N_4989,N_5502);
and U6643 (N_6643,N_5729,N_5973);
xor U6644 (N_6644,N_5163,N_4931);
xnor U6645 (N_6645,N_4836,N_5013);
xor U6646 (N_6646,N_5351,N_5032);
or U6647 (N_6647,N_4998,N_5841);
or U6648 (N_6648,N_5576,N_5274);
nand U6649 (N_6649,N_4852,N_4833);
and U6650 (N_6650,N_5635,N_4521);
nand U6651 (N_6651,N_5150,N_4651);
nor U6652 (N_6652,N_5421,N_5709);
nand U6653 (N_6653,N_5187,N_4912);
or U6654 (N_6654,N_4608,N_5116);
or U6655 (N_6655,N_5555,N_5544);
nor U6656 (N_6656,N_5693,N_4863);
xnor U6657 (N_6657,N_4911,N_5723);
or U6658 (N_6658,N_5595,N_4781);
or U6659 (N_6659,N_4902,N_5142);
and U6660 (N_6660,N_5969,N_5713);
or U6661 (N_6661,N_5161,N_5885);
and U6662 (N_6662,N_5278,N_5674);
or U6663 (N_6663,N_4838,N_5735);
nor U6664 (N_6664,N_5508,N_5612);
nand U6665 (N_6665,N_4633,N_5734);
nor U6666 (N_6666,N_5289,N_5757);
nor U6667 (N_6667,N_4992,N_5342);
nor U6668 (N_6668,N_4961,N_5042);
and U6669 (N_6669,N_5316,N_5991);
or U6670 (N_6670,N_4840,N_4851);
nand U6671 (N_6671,N_5162,N_5020);
and U6672 (N_6672,N_5519,N_4591);
xnor U6673 (N_6673,N_4985,N_4792);
and U6674 (N_6674,N_5425,N_5153);
nor U6675 (N_6675,N_5159,N_4744);
and U6676 (N_6676,N_4724,N_5507);
or U6677 (N_6677,N_4554,N_4871);
nand U6678 (N_6678,N_5731,N_5313);
xnor U6679 (N_6679,N_4716,N_5777);
nor U6680 (N_6680,N_5191,N_5224);
nor U6681 (N_6681,N_4537,N_4841);
or U6682 (N_6682,N_5174,N_4766);
nor U6683 (N_6683,N_5811,N_4906);
and U6684 (N_6684,N_5372,N_5630);
nor U6685 (N_6685,N_5550,N_4549);
or U6686 (N_6686,N_4696,N_5858);
and U6687 (N_6687,N_4940,N_4713);
or U6688 (N_6688,N_5802,N_5138);
nand U6689 (N_6689,N_4694,N_4819);
xnor U6690 (N_6690,N_5386,N_5139);
nor U6691 (N_6691,N_5299,N_4823);
xnor U6692 (N_6692,N_5022,N_4780);
and U6693 (N_6693,N_5240,N_4790);
nand U6694 (N_6694,N_5166,N_5048);
xor U6695 (N_6695,N_4935,N_5428);
and U6696 (N_6696,N_4930,N_5024);
nor U6697 (N_6697,N_5027,N_5642);
or U6698 (N_6698,N_5186,N_5911);
nor U6699 (N_6699,N_4726,N_5089);
xor U6700 (N_6700,N_5040,N_5026);
or U6701 (N_6701,N_5748,N_5101);
nor U6702 (N_6702,N_5591,N_5338);
nor U6703 (N_6703,N_5193,N_5718);
or U6704 (N_6704,N_4933,N_5685);
or U6705 (N_6705,N_5312,N_4947);
xnor U6706 (N_6706,N_5938,N_5281);
xnor U6707 (N_6707,N_5741,N_4835);
nand U6708 (N_6708,N_5730,N_5241);
nand U6709 (N_6709,N_4799,N_5077);
xnor U6710 (N_6710,N_5934,N_5909);
xnor U6711 (N_6711,N_5489,N_5949);
nand U6712 (N_6712,N_4865,N_5475);
or U6713 (N_6713,N_5926,N_5970);
and U6714 (N_6714,N_5285,N_5606);
xor U6715 (N_6715,N_4958,N_4842);
nand U6716 (N_6716,N_5258,N_5828);
and U6717 (N_6717,N_5137,N_5711);
or U6718 (N_6718,N_5412,N_5574);
nor U6719 (N_6719,N_5798,N_4893);
nand U6720 (N_6720,N_5483,N_5810);
xnor U6721 (N_6721,N_4905,N_5357);
nand U6722 (N_6722,N_5106,N_4507);
nor U6723 (N_6723,N_4803,N_5504);
xnor U6724 (N_6724,N_5639,N_4606);
and U6725 (N_6725,N_5940,N_4504);
and U6726 (N_6726,N_4769,N_5835);
nor U6727 (N_6727,N_5094,N_5222);
or U6728 (N_6728,N_4646,N_5721);
and U6729 (N_6729,N_4518,N_5214);
nand U6730 (N_6730,N_5697,N_5488);
or U6731 (N_6731,N_5124,N_5322);
nor U6732 (N_6732,N_5130,N_5339);
xnor U6733 (N_6733,N_4826,N_5720);
xor U6734 (N_6734,N_5125,N_5418);
nand U6735 (N_6735,N_5053,N_4725);
nor U6736 (N_6736,N_4612,N_4683);
nand U6737 (N_6737,N_5490,N_4858);
and U6738 (N_6738,N_5432,N_4814);
nand U6739 (N_6739,N_5902,N_4831);
or U6740 (N_6740,N_4563,N_5919);
xor U6741 (N_6741,N_5795,N_4943);
and U6742 (N_6742,N_4806,N_5081);
or U6743 (N_6743,N_5356,N_4941);
nor U6744 (N_6744,N_5898,N_5208);
nand U6745 (N_6745,N_5839,N_4519);
nor U6746 (N_6746,N_5052,N_5797);
xnor U6747 (N_6747,N_5862,N_5854);
nor U6748 (N_6748,N_4710,N_4503);
and U6749 (N_6749,N_5669,N_5582);
and U6750 (N_6750,N_5376,N_5639);
or U6751 (N_6751,N_5835,N_4861);
or U6752 (N_6752,N_5107,N_5055);
nand U6753 (N_6753,N_5930,N_4693);
or U6754 (N_6754,N_5367,N_5632);
xnor U6755 (N_6755,N_5451,N_5144);
xor U6756 (N_6756,N_5134,N_5617);
nor U6757 (N_6757,N_4748,N_5088);
xnor U6758 (N_6758,N_5354,N_4975);
nand U6759 (N_6759,N_5146,N_4869);
nand U6760 (N_6760,N_5637,N_4953);
or U6761 (N_6761,N_5252,N_4681);
or U6762 (N_6762,N_4799,N_5724);
or U6763 (N_6763,N_4621,N_5894);
or U6764 (N_6764,N_4584,N_5539);
xnor U6765 (N_6765,N_5857,N_4902);
nor U6766 (N_6766,N_4969,N_5406);
xor U6767 (N_6767,N_5841,N_5056);
or U6768 (N_6768,N_5506,N_5988);
nand U6769 (N_6769,N_5812,N_4841);
or U6770 (N_6770,N_5711,N_4915);
nand U6771 (N_6771,N_5792,N_5920);
nand U6772 (N_6772,N_5190,N_5599);
nor U6773 (N_6773,N_5803,N_5263);
nand U6774 (N_6774,N_4677,N_5637);
and U6775 (N_6775,N_5485,N_5234);
and U6776 (N_6776,N_4834,N_5349);
xor U6777 (N_6777,N_5644,N_4777);
or U6778 (N_6778,N_5310,N_5157);
nor U6779 (N_6779,N_5227,N_4542);
xor U6780 (N_6780,N_4761,N_5507);
nand U6781 (N_6781,N_5220,N_4602);
nand U6782 (N_6782,N_4724,N_5790);
nand U6783 (N_6783,N_5377,N_4677);
xor U6784 (N_6784,N_4623,N_4933);
and U6785 (N_6785,N_5967,N_4957);
nand U6786 (N_6786,N_5808,N_4764);
xnor U6787 (N_6787,N_5299,N_5920);
nand U6788 (N_6788,N_4729,N_4777);
or U6789 (N_6789,N_5575,N_4673);
or U6790 (N_6790,N_5790,N_5163);
xor U6791 (N_6791,N_5615,N_5125);
and U6792 (N_6792,N_5092,N_5429);
nor U6793 (N_6793,N_5746,N_5774);
nor U6794 (N_6794,N_5260,N_5570);
nor U6795 (N_6795,N_5684,N_5089);
xor U6796 (N_6796,N_5270,N_5089);
nor U6797 (N_6797,N_5176,N_5304);
nand U6798 (N_6798,N_4761,N_4546);
or U6799 (N_6799,N_5452,N_4915);
and U6800 (N_6800,N_4700,N_5007);
nand U6801 (N_6801,N_5780,N_4902);
and U6802 (N_6802,N_5950,N_5486);
nor U6803 (N_6803,N_5574,N_5180);
and U6804 (N_6804,N_5095,N_4518);
nor U6805 (N_6805,N_4929,N_5608);
nand U6806 (N_6806,N_5379,N_4729);
nand U6807 (N_6807,N_5905,N_5104);
nor U6808 (N_6808,N_5589,N_4710);
nor U6809 (N_6809,N_5134,N_4720);
nor U6810 (N_6810,N_4954,N_5940);
nand U6811 (N_6811,N_4892,N_4755);
nor U6812 (N_6812,N_4909,N_4882);
nor U6813 (N_6813,N_5744,N_5438);
xor U6814 (N_6814,N_4718,N_5458);
nand U6815 (N_6815,N_5386,N_5865);
nor U6816 (N_6816,N_5410,N_5315);
and U6817 (N_6817,N_4606,N_4891);
xnor U6818 (N_6818,N_5148,N_5567);
xor U6819 (N_6819,N_5535,N_5980);
nand U6820 (N_6820,N_5945,N_4730);
or U6821 (N_6821,N_5766,N_4963);
and U6822 (N_6822,N_5128,N_4751);
xor U6823 (N_6823,N_5748,N_4805);
and U6824 (N_6824,N_5618,N_4842);
nor U6825 (N_6825,N_5119,N_5969);
xnor U6826 (N_6826,N_5658,N_5530);
xor U6827 (N_6827,N_5803,N_5974);
nor U6828 (N_6828,N_5115,N_5022);
nand U6829 (N_6829,N_5012,N_5414);
xor U6830 (N_6830,N_4633,N_5075);
xor U6831 (N_6831,N_5278,N_5611);
or U6832 (N_6832,N_5333,N_5954);
xnor U6833 (N_6833,N_4534,N_5613);
or U6834 (N_6834,N_5846,N_5380);
or U6835 (N_6835,N_5719,N_5522);
nor U6836 (N_6836,N_5446,N_4827);
nor U6837 (N_6837,N_4932,N_5076);
or U6838 (N_6838,N_4588,N_5462);
or U6839 (N_6839,N_4528,N_5001);
or U6840 (N_6840,N_5237,N_5594);
xor U6841 (N_6841,N_4773,N_5443);
nand U6842 (N_6842,N_4522,N_5228);
nand U6843 (N_6843,N_4990,N_5906);
and U6844 (N_6844,N_4836,N_4907);
nor U6845 (N_6845,N_5567,N_5244);
or U6846 (N_6846,N_4654,N_5251);
nand U6847 (N_6847,N_5112,N_5629);
nor U6848 (N_6848,N_4710,N_5746);
xnor U6849 (N_6849,N_5251,N_5337);
and U6850 (N_6850,N_5661,N_5307);
or U6851 (N_6851,N_4631,N_5731);
and U6852 (N_6852,N_5173,N_5448);
or U6853 (N_6853,N_5727,N_5392);
nand U6854 (N_6854,N_5006,N_4823);
nand U6855 (N_6855,N_5630,N_5276);
and U6856 (N_6856,N_5273,N_5299);
xor U6857 (N_6857,N_4955,N_5398);
xnor U6858 (N_6858,N_5731,N_4827);
or U6859 (N_6859,N_5755,N_4929);
nor U6860 (N_6860,N_4827,N_5770);
or U6861 (N_6861,N_5822,N_5989);
nand U6862 (N_6862,N_4872,N_4811);
and U6863 (N_6863,N_4748,N_4743);
or U6864 (N_6864,N_5190,N_4582);
nand U6865 (N_6865,N_5060,N_5019);
xor U6866 (N_6866,N_5797,N_5408);
nand U6867 (N_6867,N_5489,N_5899);
nand U6868 (N_6868,N_4690,N_5178);
xor U6869 (N_6869,N_4824,N_4859);
and U6870 (N_6870,N_5197,N_4844);
and U6871 (N_6871,N_5110,N_5610);
and U6872 (N_6872,N_5911,N_4896);
xor U6873 (N_6873,N_5999,N_5725);
xnor U6874 (N_6874,N_4857,N_5436);
nor U6875 (N_6875,N_5593,N_4686);
nor U6876 (N_6876,N_5908,N_4971);
or U6877 (N_6877,N_5097,N_5619);
nor U6878 (N_6878,N_5249,N_4807);
nor U6879 (N_6879,N_5106,N_5041);
nand U6880 (N_6880,N_5263,N_5412);
xnor U6881 (N_6881,N_5158,N_5421);
or U6882 (N_6882,N_4940,N_5363);
nand U6883 (N_6883,N_4569,N_4999);
xor U6884 (N_6884,N_4785,N_4529);
xnor U6885 (N_6885,N_5889,N_5761);
or U6886 (N_6886,N_4595,N_4538);
nor U6887 (N_6887,N_5324,N_5556);
nand U6888 (N_6888,N_5585,N_5569);
or U6889 (N_6889,N_5917,N_5214);
nand U6890 (N_6890,N_5511,N_5698);
nor U6891 (N_6891,N_4942,N_4940);
nand U6892 (N_6892,N_4587,N_4679);
and U6893 (N_6893,N_4919,N_5256);
nand U6894 (N_6894,N_4655,N_5282);
or U6895 (N_6895,N_5630,N_5318);
or U6896 (N_6896,N_4725,N_5019);
nand U6897 (N_6897,N_5548,N_5509);
and U6898 (N_6898,N_5400,N_5126);
or U6899 (N_6899,N_4666,N_5815);
or U6900 (N_6900,N_5038,N_5831);
or U6901 (N_6901,N_5537,N_5531);
xor U6902 (N_6902,N_5809,N_5007);
or U6903 (N_6903,N_5960,N_5583);
nand U6904 (N_6904,N_5989,N_5913);
and U6905 (N_6905,N_5316,N_5404);
or U6906 (N_6906,N_5305,N_5203);
or U6907 (N_6907,N_5620,N_4689);
nand U6908 (N_6908,N_5035,N_5899);
nor U6909 (N_6909,N_5801,N_5447);
or U6910 (N_6910,N_5670,N_5330);
xnor U6911 (N_6911,N_5100,N_4786);
and U6912 (N_6912,N_5332,N_4858);
or U6913 (N_6913,N_5177,N_5366);
and U6914 (N_6914,N_5169,N_4660);
or U6915 (N_6915,N_4622,N_4595);
nand U6916 (N_6916,N_5846,N_4840);
xor U6917 (N_6917,N_4570,N_5483);
and U6918 (N_6918,N_5882,N_5614);
or U6919 (N_6919,N_4536,N_5221);
nand U6920 (N_6920,N_4849,N_5039);
or U6921 (N_6921,N_5444,N_4985);
xor U6922 (N_6922,N_5143,N_4930);
nand U6923 (N_6923,N_4783,N_5363);
and U6924 (N_6924,N_4886,N_5830);
xor U6925 (N_6925,N_4727,N_4564);
xor U6926 (N_6926,N_5451,N_4560);
xor U6927 (N_6927,N_5518,N_5930);
nand U6928 (N_6928,N_5434,N_4550);
nand U6929 (N_6929,N_4593,N_5274);
or U6930 (N_6930,N_4861,N_4926);
xnor U6931 (N_6931,N_4784,N_5404);
or U6932 (N_6932,N_5922,N_5665);
and U6933 (N_6933,N_5085,N_5161);
xnor U6934 (N_6934,N_4528,N_5432);
or U6935 (N_6935,N_5652,N_4941);
and U6936 (N_6936,N_4955,N_5315);
nand U6937 (N_6937,N_5120,N_4924);
nand U6938 (N_6938,N_5794,N_5182);
and U6939 (N_6939,N_5911,N_5480);
xnor U6940 (N_6940,N_5246,N_5952);
nand U6941 (N_6941,N_4843,N_4522);
nand U6942 (N_6942,N_5242,N_4867);
or U6943 (N_6943,N_4536,N_5528);
xnor U6944 (N_6944,N_5323,N_5574);
xor U6945 (N_6945,N_4609,N_4936);
xor U6946 (N_6946,N_5356,N_4914);
and U6947 (N_6947,N_5483,N_4659);
xor U6948 (N_6948,N_5070,N_5780);
and U6949 (N_6949,N_4962,N_5944);
xor U6950 (N_6950,N_5647,N_5928);
and U6951 (N_6951,N_5981,N_5614);
and U6952 (N_6952,N_4684,N_5686);
or U6953 (N_6953,N_4878,N_5655);
xnor U6954 (N_6954,N_4658,N_5045);
and U6955 (N_6955,N_5614,N_5373);
nor U6956 (N_6956,N_5613,N_5998);
and U6957 (N_6957,N_5294,N_5217);
xor U6958 (N_6958,N_4726,N_4637);
and U6959 (N_6959,N_5877,N_5762);
and U6960 (N_6960,N_5279,N_5209);
or U6961 (N_6961,N_4985,N_5408);
and U6962 (N_6962,N_5878,N_5788);
or U6963 (N_6963,N_4501,N_4790);
nand U6964 (N_6964,N_5203,N_4538);
and U6965 (N_6965,N_5229,N_4986);
and U6966 (N_6966,N_4822,N_5484);
nor U6967 (N_6967,N_5798,N_5543);
and U6968 (N_6968,N_5653,N_5586);
nor U6969 (N_6969,N_5118,N_5149);
or U6970 (N_6970,N_5984,N_5589);
and U6971 (N_6971,N_4927,N_4506);
nor U6972 (N_6972,N_4689,N_4820);
nand U6973 (N_6973,N_5903,N_5975);
xor U6974 (N_6974,N_5280,N_4977);
nor U6975 (N_6975,N_4791,N_4649);
nor U6976 (N_6976,N_5262,N_5369);
and U6977 (N_6977,N_4787,N_4798);
nand U6978 (N_6978,N_4888,N_4628);
xor U6979 (N_6979,N_5054,N_5237);
xnor U6980 (N_6980,N_4501,N_5354);
xnor U6981 (N_6981,N_4716,N_5076);
xor U6982 (N_6982,N_4574,N_4991);
xor U6983 (N_6983,N_4990,N_5990);
nand U6984 (N_6984,N_5451,N_5826);
nor U6985 (N_6985,N_5854,N_5447);
nand U6986 (N_6986,N_4751,N_5460);
or U6987 (N_6987,N_4586,N_4867);
or U6988 (N_6988,N_5621,N_5861);
nor U6989 (N_6989,N_4716,N_5448);
xor U6990 (N_6990,N_4732,N_5511);
nor U6991 (N_6991,N_5105,N_5197);
and U6992 (N_6992,N_4516,N_4606);
and U6993 (N_6993,N_4559,N_4678);
and U6994 (N_6994,N_5423,N_4605);
or U6995 (N_6995,N_4923,N_4751);
and U6996 (N_6996,N_4508,N_4932);
xnor U6997 (N_6997,N_4767,N_4542);
xor U6998 (N_6998,N_5752,N_4872);
nand U6999 (N_6999,N_4944,N_5951);
and U7000 (N_7000,N_5258,N_5304);
xor U7001 (N_7001,N_4558,N_5968);
or U7002 (N_7002,N_5037,N_5855);
xor U7003 (N_7003,N_4735,N_5147);
or U7004 (N_7004,N_5644,N_5138);
nand U7005 (N_7005,N_4586,N_5606);
or U7006 (N_7006,N_5784,N_4518);
nor U7007 (N_7007,N_5905,N_5683);
xnor U7008 (N_7008,N_5407,N_5735);
nor U7009 (N_7009,N_5510,N_5049);
xnor U7010 (N_7010,N_5681,N_5476);
and U7011 (N_7011,N_5079,N_4735);
and U7012 (N_7012,N_4744,N_5905);
nand U7013 (N_7013,N_5796,N_5346);
nor U7014 (N_7014,N_5760,N_5276);
and U7015 (N_7015,N_5413,N_4747);
xor U7016 (N_7016,N_4817,N_5539);
and U7017 (N_7017,N_4609,N_5013);
nor U7018 (N_7018,N_4750,N_4825);
and U7019 (N_7019,N_4698,N_5655);
xnor U7020 (N_7020,N_5414,N_5972);
and U7021 (N_7021,N_4987,N_5311);
or U7022 (N_7022,N_5635,N_5898);
nand U7023 (N_7023,N_4836,N_5405);
nor U7024 (N_7024,N_4641,N_4515);
and U7025 (N_7025,N_5463,N_5208);
nand U7026 (N_7026,N_4559,N_5506);
nor U7027 (N_7027,N_5760,N_5991);
or U7028 (N_7028,N_5458,N_5323);
and U7029 (N_7029,N_4666,N_5103);
or U7030 (N_7030,N_5229,N_5874);
nand U7031 (N_7031,N_5850,N_5439);
or U7032 (N_7032,N_5720,N_5031);
or U7033 (N_7033,N_4934,N_4888);
nand U7034 (N_7034,N_4886,N_5966);
or U7035 (N_7035,N_5326,N_5418);
nand U7036 (N_7036,N_5688,N_4932);
and U7037 (N_7037,N_5276,N_4886);
nand U7038 (N_7038,N_5221,N_4990);
and U7039 (N_7039,N_5593,N_5620);
or U7040 (N_7040,N_4781,N_4773);
or U7041 (N_7041,N_5455,N_5580);
nor U7042 (N_7042,N_4742,N_5659);
nand U7043 (N_7043,N_5792,N_5358);
nand U7044 (N_7044,N_5461,N_5931);
nand U7045 (N_7045,N_4732,N_5761);
or U7046 (N_7046,N_5493,N_4573);
xnor U7047 (N_7047,N_5279,N_4602);
and U7048 (N_7048,N_4576,N_4644);
or U7049 (N_7049,N_5971,N_5022);
nor U7050 (N_7050,N_4521,N_4671);
or U7051 (N_7051,N_5708,N_5858);
or U7052 (N_7052,N_4711,N_5902);
and U7053 (N_7053,N_4674,N_5504);
nand U7054 (N_7054,N_5114,N_5746);
or U7055 (N_7055,N_5418,N_4715);
nor U7056 (N_7056,N_4783,N_5095);
or U7057 (N_7057,N_5633,N_5689);
nor U7058 (N_7058,N_4506,N_5170);
xor U7059 (N_7059,N_5847,N_5434);
or U7060 (N_7060,N_5168,N_5693);
xnor U7061 (N_7061,N_5084,N_5141);
xor U7062 (N_7062,N_5567,N_4657);
nand U7063 (N_7063,N_5065,N_5900);
nand U7064 (N_7064,N_4768,N_5160);
xnor U7065 (N_7065,N_4649,N_5832);
xor U7066 (N_7066,N_4783,N_4546);
nand U7067 (N_7067,N_5273,N_5628);
nor U7068 (N_7068,N_5714,N_5864);
nor U7069 (N_7069,N_5458,N_4712);
xor U7070 (N_7070,N_4950,N_5158);
xor U7071 (N_7071,N_4719,N_5131);
xnor U7072 (N_7072,N_5181,N_4858);
nand U7073 (N_7073,N_4502,N_5840);
or U7074 (N_7074,N_5574,N_5668);
nand U7075 (N_7075,N_4615,N_4733);
xnor U7076 (N_7076,N_5560,N_5524);
nor U7077 (N_7077,N_5139,N_5032);
or U7078 (N_7078,N_4786,N_5488);
xor U7079 (N_7079,N_4928,N_5876);
and U7080 (N_7080,N_5205,N_4885);
or U7081 (N_7081,N_4813,N_5178);
xnor U7082 (N_7082,N_4552,N_5592);
xnor U7083 (N_7083,N_4594,N_4977);
nor U7084 (N_7084,N_5140,N_5567);
or U7085 (N_7085,N_4808,N_4818);
and U7086 (N_7086,N_5031,N_4786);
nor U7087 (N_7087,N_5613,N_5444);
nor U7088 (N_7088,N_5926,N_5933);
xor U7089 (N_7089,N_5222,N_5343);
nand U7090 (N_7090,N_4617,N_5701);
or U7091 (N_7091,N_5256,N_5125);
nand U7092 (N_7092,N_4685,N_5525);
nor U7093 (N_7093,N_5154,N_4626);
nand U7094 (N_7094,N_4588,N_4921);
xnor U7095 (N_7095,N_4965,N_5112);
nand U7096 (N_7096,N_5318,N_4671);
nand U7097 (N_7097,N_4512,N_4964);
nor U7098 (N_7098,N_5443,N_5829);
and U7099 (N_7099,N_5972,N_5214);
and U7100 (N_7100,N_5132,N_5784);
or U7101 (N_7101,N_4904,N_5599);
or U7102 (N_7102,N_5323,N_5910);
nand U7103 (N_7103,N_4940,N_5107);
nand U7104 (N_7104,N_4591,N_5011);
xnor U7105 (N_7105,N_5350,N_5742);
xor U7106 (N_7106,N_5684,N_5357);
or U7107 (N_7107,N_5352,N_4669);
and U7108 (N_7108,N_5765,N_5337);
xor U7109 (N_7109,N_5794,N_4677);
nand U7110 (N_7110,N_4720,N_4788);
xor U7111 (N_7111,N_5248,N_5715);
xnor U7112 (N_7112,N_5753,N_5217);
nor U7113 (N_7113,N_4772,N_4885);
and U7114 (N_7114,N_4600,N_4823);
nor U7115 (N_7115,N_5193,N_5930);
nand U7116 (N_7116,N_5215,N_4645);
and U7117 (N_7117,N_5791,N_5633);
nand U7118 (N_7118,N_4951,N_5247);
nand U7119 (N_7119,N_5910,N_5321);
xnor U7120 (N_7120,N_5437,N_5934);
or U7121 (N_7121,N_4899,N_4900);
nand U7122 (N_7122,N_5851,N_4700);
or U7123 (N_7123,N_5803,N_5960);
xnor U7124 (N_7124,N_4543,N_4867);
nand U7125 (N_7125,N_4563,N_4841);
nor U7126 (N_7126,N_4686,N_4540);
nand U7127 (N_7127,N_4584,N_5595);
nand U7128 (N_7128,N_5884,N_5203);
xor U7129 (N_7129,N_5453,N_5160);
or U7130 (N_7130,N_4988,N_5308);
nand U7131 (N_7131,N_4587,N_5615);
nand U7132 (N_7132,N_5022,N_5271);
xor U7133 (N_7133,N_4597,N_5840);
nand U7134 (N_7134,N_4920,N_5437);
xor U7135 (N_7135,N_5514,N_5304);
xnor U7136 (N_7136,N_5412,N_5907);
xor U7137 (N_7137,N_5234,N_4984);
xor U7138 (N_7138,N_5075,N_5787);
or U7139 (N_7139,N_5608,N_5531);
nor U7140 (N_7140,N_5199,N_5999);
xnor U7141 (N_7141,N_5721,N_4852);
or U7142 (N_7142,N_5492,N_5408);
or U7143 (N_7143,N_4589,N_4684);
or U7144 (N_7144,N_5305,N_5984);
and U7145 (N_7145,N_5424,N_5103);
nand U7146 (N_7146,N_5383,N_5052);
nor U7147 (N_7147,N_4685,N_5761);
nand U7148 (N_7148,N_5375,N_5893);
xor U7149 (N_7149,N_5558,N_5802);
nor U7150 (N_7150,N_5675,N_5870);
xnor U7151 (N_7151,N_4680,N_4778);
xnor U7152 (N_7152,N_4972,N_4605);
nor U7153 (N_7153,N_5738,N_4542);
and U7154 (N_7154,N_4987,N_4629);
and U7155 (N_7155,N_4965,N_5368);
nor U7156 (N_7156,N_5251,N_4689);
nor U7157 (N_7157,N_5647,N_5358);
xor U7158 (N_7158,N_5653,N_5595);
and U7159 (N_7159,N_5694,N_4642);
xor U7160 (N_7160,N_4611,N_5126);
and U7161 (N_7161,N_5119,N_4804);
and U7162 (N_7162,N_4973,N_5961);
and U7163 (N_7163,N_5109,N_4910);
nor U7164 (N_7164,N_5047,N_5578);
nand U7165 (N_7165,N_5430,N_4821);
nand U7166 (N_7166,N_5209,N_5481);
nand U7167 (N_7167,N_5375,N_5409);
nor U7168 (N_7168,N_5961,N_5112);
xnor U7169 (N_7169,N_5543,N_5623);
and U7170 (N_7170,N_5730,N_5877);
xnor U7171 (N_7171,N_4808,N_5446);
nand U7172 (N_7172,N_5972,N_5879);
nor U7173 (N_7173,N_5475,N_5023);
nor U7174 (N_7174,N_5025,N_4861);
nor U7175 (N_7175,N_5477,N_5315);
xor U7176 (N_7176,N_5888,N_5557);
xor U7177 (N_7177,N_5852,N_5133);
nor U7178 (N_7178,N_5338,N_5792);
nor U7179 (N_7179,N_5976,N_4703);
nor U7180 (N_7180,N_5153,N_5737);
nand U7181 (N_7181,N_4991,N_5677);
or U7182 (N_7182,N_5748,N_5369);
or U7183 (N_7183,N_5065,N_4824);
nor U7184 (N_7184,N_5044,N_5767);
nor U7185 (N_7185,N_4877,N_4609);
xnor U7186 (N_7186,N_5908,N_4852);
xor U7187 (N_7187,N_4709,N_4721);
and U7188 (N_7188,N_5995,N_5720);
nor U7189 (N_7189,N_5122,N_5950);
nand U7190 (N_7190,N_4858,N_4744);
nor U7191 (N_7191,N_5929,N_5585);
nand U7192 (N_7192,N_5587,N_5170);
xnor U7193 (N_7193,N_5260,N_5947);
nor U7194 (N_7194,N_4610,N_5210);
xnor U7195 (N_7195,N_4826,N_5792);
xor U7196 (N_7196,N_5622,N_5791);
xor U7197 (N_7197,N_4663,N_5986);
nand U7198 (N_7198,N_5945,N_5432);
or U7199 (N_7199,N_5922,N_4669);
nor U7200 (N_7200,N_5836,N_5780);
and U7201 (N_7201,N_4707,N_5086);
and U7202 (N_7202,N_5812,N_4926);
nor U7203 (N_7203,N_5173,N_4968);
nor U7204 (N_7204,N_4804,N_5469);
or U7205 (N_7205,N_5992,N_4669);
nor U7206 (N_7206,N_5091,N_4746);
and U7207 (N_7207,N_5120,N_4646);
nor U7208 (N_7208,N_5200,N_5271);
xnor U7209 (N_7209,N_5320,N_5948);
or U7210 (N_7210,N_4774,N_5241);
xor U7211 (N_7211,N_5684,N_5572);
and U7212 (N_7212,N_5028,N_5112);
nor U7213 (N_7213,N_4829,N_5001);
nor U7214 (N_7214,N_5149,N_5307);
nor U7215 (N_7215,N_5499,N_5407);
xnor U7216 (N_7216,N_4655,N_5474);
or U7217 (N_7217,N_5111,N_4538);
nor U7218 (N_7218,N_4618,N_4811);
or U7219 (N_7219,N_4727,N_5107);
or U7220 (N_7220,N_4969,N_5804);
xor U7221 (N_7221,N_5085,N_5889);
xnor U7222 (N_7222,N_5727,N_5735);
or U7223 (N_7223,N_5290,N_5106);
or U7224 (N_7224,N_5801,N_4665);
and U7225 (N_7225,N_5513,N_4510);
xnor U7226 (N_7226,N_4760,N_5718);
xor U7227 (N_7227,N_5415,N_5460);
and U7228 (N_7228,N_4868,N_5910);
and U7229 (N_7229,N_5550,N_4967);
xnor U7230 (N_7230,N_5863,N_5742);
or U7231 (N_7231,N_5524,N_4596);
nand U7232 (N_7232,N_4546,N_5421);
or U7233 (N_7233,N_4531,N_5196);
nor U7234 (N_7234,N_4770,N_4641);
xnor U7235 (N_7235,N_4973,N_5455);
xor U7236 (N_7236,N_5253,N_4576);
xnor U7237 (N_7237,N_5293,N_4592);
nor U7238 (N_7238,N_4716,N_4891);
xor U7239 (N_7239,N_5311,N_5239);
and U7240 (N_7240,N_5220,N_5819);
xnor U7241 (N_7241,N_4949,N_5525);
or U7242 (N_7242,N_5194,N_4519);
xnor U7243 (N_7243,N_4929,N_5430);
or U7244 (N_7244,N_4576,N_5791);
nand U7245 (N_7245,N_5370,N_5605);
nor U7246 (N_7246,N_4523,N_4501);
nor U7247 (N_7247,N_5566,N_5552);
or U7248 (N_7248,N_5688,N_4520);
nor U7249 (N_7249,N_5838,N_4999);
or U7250 (N_7250,N_5841,N_4714);
nand U7251 (N_7251,N_5483,N_4660);
nor U7252 (N_7252,N_5997,N_5827);
xor U7253 (N_7253,N_5000,N_5331);
xor U7254 (N_7254,N_4983,N_4965);
xnor U7255 (N_7255,N_5984,N_5258);
nor U7256 (N_7256,N_4721,N_4845);
nor U7257 (N_7257,N_5361,N_4630);
or U7258 (N_7258,N_5026,N_5551);
nor U7259 (N_7259,N_5186,N_4662);
xor U7260 (N_7260,N_5855,N_5910);
nor U7261 (N_7261,N_5890,N_5995);
nor U7262 (N_7262,N_5151,N_5808);
or U7263 (N_7263,N_5566,N_5785);
or U7264 (N_7264,N_5962,N_5841);
nor U7265 (N_7265,N_4587,N_5514);
nand U7266 (N_7266,N_4980,N_5762);
nand U7267 (N_7267,N_5991,N_5703);
nand U7268 (N_7268,N_5610,N_4625);
nor U7269 (N_7269,N_5181,N_4537);
nor U7270 (N_7270,N_5429,N_4615);
and U7271 (N_7271,N_4508,N_5272);
or U7272 (N_7272,N_4551,N_4667);
and U7273 (N_7273,N_5973,N_4914);
nor U7274 (N_7274,N_5379,N_5690);
nor U7275 (N_7275,N_5535,N_5742);
nor U7276 (N_7276,N_5324,N_5256);
nor U7277 (N_7277,N_4751,N_5891);
nand U7278 (N_7278,N_5321,N_4537);
xor U7279 (N_7279,N_4917,N_5452);
nand U7280 (N_7280,N_5331,N_5657);
nor U7281 (N_7281,N_5563,N_4739);
xnor U7282 (N_7282,N_5308,N_5802);
and U7283 (N_7283,N_5906,N_5741);
and U7284 (N_7284,N_5358,N_4737);
nor U7285 (N_7285,N_4986,N_4701);
or U7286 (N_7286,N_4921,N_5004);
and U7287 (N_7287,N_4876,N_5056);
nor U7288 (N_7288,N_5404,N_5216);
xor U7289 (N_7289,N_5619,N_5014);
nor U7290 (N_7290,N_5085,N_5104);
xnor U7291 (N_7291,N_5782,N_5188);
or U7292 (N_7292,N_4924,N_5008);
or U7293 (N_7293,N_5926,N_5297);
nand U7294 (N_7294,N_5460,N_5393);
xnor U7295 (N_7295,N_5391,N_5965);
xnor U7296 (N_7296,N_5634,N_4710);
and U7297 (N_7297,N_5194,N_5505);
and U7298 (N_7298,N_5012,N_5604);
nand U7299 (N_7299,N_5660,N_5893);
xnor U7300 (N_7300,N_5692,N_5883);
nor U7301 (N_7301,N_5889,N_4973);
or U7302 (N_7302,N_4681,N_4915);
nand U7303 (N_7303,N_5398,N_5624);
and U7304 (N_7304,N_5421,N_4595);
xnor U7305 (N_7305,N_5882,N_5699);
nor U7306 (N_7306,N_4780,N_5110);
and U7307 (N_7307,N_5988,N_5162);
nor U7308 (N_7308,N_4525,N_5032);
nor U7309 (N_7309,N_4615,N_4875);
or U7310 (N_7310,N_5909,N_5273);
and U7311 (N_7311,N_4593,N_5786);
nand U7312 (N_7312,N_5493,N_5799);
and U7313 (N_7313,N_4732,N_5089);
or U7314 (N_7314,N_4809,N_5565);
nor U7315 (N_7315,N_5335,N_5060);
or U7316 (N_7316,N_4507,N_5132);
xor U7317 (N_7317,N_5202,N_5275);
nand U7318 (N_7318,N_5294,N_4517);
and U7319 (N_7319,N_5446,N_4753);
and U7320 (N_7320,N_4769,N_4817);
nand U7321 (N_7321,N_5748,N_4983);
xnor U7322 (N_7322,N_5484,N_5375);
and U7323 (N_7323,N_5789,N_5821);
nand U7324 (N_7324,N_5624,N_4693);
xor U7325 (N_7325,N_5213,N_5569);
nand U7326 (N_7326,N_5156,N_5119);
or U7327 (N_7327,N_4600,N_5034);
nand U7328 (N_7328,N_5017,N_4755);
nand U7329 (N_7329,N_5025,N_4720);
xnor U7330 (N_7330,N_5755,N_4547);
or U7331 (N_7331,N_4621,N_5405);
or U7332 (N_7332,N_5094,N_4564);
or U7333 (N_7333,N_5032,N_5996);
nor U7334 (N_7334,N_5687,N_5432);
nand U7335 (N_7335,N_5661,N_5679);
or U7336 (N_7336,N_5318,N_5597);
nand U7337 (N_7337,N_4993,N_5472);
and U7338 (N_7338,N_4994,N_5972);
nor U7339 (N_7339,N_4869,N_5425);
nand U7340 (N_7340,N_5016,N_4710);
nor U7341 (N_7341,N_4778,N_5035);
and U7342 (N_7342,N_5417,N_5686);
or U7343 (N_7343,N_4642,N_4991);
nor U7344 (N_7344,N_4666,N_5015);
or U7345 (N_7345,N_5126,N_4693);
nor U7346 (N_7346,N_5237,N_5538);
xor U7347 (N_7347,N_5050,N_5064);
and U7348 (N_7348,N_5308,N_5255);
or U7349 (N_7349,N_4851,N_5820);
and U7350 (N_7350,N_4505,N_5914);
and U7351 (N_7351,N_5452,N_4954);
nor U7352 (N_7352,N_4892,N_5335);
xor U7353 (N_7353,N_5912,N_4910);
and U7354 (N_7354,N_5932,N_5843);
and U7355 (N_7355,N_5675,N_5093);
and U7356 (N_7356,N_4930,N_5994);
or U7357 (N_7357,N_5606,N_5755);
or U7358 (N_7358,N_5270,N_5447);
and U7359 (N_7359,N_5322,N_5877);
xnor U7360 (N_7360,N_5107,N_5095);
or U7361 (N_7361,N_5170,N_5407);
nor U7362 (N_7362,N_4631,N_4890);
xor U7363 (N_7363,N_4586,N_4680);
and U7364 (N_7364,N_5202,N_5519);
nor U7365 (N_7365,N_5707,N_5153);
nor U7366 (N_7366,N_5957,N_5656);
nand U7367 (N_7367,N_5078,N_4901);
nand U7368 (N_7368,N_4950,N_5116);
xnor U7369 (N_7369,N_5201,N_4607);
and U7370 (N_7370,N_5130,N_5939);
nand U7371 (N_7371,N_5897,N_4568);
and U7372 (N_7372,N_5651,N_5180);
xnor U7373 (N_7373,N_5280,N_5071);
nor U7374 (N_7374,N_5998,N_5318);
xor U7375 (N_7375,N_4526,N_4906);
or U7376 (N_7376,N_5709,N_4982);
nor U7377 (N_7377,N_5927,N_5123);
or U7378 (N_7378,N_5478,N_5924);
nor U7379 (N_7379,N_5541,N_5659);
xnor U7380 (N_7380,N_4673,N_5820);
nor U7381 (N_7381,N_5654,N_4989);
or U7382 (N_7382,N_4514,N_5293);
and U7383 (N_7383,N_5215,N_5791);
and U7384 (N_7384,N_4985,N_5778);
and U7385 (N_7385,N_4784,N_4654);
or U7386 (N_7386,N_4858,N_5379);
and U7387 (N_7387,N_5750,N_5993);
nand U7388 (N_7388,N_4757,N_5797);
nor U7389 (N_7389,N_4887,N_4506);
nand U7390 (N_7390,N_4529,N_4660);
nor U7391 (N_7391,N_4529,N_5118);
or U7392 (N_7392,N_5958,N_5579);
and U7393 (N_7393,N_5598,N_5337);
or U7394 (N_7394,N_5751,N_5904);
and U7395 (N_7395,N_4550,N_4586);
and U7396 (N_7396,N_5229,N_5838);
and U7397 (N_7397,N_5305,N_5898);
or U7398 (N_7398,N_5217,N_5454);
xnor U7399 (N_7399,N_4903,N_5983);
or U7400 (N_7400,N_5543,N_4621);
nand U7401 (N_7401,N_4786,N_5905);
nand U7402 (N_7402,N_4614,N_4979);
nor U7403 (N_7403,N_4759,N_5062);
and U7404 (N_7404,N_5121,N_5055);
xor U7405 (N_7405,N_5310,N_5170);
xor U7406 (N_7406,N_4872,N_4635);
xnor U7407 (N_7407,N_5587,N_5626);
and U7408 (N_7408,N_5705,N_5912);
nor U7409 (N_7409,N_4566,N_4934);
xor U7410 (N_7410,N_5526,N_5076);
nor U7411 (N_7411,N_4957,N_4656);
and U7412 (N_7412,N_5123,N_5365);
nor U7413 (N_7413,N_5651,N_5781);
and U7414 (N_7414,N_5221,N_4611);
or U7415 (N_7415,N_5571,N_5602);
nand U7416 (N_7416,N_5481,N_5726);
nor U7417 (N_7417,N_5159,N_4828);
and U7418 (N_7418,N_5852,N_4640);
and U7419 (N_7419,N_5801,N_5287);
nand U7420 (N_7420,N_5477,N_5139);
and U7421 (N_7421,N_5592,N_5593);
and U7422 (N_7422,N_4806,N_5631);
nor U7423 (N_7423,N_4744,N_4910);
xnor U7424 (N_7424,N_5397,N_5065);
nand U7425 (N_7425,N_5130,N_5798);
or U7426 (N_7426,N_4698,N_5848);
nand U7427 (N_7427,N_5657,N_5520);
or U7428 (N_7428,N_5024,N_5913);
and U7429 (N_7429,N_5112,N_5818);
xor U7430 (N_7430,N_5350,N_5463);
or U7431 (N_7431,N_5578,N_4560);
xnor U7432 (N_7432,N_5672,N_4959);
nand U7433 (N_7433,N_4580,N_5978);
nand U7434 (N_7434,N_4619,N_5297);
nor U7435 (N_7435,N_5255,N_4717);
nand U7436 (N_7436,N_5454,N_5408);
nand U7437 (N_7437,N_4935,N_5415);
nor U7438 (N_7438,N_5162,N_4563);
nand U7439 (N_7439,N_5792,N_5055);
or U7440 (N_7440,N_5612,N_4662);
or U7441 (N_7441,N_4512,N_5886);
nor U7442 (N_7442,N_5679,N_4917);
xor U7443 (N_7443,N_4652,N_5575);
nand U7444 (N_7444,N_5045,N_5584);
and U7445 (N_7445,N_4941,N_5475);
nand U7446 (N_7446,N_5245,N_5230);
nand U7447 (N_7447,N_5570,N_5978);
and U7448 (N_7448,N_5961,N_5104);
xor U7449 (N_7449,N_4921,N_5315);
or U7450 (N_7450,N_5491,N_5715);
and U7451 (N_7451,N_4595,N_4926);
nor U7452 (N_7452,N_5397,N_4539);
or U7453 (N_7453,N_4718,N_5186);
nand U7454 (N_7454,N_5307,N_5300);
xnor U7455 (N_7455,N_4680,N_5059);
nand U7456 (N_7456,N_5545,N_4558);
nor U7457 (N_7457,N_5639,N_5948);
xor U7458 (N_7458,N_5674,N_5991);
or U7459 (N_7459,N_5396,N_5591);
and U7460 (N_7460,N_5911,N_4902);
xor U7461 (N_7461,N_5252,N_5435);
or U7462 (N_7462,N_5254,N_5190);
xor U7463 (N_7463,N_4728,N_5434);
and U7464 (N_7464,N_5250,N_4563);
nand U7465 (N_7465,N_4555,N_5113);
xor U7466 (N_7466,N_5882,N_5459);
nand U7467 (N_7467,N_5630,N_4981);
nand U7468 (N_7468,N_4822,N_5998);
or U7469 (N_7469,N_5948,N_5555);
or U7470 (N_7470,N_5282,N_4919);
xor U7471 (N_7471,N_4726,N_5000);
xor U7472 (N_7472,N_5518,N_5902);
nand U7473 (N_7473,N_5500,N_5186);
nand U7474 (N_7474,N_5765,N_5889);
xnor U7475 (N_7475,N_4510,N_4502);
xnor U7476 (N_7476,N_4741,N_4718);
xor U7477 (N_7477,N_5260,N_5246);
and U7478 (N_7478,N_5471,N_5433);
and U7479 (N_7479,N_5241,N_4886);
xnor U7480 (N_7480,N_5086,N_4729);
or U7481 (N_7481,N_4804,N_5354);
or U7482 (N_7482,N_5254,N_5841);
nand U7483 (N_7483,N_4850,N_5671);
and U7484 (N_7484,N_5567,N_5357);
nor U7485 (N_7485,N_5175,N_5393);
xor U7486 (N_7486,N_4520,N_4819);
xnor U7487 (N_7487,N_5328,N_5951);
nand U7488 (N_7488,N_5382,N_5632);
xor U7489 (N_7489,N_5230,N_5946);
and U7490 (N_7490,N_5823,N_5293);
nand U7491 (N_7491,N_5141,N_4796);
xnor U7492 (N_7492,N_5568,N_5170);
nand U7493 (N_7493,N_5849,N_4948);
xnor U7494 (N_7494,N_5041,N_5208);
xnor U7495 (N_7495,N_5794,N_5286);
nand U7496 (N_7496,N_4717,N_5747);
nor U7497 (N_7497,N_5615,N_4594);
and U7498 (N_7498,N_5567,N_5740);
or U7499 (N_7499,N_5125,N_4850);
nor U7500 (N_7500,N_6759,N_6625);
or U7501 (N_7501,N_6844,N_7019);
and U7502 (N_7502,N_6539,N_6374);
nor U7503 (N_7503,N_6371,N_6086);
or U7504 (N_7504,N_7236,N_6803);
nand U7505 (N_7505,N_6834,N_7397);
and U7506 (N_7506,N_6973,N_6248);
xnor U7507 (N_7507,N_6115,N_7297);
and U7508 (N_7508,N_7263,N_6001);
nor U7509 (N_7509,N_7152,N_7206);
and U7510 (N_7510,N_7150,N_7340);
xor U7511 (N_7511,N_6024,N_6111);
nor U7512 (N_7512,N_7444,N_7038);
and U7513 (N_7513,N_6981,N_6090);
and U7514 (N_7514,N_6733,N_6801);
xnor U7515 (N_7515,N_6336,N_7300);
nor U7516 (N_7516,N_6767,N_7497);
or U7517 (N_7517,N_7454,N_6937);
or U7518 (N_7518,N_7187,N_6309);
nor U7519 (N_7519,N_6396,N_6757);
nor U7520 (N_7520,N_7081,N_7101);
or U7521 (N_7521,N_6318,N_7198);
nor U7522 (N_7522,N_6067,N_7111);
nand U7523 (N_7523,N_6059,N_7359);
xor U7524 (N_7524,N_6601,N_6101);
xor U7525 (N_7525,N_6746,N_6291);
xor U7526 (N_7526,N_7115,N_7186);
nand U7527 (N_7527,N_6492,N_6949);
xnor U7528 (N_7528,N_6738,N_7455);
xnor U7529 (N_7529,N_6139,N_6326);
nand U7530 (N_7530,N_6109,N_6648);
and U7531 (N_7531,N_6679,N_7469);
nand U7532 (N_7532,N_6382,N_7345);
nand U7533 (N_7533,N_6631,N_6510);
and U7534 (N_7534,N_6168,N_7217);
xor U7535 (N_7535,N_7292,N_6487);
nor U7536 (N_7536,N_6119,N_6924);
nand U7537 (N_7537,N_7388,N_7114);
and U7538 (N_7538,N_7471,N_6183);
or U7539 (N_7539,N_6297,N_7041);
and U7540 (N_7540,N_6349,N_6047);
nor U7541 (N_7541,N_7348,N_6609);
and U7542 (N_7542,N_7481,N_6445);
and U7543 (N_7543,N_6589,N_7383);
and U7544 (N_7544,N_6152,N_7456);
nor U7545 (N_7545,N_7441,N_7268);
and U7546 (N_7546,N_6706,N_6508);
nor U7547 (N_7547,N_6945,N_7299);
and U7548 (N_7548,N_6925,N_6319);
and U7549 (N_7549,N_7210,N_6192);
xor U7550 (N_7550,N_6365,N_7247);
nand U7551 (N_7551,N_6028,N_7403);
xnor U7552 (N_7552,N_6489,N_7160);
or U7553 (N_7553,N_6369,N_7037);
and U7554 (N_7554,N_6308,N_6677);
or U7555 (N_7555,N_6979,N_6082);
nor U7556 (N_7556,N_6624,N_6294);
or U7557 (N_7557,N_7404,N_6635);
xor U7558 (N_7558,N_6726,N_6507);
or U7559 (N_7559,N_7096,N_6091);
nor U7560 (N_7560,N_6418,N_6722);
nor U7561 (N_7561,N_7136,N_6633);
xor U7562 (N_7562,N_6840,N_6135);
xor U7563 (N_7563,N_6393,N_7201);
and U7564 (N_7564,N_6450,N_6640);
and U7565 (N_7565,N_7169,N_6831);
and U7566 (N_7566,N_7087,N_6138);
nor U7567 (N_7567,N_7306,N_7398);
nor U7568 (N_7568,N_6441,N_6752);
and U7569 (N_7569,N_7011,N_6343);
and U7570 (N_7570,N_7237,N_6477);
or U7571 (N_7571,N_6672,N_6426);
nand U7572 (N_7572,N_6879,N_6161);
xnor U7573 (N_7573,N_6904,N_6707);
xor U7574 (N_7574,N_7302,N_6035);
and U7575 (N_7575,N_6735,N_7421);
nand U7576 (N_7576,N_7168,N_6031);
or U7577 (N_7577,N_6381,N_6912);
nor U7578 (N_7578,N_7214,N_7050);
nand U7579 (N_7579,N_6121,N_7226);
xnor U7580 (N_7580,N_6743,N_6804);
nor U7581 (N_7581,N_7080,N_6357);
nand U7582 (N_7582,N_6780,N_6292);
nor U7583 (N_7583,N_6199,N_6252);
or U7584 (N_7584,N_6742,N_6802);
nand U7585 (N_7585,N_6040,N_6277);
nand U7586 (N_7586,N_6272,N_6874);
nor U7587 (N_7587,N_6200,N_7477);
nand U7588 (N_7588,N_7307,N_7466);
nand U7589 (N_7589,N_6570,N_6485);
and U7590 (N_7590,N_7233,N_6943);
nand U7591 (N_7591,N_7183,N_7155);
nand U7592 (N_7592,N_6709,N_6270);
or U7593 (N_7593,N_6600,N_6221);
or U7594 (N_7594,N_7392,N_7439);
nor U7595 (N_7595,N_6727,N_6156);
and U7596 (N_7596,N_7241,N_6258);
nand U7597 (N_7597,N_7377,N_7014);
or U7598 (N_7598,N_7109,N_6712);
nor U7599 (N_7599,N_6043,N_6212);
or U7600 (N_7600,N_6744,N_6875);
nand U7601 (N_7601,N_6269,N_6359);
xnor U7602 (N_7602,N_7303,N_6063);
xnor U7603 (N_7603,N_6339,N_6967);
or U7604 (N_7604,N_6867,N_6290);
nand U7605 (N_7605,N_7369,N_6254);
nand U7606 (N_7606,N_6122,N_6069);
and U7607 (N_7607,N_7132,N_6053);
nand U7608 (N_7608,N_6006,N_7026);
nor U7609 (N_7609,N_6375,N_6705);
or U7610 (N_7610,N_6584,N_7068);
or U7611 (N_7611,N_6900,N_6678);
or U7612 (N_7612,N_7364,N_7020);
nand U7613 (N_7613,N_6351,N_6658);
or U7614 (N_7614,N_7266,N_6021);
nand U7615 (N_7615,N_6986,N_6453);
xnor U7616 (N_7616,N_6203,N_6926);
or U7617 (N_7617,N_7259,N_7270);
xnor U7618 (N_7618,N_7324,N_6358);
xor U7619 (N_7619,N_7039,N_6009);
nand U7620 (N_7620,N_7427,N_6230);
xnor U7621 (N_7621,N_6284,N_6264);
nand U7622 (N_7622,N_6923,N_6094);
nor U7623 (N_7623,N_6467,N_6494);
nor U7624 (N_7624,N_6675,N_6253);
xor U7625 (N_7625,N_6545,N_6194);
xor U7626 (N_7626,N_6348,N_6894);
or U7627 (N_7627,N_6054,N_6603);
or U7628 (N_7628,N_6162,N_7119);
or U7629 (N_7629,N_6626,N_7298);
nor U7630 (N_7630,N_7476,N_6449);
xnor U7631 (N_7631,N_7229,N_6927);
xor U7632 (N_7632,N_6907,N_6583);
and U7633 (N_7633,N_6863,N_6432);
xor U7634 (N_7634,N_6618,N_6990);
and U7635 (N_7635,N_6577,N_7128);
xnor U7636 (N_7636,N_6548,N_7488);
nand U7637 (N_7637,N_7148,N_7432);
or U7638 (N_7638,N_7293,N_6792);
nand U7639 (N_7639,N_7326,N_6881);
or U7640 (N_7640,N_6224,N_6946);
or U7641 (N_7641,N_7443,N_6242);
nand U7642 (N_7642,N_6092,N_6022);
nand U7643 (N_7643,N_6807,N_6887);
nor U7644 (N_7644,N_6516,N_7277);
and U7645 (N_7645,N_7204,N_6182);
and U7646 (N_7646,N_6773,N_6352);
or U7647 (N_7647,N_7437,N_7314);
xor U7648 (N_7648,N_7106,N_6049);
and U7649 (N_7649,N_6632,N_6276);
nand U7650 (N_7650,N_7116,N_6234);
and U7651 (N_7651,N_6698,N_6715);
or U7652 (N_7652,N_6565,N_6533);
nor U7653 (N_7653,N_6651,N_6615);
and U7654 (N_7654,N_7336,N_6419);
nand U7655 (N_7655,N_6935,N_7342);
nand U7656 (N_7656,N_6806,N_7405);
or U7657 (N_7657,N_6231,N_6643);
nand U7658 (N_7658,N_6197,N_6141);
or U7659 (N_7659,N_7166,N_7353);
nor U7660 (N_7660,N_7227,N_6273);
nor U7661 (N_7661,N_6888,N_6446);
or U7662 (N_7662,N_7375,N_7366);
and U7663 (N_7663,N_6066,N_6072);
and U7664 (N_7664,N_6576,N_6033);
and U7665 (N_7665,N_6826,N_6535);
or U7666 (N_7666,N_6262,N_6560);
and U7667 (N_7667,N_6997,N_6951);
nor U7668 (N_7668,N_7249,N_6649);
xnor U7669 (N_7669,N_6886,N_7315);
nor U7670 (N_7670,N_6263,N_6719);
nand U7671 (N_7671,N_7018,N_7117);
and U7672 (N_7672,N_7275,N_6282);
or U7673 (N_7673,N_6172,N_7190);
xor U7674 (N_7674,N_7489,N_6641);
nand U7675 (N_7675,N_6266,N_6922);
or U7676 (N_7676,N_6459,N_6984);
nor U7677 (N_7677,N_7154,N_6112);
nor U7678 (N_7678,N_7402,N_6580);
nor U7679 (N_7679,N_6051,N_6730);
and U7680 (N_7680,N_7023,N_7258);
nand U7681 (N_7681,N_6865,N_6146);
nor U7682 (N_7682,N_6233,N_7180);
nand U7683 (N_7683,N_7007,N_7250);
nor U7684 (N_7684,N_6469,N_6283);
nor U7685 (N_7685,N_6075,N_7222);
nor U7686 (N_7686,N_6686,N_6612);
nand U7687 (N_7687,N_6753,N_7341);
or U7688 (N_7688,N_6448,N_6324);
nor U7689 (N_7689,N_6171,N_6760);
xnor U7690 (N_7690,N_7086,N_7122);
and U7691 (N_7691,N_6607,N_6519);
xnor U7692 (N_7692,N_6818,N_7358);
nand U7693 (N_7693,N_7487,N_7478);
or U7694 (N_7694,N_6205,N_6003);
xnor U7695 (N_7695,N_6454,N_7009);
xnor U7696 (N_7696,N_6041,N_6980);
xnor U7697 (N_7697,N_6341,N_6064);
nand U7698 (N_7698,N_6963,N_7351);
nor U7699 (N_7699,N_7267,N_6741);
xor U7700 (N_7700,N_6256,N_6137);
nand U7701 (N_7701,N_6097,N_6598);
and U7702 (N_7702,N_6196,N_6206);
and U7703 (N_7703,N_6713,N_7135);
xnor U7704 (N_7704,N_6910,N_7442);
nand U7705 (N_7705,N_7378,N_6825);
and U7706 (N_7706,N_6364,N_6209);
nor U7707 (N_7707,N_6638,N_7093);
and U7708 (N_7708,N_7322,N_6895);
nor U7709 (N_7709,N_7418,N_6045);
xnor U7710 (N_7710,N_7460,N_6915);
xnor U7711 (N_7711,N_6856,N_7486);
nor U7712 (N_7712,N_7173,N_6655);
xor U7713 (N_7713,N_7124,N_6968);
or U7714 (N_7714,N_7269,N_7446);
or U7715 (N_7715,N_6311,N_6559);
nand U7716 (N_7716,N_7063,N_6439);
nor U7717 (N_7717,N_6656,N_6662);
and U7718 (N_7718,N_7339,N_6739);
or U7719 (N_7719,N_7057,N_7414);
nand U7720 (N_7720,N_7045,N_6764);
and U7721 (N_7721,N_7447,N_6346);
nand U7722 (N_7722,N_7458,N_6646);
xor U7723 (N_7723,N_6571,N_6794);
xor U7724 (N_7724,N_7098,N_6186);
nand U7725 (N_7725,N_7196,N_6244);
nand U7726 (N_7726,N_6717,N_7029);
nand U7727 (N_7727,N_7436,N_6301);
and U7728 (N_7728,N_7246,N_7327);
or U7729 (N_7729,N_6330,N_6239);
or U7730 (N_7730,N_6288,N_7301);
nand U7731 (N_7731,N_6541,N_7271);
nand U7732 (N_7732,N_6890,N_6971);
nand U7733 (N_7733,N_7376,N_6827);
and U7734 (N_7734,N_7467,N_7102);
xor U7735 (N_7735,N_6473,N_6718);
or U7736 (N_7736,N_7012,N_6666);
nor U7737 (N_7737,N_6249,N_6157);
and U7738 (N_7738,N_6564,N_6914);
and U7739 (N_7739,N_6383,N_6228);
xor U7740 (N_7740,N_6399,N_6246);
and U7741 (N_7741,N_6563,N_6538);
and U7742 (N_7742,N_7395,N_7239);
or U7743 (N_7743,N_6460,N_6562);
xnor U7744 (N_7744,N_7197,N_7162);
xor U7745 (N_7745,N_6782,N_6514);
nand U7746 (N_7746,N_6880,N_6855);
or U7747 (N_7747,N_7094,N_6065);
nor U7748 (N_7748,N_6251,N_6398);
nand U7749 (N_7749,N_7017,N_6464);
or U7750 (N_7750,N_7043,N_6474);
nand U7751 (N_7751,N_6745,N_6384);
xor U7752 (N_7752,N_7084,N_6850);
nand U7753 (N_7753,N_6405,N_6496);
and U7754 (N_7754,N_6227,N_7123);
nor U7755 (N_7755,N_6594,N_7044);
nand U7756 (N_7756,N_6755,N_6777);
or U7757 (N_7757,N_6201,N_7046);
or U7758 (N_7758,N_7372,N_7479);
nor U7759 (N_7759,N_7363,N_7408);
or U7760 (N_7760,N_7199,N_6805);
or U7761 (N_7761,N_7289,N_7031);
nand U7762 (N_7762,N_7099,N_6312);
xnor U7763 (N_7763,N_6593,N_6068);
nand U7764 (N_7764,N_6518,N_6847);
nor U7765 (N_7765,N_6702,N_6965);
xor U7766 (N_7766,N_6761,N_6370);
and U7767 (N_7767,N_7416,N_7420);
xor U7768 (N_7768,N_7498,N_6768);
nand U7769 (N_7769,N_6431,N_6160);
nor U7770 (N_7770,N_6824,N_6440);
and U7771 (N_7771,N_6353,N_6788);
nor U7772 (N_7772,N_6355,N_6634);
and U7773 (N_7773,N_7272,N_6081);
nor U7774 (N_7774,N_6588,N_6150);
and U7775 (N_7775,N_6837,N_6173);
xor U7776 (N_7776,N_6941,N_6750);
nand U7777 (N_7777,N_7105,N_6578);
and U7778 (N_7778,N_6653,N_6340);
or U7779 (N_7779,N_6463,N_6822);
or U7780 (N_7780,N_6958,N_6723);
and U7781 (N_7781,N_7473,N_6857);
xor U7782 (N_7782,N_6211,N_7433);
nand U7783 (N_7783,N_6388,N_7244);
nand U7784 (N_7784,N_7278,N_6223);
or U7785 (N_7785,N_6002,N_6621);
or U7786 (N_7786,N_6749,N_7354);
nand U7787 (N_7787,N_7205,N_7171);
xor U7788 (N_7788,N_7357,N_6959);
nand U7789 (N_7789,N_6556,N_7185);
or U7790 (N_7790,N_6088,N_7113);
xor U7791 (N_7791,N_6151,N_7151);
or U7792 (N_7792,N_6052,N_6004);
xnor U7793 (N_7793,N_6279,N_6547);
and U7794 (N_7794,N_6862,N_6637);
or U7795 (N_7795,N_7368,N_7318);
xnor U7796 (N_7796,N_6903,N_6126);
and U7797 (N_7797,N_6079,N_6245);
nor U7798 (N_7798,N_6501,N_7330);
nand U7799 (N_7799,N_6046,N_6729);
nand U7800 (N_7800,N_7328,N_6710);
or U7801 (N_7801,N_6188,N_7110);
xor U7802 (N_7802,N_6697,N_7282);
xnor U7803 (N_7803,N_7143,N_7255);
xor U7804 (N_7804,N_6178,N_6229);
xnor U7805 (N_7805,N_6165,N_7073);
or U7806 (N_7806,N_7200,N_6933);
or U7807 (N_7807,N_6861,N_7193);
or U7808 (N_7808,N_7248,N_6839);
xnor U7809 (N_7809,N_6363,N_7323);
nand U7810 (N_7810,N_7465,N_7156);
xnor U7811 (N_7811,N_6295,N_6969);
xnor U7812 (N_7812,N_7228,N_6766);
or U7813 (N_7813,N_6176,N_6549);
or U7814 (N_7814,N_6608,N_6740);
xnor U7815 (N_7815,N_6934,N_7426);
xnor U7816 (N_7816,N_7361,N_7265);
xor U7817 (N_7817,N_6572,N_6599);
and U7818 (N_7818,N_7344,N_7161);
or U7819 (N_7819,N_6829,N_7371);
nor U7820 (N_7820,N_6523,N_6032);
xnor U7821 (N_7821,N_7220,N_6846);
or U7822 (N_7822,N_6521,N_6978);
and U7823 (N_7823,N_7066,N_7047);
xnor U7824 (N_7824,N_6387,N_6403);
or U7825 (N_7825,N_6701,N_7313);
nor U7826 (N_7826,N_7243,N_6397);
nand U7827 (N_7827,N_6763,N_6498);
nor U7828 (N_7828,N_6402,N_6567);
nor U7829 (N_7829,N_6869,N_6614);
and U7830 (N_7830,N_6669,N_6333);
xnor U7831 (N_7831,N_6404,N_6106);
or U7832 (N_7832,N_6784,N_7022);
nor U7833 (N_7833,N_6281,N_7212);
nand U7834 (N_7834,N_6039,N_6342);
nand U7835 (N_7835,N_7312,N_6015);
nor U7836 (N_7836,N_6622,N_6430);
or U7837 (N_7837,N_6191,N_6823);
nand U7838 (N_7838,N_6232,N_6235);
or U7839 (N_7839,N_6013,N_6882);
nor U7840 (N_7840,N_7449,N_7085);
xor U7841 (N_7841,N_7253,N_6596);
nand U7842 (N_7842,N_6703,N_6293);
or U7843 (N_7843,N_6202,N_7429);
nor U7844 (N_7844,N_6849,N_6468);
nand U7845 (N_7845,N_6005,N_7251);
or U7846 (N_7846,N_6982,N_6424);
xor U7847 (N_7847,N_7349,N_6630);
or U7848 (N_7848,N_7131,N_6329);
nor U7849 (N_7849,N_6858,N_6406);
xnor U7850 (N_7850,N_7474,N_6483);
nand U7851 (N_7851,N_6007,N_6217);
and U7852 (N_7852,N_7355,N_6964);
nor U7853 (N_7853,N_7015,N_6144);
nor U7854 (N_7854,N_6321,N_6841);
nor U7855 (N_7855,N_6975,N_6673);
nor U7856 (N_7856,N_7075,N_6660);
xor U7857 (N_7857,N_6055,N_7380);
nand U7858 (N_7858,N_7033,N_6555);
nand U7859 (N_7859,N_7095,N_6167);
nand U7860 (N_7860,N_7415,N_7054);
nor U7861 (N_7861,N_7192,N_7352);
and U7862 (N_7862,N_6378,N_6961);
nor U7863 (N_7863,N_6616,N_7338);
nand U7864 (N_7864,N_6307,N_6852);
nor U7865 (N_7865,N_6238,N_6117);
or U7866 (N_7866,N_6215,N_6736);
nor U7867 (N_7867,N_7107,N_6193);
nor U7868 (N_7868,N_7202,N_6917);
and U7869 (N_7869,N_7211,N_6808);
nor U7870 (N_7870,N_6667,N_6268);
nand U7871 (N_7871,N_7092,N_6073);
and U7872 (N_7872,N_7310,N_6948);
nor U7873 (N_7873,N_6663,N_6606);
or U7874 (N_7874,N_6765,N_6956);
and U7875 (N_7875,N_6019,N_6970);
nor U7876 (N_7876,N_6048,N_6020);
and U7877 (N_7877,N_6434,N_7382);
and U7878 (N_7878,N_6195,N_7386);
or U7879 (N_7879,N_6939,N_6558);
nand U7880 (N_7880,N_6619,N_7482);
nand U7881 (N_7881,N_7295,N_6711);
nor U7882 (N_7882,N_6762,N_7280);
nand U7883 (N_7883,N_7316,N_6107);
nand U7884 (N_7884,N_6524,N_7000);
nand U7885 (N_7885,N_6931,N_6198);
nor U7886 (N_7886,N_6298,N_6515);
xnor U7887 (N_7887,N_6386,N_6422);
nor U7888 (N_7888,N_6991,N_6134);
xnor U7889 (N_7889,N_6581,N_6795);
nand U7890 (N_7890,N_7157,N_6532);
xnor U7891 (N_7891,N_6790,N_7133);
or U7892 (N_7892,N_6164,N_6550);
xor U7893 (N_7893,N_6942,N_6680);
nor U7894 (N_7894,N_6169,N_7459);
xnor U7895 (N_7895,N_7231,N_6810);
or U7896 (N_7896,N_7373,N_6906);
nor U7897 (N_7897,N_7142,N_7141);
xor U7898 (N_7898,N_6366,N_7067);
and U7899 (N_7899,N_6690,N_6921);
and U7900 (N_7900,N_6687,N_6305);
or U7901 (N_7901,N_6148,N_6350);
nor U7902 (N_7902,N_6783,N_7317);
nor U7903 (N_7903,N_7195,N_6685);
nand U7904 (N_7904,N_6287,N_6415);
and U7905 (N_7905,N_7125,N_6682);
nor U7906 (N_7906,N_6327,N_7036);
and U7907 (N_7907,N_7129,N_6930);
and U7908 (N_7908,N_6732,N_6642);
and U7909 (N_7909,N_6300,N_7130);
or U7910 (N_7910,N_6681,N_7146);
nand U7911 (N_7911,N_7091,N_7194);
or U7912 (N_7912,N_6377,N_7242);
xnor U7913 (N_7913,N_7283,N_7396);
or U7914 (N_7914,N_6796,N_6458);
or U7915 (N_7915,N_6337,N_7288);
nand U7916 (N_7916,N_6530,N_6095);
and U7917 (N_7917,N_7181,N_7435);
xor U7918 (N_7918,N_7191,N_7118);
nor U7919 (N_7919,N_6481,N_6136);
nor U7920 (N_7920,N_6758,N_7490);
and U7921 (N_7921,N_6989,N_6983);
nor U7922 (N_7922,N_6361,N_6255);
nand U7923 (N_7923,N_6817,N_6502);
and U7924 (N_7924,N_6512,N_6360);
and U7925 (N_7925,N_7216,N_7296);
xnor U7926 (N_7926,N_7175,N_6845);
and U7927 (N_7927,N_7016,N_7240);
or U7928 (N_7928,N_6799,N_7438);
or U7929 (N_7929,N_7021,N_6798);
xnor U7930 (N_7930,N_6409,N_7385);
nor U7931 (N_7931,N_6960,N_6411);
or U7932 (N_7932,N_6950,N_6362);
and U7933 (N_7933,N_6511,N_6017);
nor U7934 (N_7934,N_6820,N_6816);
nand U7935 (N_7935,N_7400,N_6476);
nand U7936 (N_7936,N_7367,N_6976);
nand U7937 (N_7937,N_7281,N_7172);
nand U7938 (N_7938,N_6553,N_7005);
nor U7939 (N_7939,N_6400,N_6695);
nand U7940 (N_7940,N_6617,N_6901);
and U7941 (N_7941,N_6423,N_6814);
or U7942 (N_7942,N_7064,N_7472);
xor U7943 (N_7943,N_6522,N_6551);
nor U7944 (N_7944,N_6071,N_7165);
and U7945 (N_7945,N_6985,N_7484);
nand U7946 (N_7946,N_6480,N_6708);
and U7947 (N_7947,N_7399,N_6417);
xnor U7948 (N_7948,N_7079,N_6602);
xnor U7949 (N_7949,N_7496,N_6591);
and U7950 (N_7950,N_6836,N_6163);
or U7951 (N_7951,N_6566,N_6133);
and U7952 (N_7952,N_6661,N_6592);
xor U7953 (N_7953,N_7139,N_7207);
and U7954 (N_7954,N_7097,N_7234);
or U7955 (N_7955,N_6528,N_6586);
nor U7956 (N_7956,N_6243,N_6513);
nor U7957 (N_7957,N_7053,N_6693);
or U7958 (N_7958,N_6652,N_7008);
xor U7959 (N_7959,N_7208,N_6219);
nand U7960 (N_7960,N_7035,N_6833);
xnor U7961 (N_7961,N_6466,N_7491);
and U7962 (N_7962,N_6775,N_6442);
and U7963 (N_7963,N_6026,N_6143);
nor U7964 (N_7964,N_6728,N_6093);
xnor U7965 (N_7965,N_7406,N_6158);
xnor U7966 (N_7966,N_6414,N_6016);
xor U7967 (N_7967,N_7218,N_7356);
nor U7968 (N_7968,N_6647,N_6873);
nand U7969 (N_7969,N_6789,N_6770);
or U7970 (N_7970,N_6316,N_7411);
or U7971 (N_7971,N_6147,N_7422);
xnor U7972 (N_7972,N_6470,N_7370);
nor U7973 (N_7973,N_6170,N_6210);
nor U7974 (N_7974,N_7027,N_6145);
and U7975 (N_7975,N_6385,N_7453);
nand U7976 (N_7976,N_7457,N_6813);
or U7977 (N_7977,N_6771,N_6714);
nand U7978 (N_7978,N_6132,N_6056);
nand U7979 (N_7979,N_6944,N_7410);
nand U7980 (N_7980,N_6499,N_7089);
and U7981 (N_7981,N_7167,N_7276);
or U7982 (N_7982,N_7252,N_6654);
xor U7983 (N_7983,N_6379,N_6042);
nor U7984 (N_7984,N_6838,N_7127);
xnor U7985 (N_7985,N_7365,N_7287);
xor U7986 (N_7986,N_6407,N_6380);
or U7987 (N_7987,N_7209,N_6843);
or U7988 (N_7988,N_7311,N_6275);
xnor U7989 (N_7989,N_6992,N_6853);
nor U7990 (N_7990,N_7056,N_6070);
and U7991 (N_7991,N_7034,N_7179);
and U7992 (N_7992,N_6484,N_7235);
nor U7993 (N_7993,N_6394,N_7335);
nor U7994 (N_7994,N_7189,N_6676);
xor U7995 (N_7995,N_6204,N_6500);
nor U7996 (N_7996,N_6911,N_7077);
nor U7997 (N_7997,N_6437,N_7028);
or U7998 (N_7998,N_7103,N_7319);
nand U7999 (N_7999,N_7174,N_6475);
nor U8000 (N_8000,N_7448,N_7176);
and U8001 (N_8001,N_6936,N_6885);
nand U8002 (N_8002,N_7412,N_6552);
nand U8003 (N_8003,N_6062,N_7452);
nor U8004 (N_8004,N_6103,N_6462);
xor U8005 (N_8005,N_7078,N_6089);
and U8006 (N_8006,N_6320,N_7480);
and U8007 (N_8007,N_6725,N_6561);
or U8008 (N_8008,N_6902,N_7121);
xnor U8009 (N_8009,N_7391,N_6889);
nand U8010 (N_8010,N_6142,N_6317);
or U8011 (N_8011,N_7256,N_6060);
xnor U8012 (N_8012,N_7334,N_7393);
nor U8013 (N_8013,N_6389,N_6113);
nor U8014 (N_8014,N_6140,N_7413);
nand U8015 (N_8015,N_7245,N_7230);
xor U8016 (N_8016,N_7048,N_6898);
and U8017 (N_8017,N_6325,N_6259);
and U8018 (N_8018,N_6977,N_7049);
nor U8019 (N_8019,N_7264,N_7213);
and U8020 (N_8020,N_6118,N_6720);
xnor U8021 (N_8021,N_6408,N_6962);
nand U8022 (N_8022,N_7360,N_7425);
nor U8023 (N_8023,N_6525,N_7450);
xor U8024 (N_8024,N_6668,N_7333);
or U8025 (N_8025,N_6787,N_6876);
xnor U8026 (N_8026,N_6368,N_6213);
or U8027 (N_8027,N_7010,N_7042);
nand U8028 (N_8028,N_7188,N_6897);
xnor U8029 (N_8029,N_6310,N_6769);
nand U8030 (N_8030,N_6038,N_6010);
nor U8031 (N_8031,N_6410,N_6313);
xnor U8032 (N_8032,N_6896,N_6947);
nor U8033 (N_8033,N_6250,N_6125);
and U8034 (N_8034,N_6776,N_7002);
xnor U8035 (N_8035,N_7494,N_6265);
nor U8036 (N_8036,N_6689,N_7284);
xor U8037 (N_8037,N_6568,N_7178);
or U8038 (N_8038,N_7219,N_6529);
and U8039 (N_8039,N_7177,N_7431);
or U8040 (N_8040,N_6546,N_6175);
xor U8041 (N_8041,N_7381,N_6891);
or U8042 (N_8042,N_6573,N_6057);
xnor U8043 (N_8043,N_7238,N_6999);
nand U8044 (N_8044,N_6108,N_7100);
or U8045 (N_8045,N_6299,N_6104);
xor U8046 (N_8046,N_6694,N_6893);
xor U8047 (N_8047,N_6884,N_6998);
xnor U8048 (N_8048,N_6216,N_6554);
and U8049 (N_8049,N_7331,N_6916);
nor U8050 (N_8050,N_6683,N_7428);
nand U8051 (N_8051,N_6665,N_6105);
and U8052 (N_8052,N_7024,N_7260);
xor U8053 (N_8053,N_7285,N_6373);
xnor U8054 (N_8054,N_6471,N_6344);
and U8055 (N_8055,N_7062,N_7164);
xnor U8056 (N_8056,N_6037,N_6582);
xor U8057 (N_8057,N_6084,N_7030);
xor U8058 (N_8058,N_6190,N_6692);
or U8059 (N_8059,N_6208,N_7158);
nand U8060 (N_8060,N_6303,N_6124);
nand U8061 (N_8061,N_6627,N_7499);
and U8062 (N_8062,N_7140,N_6261);
nor U8063 (N_8063,N_7321,N_6100);
and U8064 (N_8064,N_7138,N_7374);
or U8065 (N_8065,N_7419,N_6401);
or U8066 (N_8066,N_6751,N_7145);
nand U8067 (N_8067,N_6664,N_6443);
and U8068 (N_8068,N_6030,N_7223);
or U8069 (N_8069,N_6447,N_6000);
and U8070 (N_8070,N_7401,N_6018);
xor U8071 (N_8071,N_7051,N_6280);
or U8072 (N_8072,N_6332,N_6367);
or U8073 (N_8073,N_6639,N_6236);
nand U8074 (N_8074,N_7350,N_6899);
or U8075 (N_8075,N_7309,N_6785);
xnor U8076 (N_8076,N_6848,N_6323);
or U8077 (N_8077,N_7254,N_6304);
and U8078 (N_8078,N_7058,N_6868);
nand U8079 (N_8079,N_7379,N_6731);
xor U8080 (N_8080,N_6008,N_6854);
or U8081 (N_8081,N_6800,N_6786);
or U8082 (N_8082,N_7083,N_6864);
nor U8083 (N_8083,N_6044,N_6809);
nor U8084 (N_8084,N_6892,N_6908);
nor U8085 (N_8085,N_6179,N_6472);
or U8086 (N_8086,N_6425,N_6579);
and U8087 (N_8087,N_6486,N_6835);
and U8088 (N_8088,N_6877,N_6077);
nand U8089 (N_8089,N_6438,N_7003);
nand U8090 (N_8090,N_6534,N_6842);
and U8091 (N_8091,N_6756,N_6575);
nor U8092 (N_8092,N_6154,N_6435);
nand U8093 (N_8093,N_6478,N_7290);
and U8094 (N_8094,N_6083,N_6180);
nand U8095 (N_8095,N_6174,N_7040);
nor U8096 (N_8096,N_6153,N_6127);
nand U8097 (N_8097,N_7144,N_6098);
nor U8098 (N_8098,N_6955,N_6356);
or U8099 (N_8099,N_6257,N_6932);
xor U8100 (N_8100,N_6286,N_6347);
or U8101 (N_8101,N_6114,N_7387);
nand U8102 (N_8102,N_6605,N_6306);
xnor U8103 (N_8103,N_7409,N_6954);
xor U8104 (N_8104,N_6050,N_6670);
or U8105 (N_8105,N_6928,N_6096);
xnor U8106 (N_8106,N_6260,N_6428);
nor U8107 (N_8107,N_6011,N_7052);
or U8108 (N_8108,N_6920,N_6421);
and U8109 (N_8109,N_6509,N_6338);
and U8110 (N_8110,N_6451,N_6110);
or U8111 (N_8111,N_6335,N_6274);
and U8112 (N_8112,N_6866,N_6495);
nor U8113 (N_8113,N_7394,N_6078);
or U8114 (N_8114,N_6716,N_7088);
nand U8115 (N_8115,N_6748,N_6345);
nor U8116 (N_8116,N_7065,N_6116);
nor U8117 (N_8117,N_6721,N_6544);
and U8118 (N_8118,N_7163,N_6302);
nand U8119 (N_8119,N_6159,N_6613);
nor U8120 (N_8120,N_6166,N_6734);
nor U8121 (N_8121,N_6793,N_7006);
nor U8122 (N_8122,N_7362,N_7463);
nand U8123 (N_8123,N_7325,N_7308);
xor U8124 (N_8124,N_6747,N_6691);
or U8125 (N_8125,N_6207,N_6220);
xor U8126 (N_8126,N_6413,N_7470);
xnor U8127 (N_8127,N_6859,N_6754);
and U8128 (N_8128,N_6797,N_6688);
nand U8129 (N_8129,N_6058,N_7001);
nor U8130 (N_8130,N_7076,N_6779);
nor U8131 (N_8131,N_6267,N_6184);
nor U8132 (N_8132,N_6372,N_6420);
nand U8133 (N_8133,N_6131,N_6177);
and U8134 (N_8134,N_6611,N_7485);
nand U8135 (N_8135,N_6099,N_7424);
nand U8136 (N_8136,N_6629,N_6036);
nor U8137 (N_8137,N_6811,N_7072);
nor U8138 (N_8138,N_6871,N_6085);
and U8139 (N_8139,N_7468,N_6585);
nand U8140 (N_8140,N_6517,N_7430);
nand U8141 (N_8141,N_6953,N_6540);
xnor U8142 (N_8142,N_6181,N_6918);
nand U8143 (N_8143,N_7074,N_6938);
nand U8144 (N_8144,N_6737,N_7337);
nor U8145 (N_8145,N_7320,N_7294);
nor U8146 (N_8146,N_6322,N_7407);
or U8147 (N_8147,N_6023,N_6416);
and U8148 (N_8148,N_6929,N_7120);
or U8149 (N_8149,N_7347,N_7215);
and U8150 (N_8150,N_7232,N_6237);
or U8151 (N_8151,N_6456,N_6952);
nand U8152 (N_8152,N_6493,N_6832);
xor U8153 (N_8153,N_7332,N_6940);
and U8154 (N_8154,N_6644,N_6189);
nor U8155 (N_8155,N_6289,N_7286);
or U8156 (N_8156,N_6812,N_7149);
nor U8157 (N_8157,N_6684,N_7273);
and U8158 (N_8158,N_6391,N_6129);
and U8159 (N_8159,N_7104,N_7025);
nor U8160 (N_8160,N_6995,N_6569);
nand U8161 (N_8161,N_7423,N_6328);
xnor U8162 (N_8162,N_6455,N_7493);
or U8163 (N_8163,N_6427,N_6791);
nand U8164 (N_8164,N_6781,N_7224);
nor U8165 (N_8165,N_6505,N_6974);
nor U8166 (N_8166,N_7462,N_7203);
nor U8167 (N_8167,N_7305,N_6543);
and U8168 (N_8168,N_6029,N_6815);
xnor U8169 (N_8169,N_6061,N_7182);
nor U8170 (N_8170,N_6128,N_6604);
or U8171 (N_8171,N_6883,N_7343);
xnor U8172 (N_8172,N_7112,N_6527);
xor U8173 (N_8173,N_7346,N_6074);
nand U8174 (N_8174,N_6436,N_7032);
or U8175 (N_8175,N_6870,N_7384);
and U8176 (N_8176,N_6285,N_6241);
nand U8177 (N_8177,N_6659,N_7070);
xor U8178 (N_8178,N_6699,N_6149);
and U8179 (N_8179,N_7262,N_6296);
xor U8180 (N_8180,N_7390,N_6130);
nor U8181 (N_8181,N_6392,N_7069);
and U8182 (N_8182,N_6395,N_6972);
xnor U8183 (N_8183,N_7274,N_6479);
nand U8184 (N_8184,N_6504,N_7060);
xnor U8185 (N_8185,N_6778,N_6860);
nand U8186 (N_8186,N_6025,N_6772);
or U8187 (N_8187,N_6671,N_6590);
nor U8188 (N_8188,N_6490,N_7055);
or U8189 (N_8189,N_6587,N_6657);
nor U8190 (N_8190,N_6531,N_6595);
nor U8191 (N_8191,N_7184,N_7013);
and U8192 (N_8192,N_7492,N_7329);
nand U8193 (N_8193,N_6185,N_6354);
nand U8194 (N_8194,N_6774,N_6488);
nor U8195 (N_8195,N_7159,N_6957);
nand U8196 (N_8196,N_7170,N_6724);
or U8197 (N_8197,N_7261,N_6087);
nand U8198 (N_8198,N_7451,N_7464);
or U8199 (N_8199,N_7483,N_7417);
nand U8200 (N_8200,N_6429,N_6123);
xor U8201 (N_8201,N_6996,N_6444);
or U8202 (N_8202,N_6905,N_6819);
nand U8203 (N_8203,N_7279,N_6526);
or U8204 (N_8204,N_6828,N_6315);
xor U8205 (N_8205,N_7440,N_7071);
nand U8206 (N_8206,N_6620,N_6187);
nor U8207 (N_8207,N_6821,N_6376);
or U8208 (N_8208,N_6465,N_7108);
nand U8209 (N_8209,N_6271,N_7082);
xnor U8210 (N_8210,N_6506,N_6645);
xnor U8211 (N_8211,N_7225,N_7304);
nand U8212 (N_8212,N_6919,N_6214);
nor U8213 (N_8213,N_6704,N_6014);
or U8214 (N_8214,N_6557,N_6610);
and U8215 (N_8215,N_6650,N_6331);
and U8216 (N_8216,N_6503,N_6542);
or U8217 (N_8217,N_6696,N_6314);
xnor U8218 (N_8218,N_6334,N_7291);
and U8219 (N_8219,N_6027,N_6247);
xnor U8220 (N_8220,N_6222,N_6120);
or U8221 (N_8221,N_6034,N_6993);
nand U8222 (N_8222,N_6491,N_6390);
nor U8223 (N_8223,N_7126,N_6537);
nand U8224 (N_8224,N_6913,N_6076);
nor U8225 (N_8225,N_6012,N_7257);
nor U8226 (N_8226,N_6433,N_6628);
xnor U8227 (N_8227,N_6878,N_6574);
and U8228 (N_8228,N_7434,N_6225);
nor U8229 (N_8229,N_7445,N_6452);
nor U8230 (N_8230,N_6830,N_7153);
xnor U8231 (N_8231,N_6080,N_6482);
xor U8232 (N_8232,N_7090,N_6623);
nand U8233 (N_8233,N_6636,N_7461);
and U8234 (N_8234,N_7134,N_7495);
xnor U8235 (N_8235,N_6994,N_6457);
xnor U8236 (N_8236,N_6966,N_6102);
xor U8237 (N_8237,N_6872,N_6461);
nand U8238 (N_8238,N_7137,N_6520);
and U8239 (N_8239,N_6597,N_6497);
nor U8240 (N_8240,N_6674,N_7147);
or U8241 (N_8241,N_7059,N_6155);
and U8242 (N_8242,N_6226,N_6278);
and U8243 (N_8243,N_7061,N_7221);
or U8244 (N_8244,N_7389,N_6987);
or U8245 (N_8245,N_6700,N_6240);
xor U8246 (N_8246,N_6851,N_6412);
nand U8247 (N_8247,N_7004,N_7475);
or U8248 (N_8248,N_6909,N_6218);
and U8249 (N_8249,N_6988,N_6536);
xor U8250 (N_8250,N_6889,N_6439);
xnor U8251 (N_8251,N_6126,N_6298);
xor U8252 (N_8252,N_6868,N_6074);
nand U8253 (N_8253,N_6503,N_7240);
nand U8254 (N_8254,N_6934,N_7253);
and U8255 (N_8255,N_7058,N_7042);
or U8256 (N_8256,N_6411,N_7394);
xnor U8257 (N_8257,N_6467,N_6244);
xnor U8258 (N_8258,N_6854,N_6690);
nor U8259 (N_8259,N_6137,N_6080);
xor U8260 (N_8260,N_7215,N_6653);
nand U8261 (N_8261,N_7425,N_6086);
nand U8262 (N_8262,N_7023,N_6520);
nand U8263 (N_8263,N_6937,N_6740);
xnor U8264 (N_8264,N_6287,N_7279);
and U8265 (N_8265,N_6387,N_6700);
nor U8266 (N_8266,N_6124,N_7135);
and U8267 (N_8267,N_6458,N_7069);
and U8268 (N_8268,N_6346,N_7209);
nand U8269 (N_8269,N_6178,N_6503);
nor U8270 (N_8270,N_7459,N_7135);
nand U8271 (N_8271,N_6422,N_7404);
nand U8272 (N_8272,N_6486,N_7044);
nand U8273 (N_8273,N_6407,N_7355);
and U8274 (N_8274,N_6931,N_7268);
nand U8275 (N_8275,N_6243,N_6566);
or U8276 (N_8276,N_6030,N_6662);
nor U8277 (N_8277,N_7216,N_6992);
and U8278 (N_8278,N_6343,N_6179);
xnor U8279 (N_8279,N_6931,N_6604);
and U8280 (N_8280,N_6783,N_6202);
and U8281 (N_8281,N_6033,N_6578);
or U8282 (N_8282,N_7158,N_6877);
nand U8283 (N_8283,N_7303,N_6563);
and U8284 (N_8284,N_6032,N_6734);
nand U8285 (N_8285,N_6701,N_6747);
and U8286 (N_8286,N_6541,N_7287);
and U8287 (N_8287,N_6967,N_7368);
and U8288 (N_8288,N_6871,N_7201);
and U8289 (N_8289,N_6892,N_6909);
or U8290 (N_8290,N_7323,N_6755);
or U8291 (N_8291,N_7359,N_6539);
xnor U8292 (N_8292,N_6051,N_6008);
nor U8293 (N_8293,N_6784,N_6548);
nand U8294 (N_8294,N_6870,N_7188);
nor U8295 (N_8295,N_7123,N_6532);
xor U8296 (N_8296,N_6040,N_7467);
and U8297 (N_8297,N_7036,N_6311);
xor U8298 (N_8298,N_6196,N_7423);
nand U8299 (N_8299,N_6788,N_7056);
or U8300 (N_8300,N_6315,N_6079);
or U8301 (N_8301,N_6194,N_7069);
or U8302 (N_8302,N_6253,N_6204);
nand U8303 (N_8303,N_6847,N_7138);
and U8304 (N_8304,N_6274,N_6569);
and U8305 (N_8305,N_7351,N_7224);
or U8306 (N_8306,N_6191,N_6183);
or U8307 (N_8307,N_6883,N_6256);
nand U8308 (N_8308,N_6012,N_6072);
nor U8309 (N_8309,N_6237,N_7392);
or U8310 (N_8310,N_7381,N_6369);
xnor U8311 (N_8311,N_6534,N_6962);
nand U8312 (N_8312,N_6006,N_7280);
and U8313 (N_8313,N_6246,N_6081);
xnor U8314 (N_8314,N_6192,N_6416);
xor U8315 (N_8315,N_6060,N_6450);
nor U8316 (N_8316,N_6948,N_6582);
nor U8317 (N_8317,N_6112,N_6357);
nor U8318 (N_8318,N_6791,N_6870);
nand U8319 (N_8319,N_7193,N_7300);
xor U8320 (N_8320,N_6110,N_6132);
or U8321 (N_8321,N_6053,N_6744);
nand U8322 (N_8322,N_7487,N_7300);
nand U8323 (N_8323,N_6265,N_6203);
or U8324 (N_8324,N_7191,N_6305);
and U8325 (N_8325,N_6531,N_6700);
xor U8326 (N_8326,N_6979,N_7031);
xor U8327 (N_8327,N_6866,N_7095);
xnor U8328 (N_8328,N_6395,N_7226);
or U8329 (N_8329,N_6378,N_6010);
and U8330 (N_8330,N_7398,N_6695);
and U8331 (N_8331,N_6321,N_6930);
xor U8332 (N_8332,N_7025,N_6661);
or U8333 (N_8333,N_6141,N_6649);
and U8334 (N_8334,N_6081,N_6041);
and U8335 (N_8335,N_7066,N_7027);
or U8336 (N_8336,N_6214,N_6783);
nand U8337 (N_8337,N_7008,N_6762);
or U8338 (N_8338,N_7083,N_7397);
and U8339 (N_8339,N_6436,N_6074);
nor U8340 (N_8340,N_6628,N_6794);
nand U8341 (N_8341,N_6710,N_7142);
xor U8342 (N_8342,N_6858,N_6047);
nand U8343 (N_8343,N_6211,N_7482);
xnor U8344 (N_8344,N_6289,N_7045);
and U8345 (N_8345,N_7306,N_6669);
nand U8346 (N_8346,N_6150,N_6781);
and U8347 (N_8347,N_7370,N_6435);
nor U8348 (N_8348,N_6291,N_7460);
nand U8349 (N_8349,N_6938,N_7058);
and U8350 (N_8350,N_6449,N_7013);
nand U8351 (N_8351,N_7388,N_6741);
or U8352 (N_8352,N_6382,N_7137);
xnor U8353 (N_8353,N_6084,N_6421);
or U8354 (N_8354,N_6448,N_6081);
nand U8355 (N_8355,N_7223,N_6371);
xor U8356 (N_8356,N_6656,N_7093);
xor U8357 (N_8357,N_7123,N_6956);
nand U8358 (N_8358,N_6120,N_6988);
xor U8359 (N_8359,N_6356,N_6462);
or U8360 (N_8360,N_7354,N_6944);
or U8361 (N_8361,N_6291,N_6233);
nand U8362 (N_8362,N_7225,N_6932);
xnor U8363 (N_8363,N_6460,N_6091);
nor U8364 (N_8364,N_6243,N_6555);
xor U8365 (N_8365,N_6160,N_6687);
and U8366 (N_8366,N_7235,N_6737);
or U8367 (N_8367,N_6647,N_6886);
and U8368 (N_8368,N_6106,N_7298);
xnor U8369 (N_8369,N_6066,N_6259);
and U8370 (N_8370,N_6242,N_6625);
nor U8371 (N_8371,N_6631,N_7386);
nor U8372 (N_8372,N_7358,N_7494);
or U8373 (N_8373,N_6274,N_6928);
or U8374 (N_8374,N_6408,N_6293);
or U8375 (N_8375,N_6534,N_6022);
nand U8376 (N_8376,N_7055,N_6172);
or U8377 (N_8377,N_6191,N_6372);
and U8378 (N_8378,N_7427,N_7139);
or U8379 (N_8379,N_6588,N_6501);
or U8380 (N_8380,N_6378,N_6503);
xnor U8381 (N_8381,N_6727,N_7214);
or U8382 (N_8382,N_7157,N_7308);
nor U8383 (N_8383,N_6199,N_7151);
nor U8384 (N_8384,N_6681,N_6645);
nor U8385 (N_8385,N_7041,N_6319);
nor U8386 (N_8386,N_7215,N_6147);
xnor U8387 (N_8387,N_7289,N_6631);
nor U8388 (N_8388,N_6188,N_6793);
and U8389 (N_8389,N_6966,N_7177);
nor U8390 (N_8390,N_6539,N_7196);
and U8391 (N_8391,N_6435,N_6381);
nand U8392 (N_8392,N_6403,N_6424);
or U8393 (N_8393,N_6632,N_6652);
xnor U8394 (N_8394,N_6198,N_6039);
nand U8395 (N_8395,N_6856,N_6013);
xnor U8396 (N_8396,N_7322,N_7415);
and U8397 (N_8397,N_7150,N_6400);
nand U8398 (N_8398,N_7155,N_6722);
or U8399 (N_8399,N_6592,N_6618);
nor U8400 (N_8400,N_6647,N_6724);
or U8401 (N_8401,N_6684,N_6484);
or U8402 (N_8402,N_7153,N_7318);
nor U8403 (N_8403,N_6290,N_6492);
nand U8404 (N_8404,N_6955,N_7226);
or U8405 (N_8405,N_7458,N_6749);
and U8406 (N_8406,N_6104,N_6062);
nor U8407 (N_8407,N_6288,N_7443);
nand U8408 (N_8408,N_6107,N_7044);
or U8409 (N_8409,N_7270,N_7214);
nor U8410 (N_8410,N_6335,N_6158);
nor U8411 (N_8411,N_6001,N_6099);
or U8412 (N_8412,N_7253,N_7133);
nand U8413 (N_8413,N_6999,N_6826);
xor U8414 (N_8414,N_6131,N_7326);
nand U8415 (N_8415,N_7179,N_7430);
xor U8416 (N_8416,N_6176,N_6638);
or U8417 (N_8417,N_6431,N_7449);
or U8418 (N_8418,N_6664,N_6879);
nand U8419 (N_8419,N_6047,N_6131);
and U8420 (N_8420,N_6468,N_6445);
xor U8421 (N_8421,N_6704,N_7143);
xnor U8422 (N_8422,N_6217,N_6883);
and U8423 (N_8423,N_6633,N_6258);
and U8424 (N_8424,N_7197,N_6947);
nor U8425 (N_8425,N_6985,N_6571);
xnor U8426 (N_8426,N_6113,N_6315);
nand U8427 (N_8427,N_7448,N_7352);
nor U8428 (N_8428,N_6331,N_6615);
xor U8429 (N_8429,N_7191,N_7310);
and U8430 (N_8430,N_6253,N_6374);
nor U8431 (N_8431,N_7012,N_7262);
or U8432 (N_8432,N_6960,N_6206);
nand U8433 (N_8433,N_6650,N_6497);
nor U8434 (N_8434,N_6486,N_6032);
nand U8435 (N_8435,N_6414,N_7052);
nor U8436 (N_8436,N_6820,N_6223);
and U8437 (N_8437,N_6613,N_7352);
or U8438 (N_8438,N_6396,N_6088);
or U8439 (N_8439,N_6145,N_6092);
or U8440 (N_8440,N_6698,N_6890);
and U8441 (N_8441,N_6084,N_6590);
and U8442 (N_8442,N_7014,N_6884);
nor U8443 (N_8443,N_6784,N_7097);
nand U8444 (N_8444,N_6052,N_6605);
nand U8445 (N_8445,N_6584,N_7100);
nand U8446 (N_8446,N_7036,N_6985);
or U8447 (N_8447,N_6461,N_6267);
nor U8448 (N_8448,N_7312,N_7499);
or U8449 (N_8449,N_6641,N_6447);
nand U8450 (N_8450,N_6084,N_6952);
nor U8451 (N_8451,N_6584,N_7382);
nor U8452 (N_8452,N_6569,N_6003);
or U8453 (N_8453,N_6920,N_6340);
and U8454 (N_8454,N_6801,N_6451);
nand U8455 (N_8455,N_6695,N_6897);
nor U8456 (N_8456,N_6183,N_6178);
xnor U8457 (N_8457,N_6560,N_6416);
and U8458 (N_8458,N_6443,N_6668);
or U8459 (N_8459,N_6500,N_7322);
or U8460 (N_8460,N_7071,N_6852);
xor U8461 (N_8461,N_7131,N_6870);
nor U8462 (N_8462,N_6714,N_7018);
xor U8463 (N_8463,N_6318,N_7206);
nand U8464 (N_8464,N_7164,N_6865);
xnor U8465 (N_8465,N_7044,N_6939);
and U8466 (N_8466,N_6269,N_7071);
nand U8467 (N_8467,N_6652,N_6544);
nor U8468 (N_8468,N_6306,N_6365);
xnor U8469 (N_8469,N_6507,N_7123);
or U8470 (N_8470,N_6273,N_6739);
nor U8471 (N_8471,N_7102,N_6479);
xnor U8472 (N_8472,N_6867,N_7339);
xnor U8473 (N_8473,N_6371,N_6790);
or U8474 (N_8474,N_7054,N_7357);
xor U8475 (N_8475,N_6833,N_6301);
and U8476 (N_8476,N_6735,N_6082);
nor U8477 (N_8477,N_7199,N_6598);
nor U8478 (N_8478,N_7138,N_6160);
nand U8479 (N_8479,N_6976,N_7036);
and U8480 (N_8480,N_6855,N_6917);
nand U8481 (N_8481,N_6288,N_6906);
xor U8482 (N_8482,N_6817,N_6100);
nor U8483 (N_8483,N_6901,N_6385);
xnor U8484 (N_8484,N_7314,N_6561);
or U8485 (N_8485,N_7300,N_6420);
xor U8486 (N_8486,N_6778,N_6269);
nand U8487 (N_8487,N_7274,N_6698);
nor U8488 (N_8488,N_6256,N_7288);
or U8489 (N_8489,N_7323,N_7276);
xor U8490 (N_8490,N_6101,N_6188);
nand U8491 (N_8491,N_6034,N_6331);
or U8492 (N_8492,N_7310,N_7388);
nand U8493 (N_8493,N_7199,N_7489);
or U8494 (N_8494,N_7054,N_6478);
and U8495 (N_8495,N_7455,N_6686);
nor U8496 (N_8496,N_6270,N_6224);
or U8497 (N_8497,N_6352,N_7444);
xor U8498 (N_8498,N_6958,N_6668);
or U8499 (N_8499,N_6327,N_6450);
xnor U8500 (N_8500,N_6802,N_6550);
or U8501 (N_8501,N_7303,N_6279);
and U8502 (N_8502,N_7240,N_6077);
xnor U8503 (N_8503,N_6334,N_6016);
nor U8504 (N_8504,N_6168,N_6182);
and U8505 (N_8505,N_6749,N_6532);
or U8506 (N_8506,N_6279,N_7002);
nor U8507 (N_8507,N_6567,N_7023);
or U8508 (N_8508,N_6751,N_6701);
nor U8509 (N_8509,N_6907,N_6004);
nor U8510 (N_8510,N_6252,N_7186);
or U8511 (N_8511,N_7037,N_6692);
nor U8512 (N_8512,N_6042,N_6391);
xor U8513 (N_8513,N_7009,N_6739);
and U8514 (N_8514,N_6316,N_6055);
and U8515 (N_8515,N_6179,N_6208);
or U8516 (N_8516,N_7068,N_6243);
and U8517 (N_8517,N_6539,N_7173);
nor U8518 (N_8518,N_7153,N_6592);
nand U8519 (N_8519,N_6350,N_6723);
nor U8520 (N_8520,N_6031,N_6991);
nor U8521 (N_8521,N_7211,N_6448);
xnor U8522 (N_8522,N_6501,N_6788);
xnor U8523 (N_8523,N_7403,N_7434);
nor U8524 (N_8524,N_6818,N_6796);
or U8525 (N_8525,N_6688,N_6500);
or U8526 (N_8526,N_6473,N_7422);
nor U8527 (N_8527,N_7376,N_6366);
xnor U8528 (N_8528,N_7443,N_7110);
or U8529 (N_8529,N_6458,N_7422);
and U8530 (N_8530,N_6885,N_6728);
nand U8531 (N_8531,N_6318,N_6349);
xor U8532 (N_8532,N_6250,N_6075);
nand U8533 (N_8533,N_7132,N_7167);
nor U8534 (N_8534,N_7088,N_6930);
nand U8535 (N_8535,N_6365,N_7277);
and U8536 (N_8536,N_7108,N_6283);
or U8537 (N_8537,N_6986,N_6778);
or U8538 (N_8538,N_6386,N_7108);
nand U8539 (N_8539,N_6581,N_6316);
and U8540 (N_8540,N_7240,N_7409);
or U8541 (N_8541,N_7121,N_6486);
nand U8542 (N_8542,N_6307,N_6864);
or U8543 (N_8543,N_7423,N_6063);
nand U8544 (N_8544,N_6644,N_7294);
nor U8545 (N_8545,N_6441,N_6477);
nor U8546 (N_8546,N_7232,N_7382);
and U8547 (N_8547,N_6582,N_6885);
and U8548 (N_8548,N_7443,N_6060);
and U8549 (N_8549,N_6920,N_6942);
xnor U8550 (N_8550,N_6848,N_6804);
nor U8551 (N_8551,N_7417,N_6433);
or U8552 (N_8552,N_6385,N_7273);
xnor U8553 (N_8553,N_6885,N_7330);
nor U8554 (N_8554,N_6218,N_6717);
or U8555 (N_8555,N_6719,N_7379);
and U8556 (N_8556,N_6884,N_7369);
and U8557 (N_8557,N_7124,N_6026);
or U8558 (N_8558,N_6960,N_6898);
or U8559 (N_8559,N_6286,N_6245);
xnor U8560 (N_8560,N_6309,N_7250);
or U8561 (N_8561,N_6219,N_7082);
nand U8562 (N_8562,N_6066,N_6832);
or U8563 (N_8563,N_7115,N_7432);
nand U8564 (N_8564,N_7099,N_7113);
nand U8565 (N_8565,N_7064,N_7002);
or U8566 (N_8566,N_6527,N_6894);
or U8567 (N_8567,N_6195,N_6816);
nor U8568 (N_8568,N_7409,N_6624);
xor U8569 (N_8569,N_7393,N_6256);
and U8570 (N_8570,N_6884,N_6802);
nor U8571 (N_8571,N_6661,N_6863);
and U8572 (N_8572,N_6627,N_6803);
or U8573 (N_8573,N_7027,N_6425);
nor U8574 (N_8574,N_6040,N_7377);
nand U8575 (N_8575,N_6985,N_6453);
and U8576 (N_8576,N_7222,N_7494);
xor U8577 (N_8577,N_7034,N_6714);
xor U8578 (N_8578,N_7432,N_6000);
nand U8579 (N_8579,N_6428,N_7290);
or U8580 (N_8580,N_7080,N_7173);
xor U8581 (N_8581,N_6052,N_7414);
and U8582 (N_8582,N_6901,N_6211);
xor U8583 (N_8583,N_6903,N_6493);
xor U8584 (N_8584,N_6809,N_7307);
nor U8585 (N_8585,N_7439,N_7017);
xnor U8586 (N_8586,N_6374,N_6757);
nor U8587 (N_8587,N_6372,N_7344);
xnor U8588 (N_8588,N_6487,N_7308);
nor U8589 (N_8589,N_6964,N_7186);
xor U8590 (N_8590,N_6853,N_6151);
nand U8591 (N_8591,N_6011,N_6022);
nand U8592 (N_8592,N_7034,N_7091);
nor U8593 (N_8593,N_7394,N_7148);
and U8594 (N_8594,N_6892,N_6343);
xor U8595 (N_8595,N_6903,N_7474);
xnor U8596 (N_8596,N_6721,N_6327);
or U8597 (N_8597,N_6127,N_7302);
xnor U8598 (N_8598,N_6963,N_6546);
nor U8599 (N_8599,N_7159,N_7448);
or U8600 (N_8600,N_6395,N_6164);
or U8601 (N_8601,N_7117,N_7392);
or U8602 (N_8602,N_7134,N_6069);
xor U8603 (N_8603,N_6913,N_6026);
or U8604 (N_8604,N_7232,N_6655);
nand U8605 (N_8605,N_6045,N_7136);
and U8606 (N_8606,N_6537,N_6996);
xnor U8607 (N_8607,N_7427,N_6339);
and U8608 (N_8608,N_6993,N_6624);
nand U8609 (N_8609,N_6071,N_7244);
xnor U8610 (N_8610,N_6648,N_6820);
xnor U8611 (N_8611,N_7375,N_6288);
xnor U8612 (N_8612,N_6471,N_6105);
nand U8613 (N_8613,N_7202,N_6339);
nor U8614 (N_8614,N_6027,N_7021);
and U8615 (N_8615,N_7282,N_6273);
or U8616 (N_8616,N_7393,N_6131);
xor U8617 (N_8617,N_6296,N_7007);
nand U8618 (N_8618,N_7235,N_6229);
nand U8619 (N_8619,N_6533,N_6332);
or U8620 (N_8620,N_7444,N_6407);
or U8621 (N_8621,N_7340,N_7332);
or U8622 (N_8622,N_6524,N_6061);
nand U8623 (N_8623,N_6753,N_7156);
nand U8624 (N_8624,N_6164,N_6373);
or U8625 (N_8625,N_7393,N_7001);
and U8626 (N_8626,N_6981,N_6297);
nand U8627 (N_8627,N_6990,N_6518);
xnor U8628 (N_8628,N_6245,N_6722);
or U8629 (N_8629,N_6235,N_6123);
or U8630 (N_8630,N_6251,N_6264);
nor U8631 (N_8631,N_6865,N_6810);
nor U8632 (N_8632,N_6051,N_7130);
or U8633 (N_8633,N_6792,N_6294);
xnor U8634 (N_8634,N_6267,N_6171);
nor U8635 (N_8635,N_6674,N_6414);
and U8636 (N_8636,N_6089,N_7248);
nor U8637 (N_8637,N_7435,N_6775);
or U8638 (N_8638,N_6874,N_6316);
nor U8639 (N_8639,N_7421,N_7164);
nand U8640 (N_8640,N_6920,N_6957);
and U8641 (N_8641,N_6190,N_6845);
nor U8642 (N_8642,N_6101,N_6897);
and U8643 (N_8643,N_6253,N_6492);
or U8644 (N_8644,N_6969,N_7012);
xnor U8645 (N_8645,N_7078,N_7263);
nor U8646 (N_8646,N_6754,N_6160);
nand U8647 (N_8647,N_6494,N_6548);
xor U8648 (N_8648,N_6682,N_6931);
and U8649 (N_8649,N_7495,N_6754);
nor U8650 (N_8650,N_6578,N_6171);
and U8651 (N_8651,N_6168,N_7065);
and U8652 (N_8652,N_6648,N_7339);
and U8653 (N_8653,N_6825,N_7189);
nor U8654 (N_8654,N_6680,N_6776);
nor U8655 (N_8655,N_7226,N_7371);
nand U8656 (N_8656,N_7475,N_6351);
nor U8657 (N_8657,N_7477,N_6887);
nor U8658 (N_8658,N_7256,N_7315);
nand U8659 (N_8659,N_6865,N_6122);
and U8660 (N_8660,N_7197,N_7467);
nand U8661 (N_8661,N_6369,N_6589);
or U8662 (N_8662,N_7042,N_6361);
or U8663 (N_8663,N_6034,N_7037);
and U8664 (N_8664,N_6726,N_7334);
nand U8665 (N_8665,N_7085,N_6040);
nand U8666 (N_8666,N_6410,N_6531);
and U8667 (N_8667,N_6227,N_7117);
xnor U8668 (N_8668,N_6597,N_6733);
nor U8669 (N_8669,N_6352,N_6936);
and U8670 (N_8670,N_6605,N_7289);
and U8671 (N_8671,N_7080,N_6244);
xor U8672 (N_8672,N_6290,N_6121);
and U8673 (N_8673,N_6643,N_6385);
and U8674 (N_8674,N_6146,N_6242);
or U8675 (N_8675,N_6795,N_7463);
and U8676 (N_8676,N_7373,N_7104);
xor U8677 (N_8677,N_7465,N_6475);
nor U8678 (N_8678,N_7163,N_6760);
or U8679 (N_8679,N_6882,N_6616);
nand U8680 (N_8680,N_6307,N_6093);
or U8681 (N_8681,N_6937,N_6073);
and U8682 (N_8682,N_6435,N_7272);
nor U8683 (N_8683,N_6409,N_6248);
xor U8684 (N_8684,N_7419,N_6891);
and U8685 (N_8685,N_7041,N_7259);
xnor U8686 (N_8686,N_6207,N_6953);
xor U8687 (N_8687,N_7331,N_6973);
and U8688 (N_8688,N_6148,N_7116);
nor U8689 (N_8689,N_6140,N_6391);
nor U8690 (N_8690,N_7177,N_6773);
nand U8691 (N_8691,N_6992,N_6317);
xnor U8692 (N_8692,N_7437,N_6014);
nand U8693 (N_8693,N_6407,N_6351);
or U8694 (N_8694,N_7320,N_6572);
xnor U8695 (N_8695,N_7038,N_6713);
and U8696 (N_8696,N_7356,N_7069);
or U8697 (N_8697,N_7153,N_6413);
xor U8698 (N_8698,N_6460,N_7293);
nor U8699 (N_8699,N_7036,N_7265);
and U8700 (N_8700,N_7238,N_7027);
xor U8701 (N_8701,N_7024,N_7463);
or U8702 (N_8702,N_7020,N_6959);
or U8703 (N_8703,N_6874,N_6824);
nand U8704 (N_8704,N_6291,N_7193);
or U8705 (N_8705,N_6913,N_7457);
or U8706 (N_8706,N_6441,N_6513);
xor U8707 (N_8707,N_7179,N_7284);
and U8708 (N_8708,N_6571,N_6542);
nor U8709 (N_8709,N_6508,N_7015);
nor U8710 (N_8710,N_6932,N_6984);
nand U8711 (N_8711,N_6683,N_7080);
or U8712 (N_8712,N_6887,N_6609);
nor U8713 (N_8713,N_6486,N_7090);
nand U8714 (N_8714,N_6269,N_6278);
and U8715 (N_8715,N_6185,N_6214);
and U8716 (N_8716,N_6458,N_6875);
or U8717 (N_8717,N_6763,N_7279);
xor U8718 (N_8718,N_7302,N_6693);
nor U8719 (N_8719,N_7499,N_6548);
or U8720 (N_8720,N_6904,N_7242);
and U8721 (N_8721,N_7078,N_6200);
nand U8722 (N_8722,N_6218,N_6304);
nand U8723 (N_8723,N_6036,N_6368);
nor U8724 (N_8724,N_6424,N_6338);
xnor U8725 (N_8725,N_7130,N_6458);
nand U8726 (N_8726,N_6108,N_7183);
xor U8727 (N_8727,N_6211,N_6380);
and U8728 (N_8728,N_7456,N_6334);
nor U8729 (N_8729,N_6471,N_6541);
nor U8730 (N_8730,N_7180,N_7483);
nand U8731 (N_8731,N_6740,N_6791);
or U8732 (N_8732,N_6542,N_6739);
nand U8733 (N_8733,N_7198,N_6342);
or U8734 (N_8734,N_6259,N_7355);
nor U8735 (N_8735,N_6399,N_6077);
and U8736 (N_8736,N_7258,N_6561);
nor U8737 (N_8737,N_6735,N_6262);
and U8738 (N_8738,N_7197,N_6734);
nand U8739 (N_8739,N_6810,N_6365);
nand U8740 (N_8740,N_6698,N_7389);
nor U8741 (N_8741,N_6433,N_6372);
nor U8742 (N_8742,N_6124,N_7148);
xnor U8743 (N_8743,N_6292,N_6506);
nor U8744 (N_8744,N_7172,N_6110);
xnor U8745 (N_8745,N_6673,N_7477);
and U8746 (N_8746,N_7485,N_6282);
nand U8747 (N_8747,N_7477,N_6311);
and U8748 (N_8748,N_6250,N_6172);
xor U8749 (N_8749,N_7056,N_6836);
or U8750 (N_8750,N_7281,N_6058);
or U8751 (N_8751,N_6540,N_7249);
nor U8752 (N_8752,N_6758,N_6392);
or U8753 (N_8753,N_6820,N_6285);
or U8754 (N_8754,N_6895,N_6660);
xor U8755 (N_8755,N_7019,N_6311);
or U8756 (N_8756,N_6831,N_7205);
nand U8757 (N_8757,N_7250,N_6773);
nor U8758 (N_8758,N_6407,N_6640);
nor U8759 (N_8759,N_7372,N_6220);
nor U8760 (N_8760,N_7192,N_6150);
or U8761 (N_8761,N_6552,N_6346);
nand U8762 (N_8762,N_6562,N_6265);
and U8763 (N_8763,N_6057,N_7200);
or U8764 (N_8764,N_6375,N_6971);
nor U8765 (N_8765,N_6202,N_6025);
and U8766 (N_8766,N_6525,N_7169);
or U8767 (N_8767,N_6131,N_6967);
and U8768 (N_8768,N_7462,N_6620);
xnor U8769 (N_8769,N_6740,N_7358);
or U8770 (N_8770,N_7364,N_7117);
xnor U8771 (N_8771,N_7203,N_6550);
nor U8772 (N_8772,N_7006,N_6897);
and U8773 (N_8773,N_6946,N_6876);
nor U8774 (N_8774,N_6707,N_6217);
nand U8775 (N_8775,N_7110,N_6828);
nor U8776 (N_8776,N_7140,N_6061);
nor U8777 (N_8777,N_7149,N_6644);
nor U8778 (N_8778,N_7139,N_7212);
or U8779 (N_8779,N_6893,N_6874);
nor U8780 (N_8780,N_6480,N_6377);
or U8781 (N_8781,N_7085,N_6083);
or U8782 (N_8782,N_6227,N_7270);
nor U8783 (N_8783,N_6062,N_6179);
xor U8784 (N_8784,N_6956,N_7319);
or U8785 (N_8785,N_7476,N_6089);
nand U8786 (N_8786,N_6971,N_6625);
or U8787 (N_8787,N_6420,N_6382);
or U8788 (N_8788,N_6773,N_6258);
nand U8789 (N_8789,N_6039,N_6931);
or U8790 (N_8790,N_6104,N_7072);
nor U8791 (N_8791,N_7408,N_6044);
nand U8792 (N_8792,N_7105,N_6811);
or U8793 (N_8793,N_7037,N_7283);
and U8794 (N_8794,N_7043,N_6548);
or U8795 (N_8795,N_6311,N_6508);
nor U8796 (N_8796,N_6782,N_7013);
nor U8797 (N_8797,N_6043,N_7446);
or U8798 (N_8798,N_6775,N_6525);
nor U8799 (N_8799,N_7185,N_6016);
and U8800 (N_8800,N_7177,N_7041);
xor U8801 (N_8801,N_6428,N_6698);
xnor U8802 (N_8802,N_6611,N_7037);
xor U8803 (N_8803,N_6848,N_6971);
xor U8804 (N_8804,N_6605,N_7309);
nand U8805 (N_8805,N_6379,N_7469);
or U8806 (N_8806,N_6221,N_6112);
nor U8807 (N_8807,N_7412,N_6560);
or U8808 (N_8808,N_7218,N_6614);
xnor U8809 (N_8809,N_6816,N_6695);
nand U8810 (N_8810,N_6289,N_6310);
and U8811 (N_8811,N_6382,N_6198);
xnor U8812 (N_8812,N_6409,N_6508);
and U8813 (N_8813,N_7320,N_6438);
or U8814 (N_8814,N_6369,N_6240);
nand U8815 (N_8815,N_7158,N_7073);
nor U8816 (N_8816,N_6632,N_6925);
nor U8817 (N_8817,N_7498,N_6112);
nor U8818 (N_8818,N_7363,N_6434);
xnor U8819 (N_8819,N_6039,N_6918);
and U8820 (N_8820,N_6521,N_7289);
xnor U8821 (N_8821,N_7348,N_6618);
xor U8822 (N_8822,N_6711,N_6730);
and U8823 (N_8823,N_6390,N_6468);
xnor U8824 (N_8824,N_7113,N_6466);
and U8825 (N_8825,N_6201,N_6613);
nor U8826 (N_8826,N_6634,N_6516);
nor U8827 (N_8827,N_6810,N_6467);
or U8828 (N_8828,N_6094,N_6599);
nand U8829 (N_8829,N_6253,N_6934);
nor U8830 (N_8830,N_6143,N_6103);
nand U8831 (N_8831,N_7292,N_6832);
nand U8832 (N_8832,N_6432,N_6791);
nor U8833 (N_8833,N_6348,N_7074);
nand U8834 (N_8834,N_6877,N_6364);
nor U8835 (N_8835,N_6836,N_7479);
nor U8836 (N_8836,N_6972,N_7045);
xor U8837 (N_8837,N_6177,N_7111);
nor U8838 (N_8838,N_7407,N_6186);
xor U8839 (N_8839,N_6134,N_7003);
xor U8840 (N_8840,N_6852,N_7444);
nand U8841 (N_8841,N_7013,N_6700);
nand U8842 (N_8842,N_7399,N_7368);
or U8843 (N_8843,N_6635,N_7365);
or U8844 (N_8844,N_6898,N_7357);
and U8845 (N_8845,N_7070,N_7338);
or U8846 (N_8846,N_6861,N_7281);
or U8847 (N_8847,N_6904,N_6560);
nor U8848 (N_8848,N_7455,N_6501);
and U8849 (N_8849,N_7229,N_6189);
or U8850 (N_8850,N_7014,N_6406);
nor U8851 (N_8851,N_7196,N_6547);
nor U8852 (N_8852,N_6570,N_6377);
nor U8853 (N_8853,N_6077,N_6014);
xnor U8854 (N_8854,N_6843,N_7446);
and U8855 (N_8855,N_7345,N_7349);
and U8856 (N_8856,N_6218,N_6469);
or U8857 (N_8857,N_6783,N_6986);
xnor U8858 (N_8858,N_6410,N_6310);
xor U8859 (N_8859,N_6630,N_7430);
and U8860 (N_8860,N_6644,N_7180);
nand U8861 (N_8861,N_6605,N_6776);
nand U8862 (N_8862,N_7400,N_6895);
and U8863 (N_8863,N_7364,N_6500);
or U8864 (N_8864,N_6559,N_6248);
and U8865 (N_8865,N_6563,N_7354);
or U8866 (N_8866,N_6469,N_6675);
nor U8867 (N_8867,N_7139,N_6259);
xor U8868 (N_8868,N_7472,N_6667);
nor U8869 (N_8869,N_6960,N_6430);
nand U8870 (N_8870,N_6158,N_7452);
and U8871 (N_8871,N_6284,N_6298);
xnor U8872 (N_8872,N_7299,N_7387);
and U8873 (N_8873,N_6163,N_6057);
and U8874 (N_8874,N_7308,N_6217);
xor U8875 (N_8875,N_6758,N_6480);
nor U8876 (N_8876,N_6792,N_6095);
and U8877 (N_8877,N_7281,N_6590);
nand U8878 (N_8878,N_6413,N_6036);
or U8879 (N_8879,N_6340,N_6126);
nand U8880 (N_8880,N_6017,N_6949);
nor U8881 (N_8881,N_6176,N_7160);
nor U8882 (N_8882,N_7057,N_6476);
xor U8883 (N_8883,N_6472,N_6536);
nand U8884 (N_8884,N_6107,N_6735);
and U8885 (N_8885,N_7295,N_7481);
xor U8886 (N_8886,N_6064,N_7161);
or U8887 (N_8887,N_6821,N_7129);
xor U8888 (N_8888,N_6631,N_6280);
and U8889 (N_8889,N_7039,N_6843);
and U8890 (N_8890,N_6755,N_6531);
nor U8891 (N_8891,N_6318,N_7111);
nand U8892 (N_8892,N_6306,N_6821);
nor U8893 (N_8893,N_6654,N_6077);
or U8894 (N_8894,N_6048,N_7166);
and U8895 (N_8895,N_6692,N_7042);
or U8896 (N_8896,N_6267,N_6071);
nor U8897 (N_8897,N_6585,N_6598);
and U8898 (N_8898,N_7163,N_7097);
and U8899 (N_8899,N_6209,N_6924);
nor U8900 (N_8900,N_6766,N_7066);
nand U8901 (N_8901,N_6662,N_6937);
and U8902 (N_8902,N_6738,N_6785);
nand U8903 (N_8903,N_6785,N_6633);
xor U8904 (N_8904,N_6569,N_6423);
or U8905 (N_8905,N_6502,N_6088);
nor U8906 (N_8906,N_7322,N_6443);
or U8907 (N_8907,N_6509,N_7117);
nand U8908 (N_8908,N_7475,N_6380);
nor U8909 (N_8909,N_7432,N_7031);
or U8910 (N_8910,N_6638,N_6087);
xor U8911 (N_8911,N_7208,N_6657);
or U8912 (N_8912,N_6207,N_6683);
nor U8913 (N_8913,N_6572,N_7125);
xor U8914 (N_8914,N_7289,N_6724);
and U8915 (N_8915,N_6425,N_6286);
and U8916 (N_8916,N_7246,N_6289);
or U8917 (N_8917,N_6886,N_6888);
and U8918 (N_8918,N_7048,N_6309);
xnor U8919 (N_8919,N_6337,N_6242);
nor U8920 (N_8920,N_6269,N_6466);
or U8921 (N_8921,N_6181,N_6094);
and U8922 (N_8922,N_7269,N_6701);
or U8923 (N_8923,N_6002,N_7433);
and U8924 (N_8924,N_6881,N_6606);
nand U8925 (N_8925,N_6352,N_6908);
nor U8926 (N_8926,N_6369,N_7173);
or U8927 (N_8927,N_7391,N_6187);
and U8928 (N_8928,N_6034,N_6057);
nand U8929 (N_8929,N_6538,N_6854);
or U8930 (N_8930,N_6820,N_6969);
nor U8931 (N_8931,N_7484,N_6352);
and U8932 (N_8932,N_6486,N_7159);
and U8933 (N_8933,N_7388,N_6158);
and U8934 (N_8934,N_6976,N_6470);
or U8935 (N_8935,N_6975,N_7320);
nor U8936 (N_8936,N_6944,N_6724);
nor U8937 (N_8937,N_7459,N_6517);
or U8938 (N_8938,N_7067,N_7152);
or U8939 (N_8939,N_6070,N_6124);
xnor U8940 (N_8940,N_6709,N_6073);
or U8941 (N_8941,N_7338,N_7415);
xnor U8942 (N_8942,N_6465,N_6029);
xnor U8943 (N_8943,N_7392,N_7425);
or U8944 (N_8944,N_6486,N_6800);
nor U8945 (N_8945,N_6475,N_6772);
nor U8946 (N_8946,N_7251,N_6763);
and U8947 (N_8947,N_6886,N_6042);
and U8948 (N_8948,N_7010,N_6075);
or U8949 (N_8949,N_7007,N_6476);
nand U8950 (N_8950,N_6414,N_7484);
nand U8951 (N_8951,N_6682,N_6824);
nand U8952 (N_8952,N_6458,N_7121);
nor U8953 (N_8953,N_7281,N_6716);
or U8954 (N_8954,N_6762,N_6429);
or U8955 (N_8955,N_7152,N_7462);
nor U8956 (N_8956,N_7193,N_6757);
and U8957 (N_8957,N_7144,N_7076);
and U8958 (N_8958,N_6035,N_6022);
nor U8959 (N_8959,N_7414,N_6213);
xor U8960 (N_8960,N_7145,N_7230);
or U8961 (N_8961,N_7151,N_7407);
nor U8962 (N_8962,N_7022,N_7014);
and U8963 (N_8963,N_7457,N_6312);
or U8964 (N_8964,N_7234,N_6283);
nand U8965 (N_8965,N_6405,N_6684);
xnor U8966 (N_8966,N_6060,N_6510);
xor U8967 (N_8967,N_6200,N_7111);
nor U8968 (N_8968,N_6453,N_6295);
nor U8969 (N_8969,N_7283,N_7095);
xnor U8970 (N_8970,N_6477,N_6118);
nand U8971 (N_8971,N_7058,N_7013);
or U8972 (N_8972,N_6352,N_6045);
nor U8973 (N_8973,N_7342,N_7389);
nor U8974 (N_8974,N_6325,N_6718);
nor U8975 (N_8975,N_6989,N_7333);
and U8976 (N_8976,N_6747,N_7004);
xnor U8977 (N_8977,N_7303,N_6121);
xnor U8978 (N_8978,N_7288,N_6241);
xor U8979 (N_8979,N_6352,N_6167);
nor U8980 (N_8980,N_7291,N_7195);
or U8981 (N_8981,N_6400,N_6737);
or U8982 (N_8982,N_6767,N_7346);
xnor U8983 (N_8983,N_7413,N_6411);
xnor U8984 (N_8984,N_7337,N_6341);
or U8985 (N_8985,N_6233,N_6620);
nor U8986 (N_8986,N_6067,N_6789);
or U8987 (N_8987,N_6658,N_6770);
and U8988 (N_8988,N_6501,N_6418);
and U8989 (N_8989,N_6177,N_7412);
xor U8990 (N_8990,N_6690,N_6467);
xnor U8991 (N_8991,N_6523,N_7291);
nand U8992 (N_8992,N_6574,N_7188);
nor U8993 (N_8993,N_7376,N_7289);
and U8994 (N_8994,N_6257,N_6710);
nand U8995 (N_8995,N_7302,N_7246);
xnor U8996 (N_8996,N_6743,N_6260);
nor U8997 (N_8997,N_6038,N_6753);
nor U8998 (N_8998,N_6422,N_7208);
nand U8999 (N_8999,N_7271,N_7494);
or U9000 (N_9000,N_7826,N_8490);
nand U9001 (N_9001,N_8123,N_8578);
nor U9002 (N_9002,N_8095,N_8685);
nor U9003 (N_9003,N_8950,N_8875);
xor U9004 (N_9004,N_8254,N_8883);
or U9005 (N_9005,N_7733,N_7551);
nor U9006 (N_9006,N_7856,N_8093);
and U9007 (N_9007,N_7608,N_7603);
nand U9008 (N_9008,N_7958,N_8345);
or U9009 (N_9009,N_8717,N_7898);
or U9010 (N_9010,N_7751,N_7609);
nor U9011 (N_9011,N_8487,N_7593);
xor U9012 (N_9012,N_8069,N_7872);
or U9013 (N_9013,N_8484,N_7730);
and U9014 (N_9014,N_8549,N_8369);
nand U9015 (N_9015,N_8473,N_7983);
nand U9016 (N_9016,N_8538,N_7818);
nand U9017 (N_9017,N_8469,N_8871);
or U9018 (N_9018,N_7746,N_7937);
xnor U9019 (N_9019,N_8702,N_8787);
nor U9020 (N_9020,N_8737,N_8138);
xor U9021 (N_9021,N_8979,N_7536);
or U9022 (N_9022,N_7743,N_7763);
nand U9023 (N_9023,N_8195,N_8042);
nand U9024 (N_9024,N_7945,N_8658);
nor U9025 (N_9025,N_8850,N_8418);
nand U9026 (N_9026,N_8651,N_8410);
and U9027 (N_9027,N_7654,N_8477);
nor U9028 (N_9028,N_8736,N_8684);
nand U9029 (N_9029,N_8809,N_8020);
or U9030 (N_9030,N_7615,N_7930);
xor U9031 (N_9031,N_8358,N_8947);
nand U9032 (N_9032,N_8072,N_8674);
and U9033 (N_9033,N_7601,N_8274);
nand U9034 (N_9034,N_7677,N_7700);
and U9035 (N_9035,N_7750,N_8184);
and U9036 (N_9036,N_8506,N_8117);
xor U9037 (N_9037,N_8091,N_8539);
xnor U9038 (N_9038,N_7893,N_8858);
nand U9039 (N_9039,N_8942,N_8156);
xnor U9040 (N_9040,N_8011,N_8185);
and U9041 (N_9041,N_8909,N_8232);
nand U9042 (N_9042,N_8509,N_8522);
and U9043 (N_9043,N_8854,N_7820);
nor U9044 (N_9044,N_8677,N_7765);
or U9045 (N_9045,N_8575,N_8159);
xor U9046 (N_9046,N_7690,N_7670);
and U9047 (N_9047,N_8040,N_8803);
or U9048 (N_9048,N_8439,N_8820);
xnor U9049 (N_9049,N_8552,N_7716);
nor U9050 (N_9050,N_8433,N_7920);
or U9051 (N_9051,N_7860,N_7592);
and U9052 (N_9052,N_8372,N_8328);
xor U9053 (N_9053,N_8944,N_8992);
or U9054 (N_9054,N_8000,N_7582);
and U9055 (N_9055,N_7767,N_8965);
nor U9056 (N_9056,N_8049,N_8720);
and U9057 (N_9057,N_7809,N_8083);
nand U9058 (N_9058,N_7869,N_8155);
nor U9059 (N_9059,N_8830,N_7735);
nand U9060 (N_9060,N_8876,N_7754);
and U9061 (N_9061,N_8388,N_8887);
nor U9062 (N_9062,N_7644,N_7620);
and U9063 (N_9063,N_7511,N_7600);
or U9064 (N_9064,N_8894,N_8294);
nor U9065 (N_9065,N_8526,N_8163);
and U9066 (N_9066,N_7580,N_7915);
and U9067 (N_9067,N_8716,N_7845);
and U9068 (N_9068,N_8395,N_7507);
nand U9069 (N_9069,N_8380,N_8259);
and U9070 (N_9070,N_7769,N_8943);
xnor U9071 (N_9071,N_7839,N_8569);
nor U9072 (N_9072,N_8905,N_7571);
nand U9073 (N_9073,N_8529,N_8161);
nor U9074 (N_9074,N_7969,N_7939);
nand U9075 (N_9075,N_7914,N_7770);
and U9076 (N_9076,N_7828,N_7594);
nor U9077 (N_9077,N_8305,N_7715);
nor U9078 (N_9078,N_8951,N_8107);
xor U9079 (N_9079,N_7653,N_8620);
nor U9080 (N_9080,N_8900,N_8461);
nand U9081 (N_9081,N_7755,N_8488);
and U9082 (N_9082,N_7506,N_8081);
xnor U9083 (N_9083,N_7543,N_8260);
nor U9084 (N_9084,N_8551,N_7995);
or U9085 (N_9085,N_7556,N_8622);
nor U9086 (N_9086,N_8532,N_8707);
nand U9087 (N_9087,N_7907,N_7585);
nand U9088 (N_9088,N_8176,N_8839);
nor U9089 (N_9089,N_8841,N_8981);
and U9090 (N_9090,N_8193,N_7963);
nand U9091 (N_9091,N_8590,N_8730);
and U9092 (N_9092,N_8505,N_8705);
nand U9093 (N_9093,N_7738,N_7954);
and U9094 (N_9094,N_8394,N_8659);
or U9095 (N_9095,N_8443,N_8520);
xor U9096 (N_9096,N_8824,N_8472);
nor U9097 (N_9097,N_8675,N_8719);
xnor U9098 (N_9098,N_8917,N_7897);
nand U9099 (N_9099,N_7621,N_8481);
nor U9100 (N_9100,N_8082,N_8157);
nor U9101 (N_9101,N_7870,N_7502);
nor U9102 (N_9102,N_8728,N_8941);
nand U9103 (N_9103,N_7564,N_8791);
xnor U9104 (N_9104,N_8419,N_8631);
xnor U9105 (N_9105,N_7970,N_8363);
xnor U9106 (N_9106,N_7989,N_7921);
or U9107 (N_9107,N_8657,N_8312);
xor U9108 (N_9108,N_7524,N_8370);
xnor U9109 (N_9109,N_7866,N_8119);
or U9110 (N_9110,N_7520,N_7988);
or U9111 (N_9111,N_8321,N_8226);
or U9112 (N_9112,N_7799,N_8094);
nor U9113 (N_9113,N_8351,N_7581);
and U9114 (N_9114,N_8166,N_8792);
and U9115 (N_9115,N_8374,N_8017);
and U9116 (N_9116,N_8591,N_8057);
xor U9117 (N_9117,N_7817,N_7948);
xor U9118 (N_9118,N_8493,N_7798);
and U9119 (N_9119,N_7783,N_8945);
nand U9120 (N_9120,N_7778,N_7998);
xnor U9121 (N_9121,N_8101,N_8513);
nor U9122 (N_9122,N_7660,N_8669);
or U9123 (N_9123,N_7679,N_8234);
nand U9124 (N_9124,N_7774,N_7598);
nor U9125 (N_9125,N_7786,N_7731);
or U9126 (N_9126,N_8405,N_7924);
nand U9127 (N_9127,N_8279,N_7708);
xor U9128 (N_9128,N_7905,N_8152);
nor U9129 (N_9129,N_8576,N_8333);
nor U9130 (N_9130,N_7853,N_7957);
and U9131 (N_9131,N_8001,N_8554);
and U9132 (N_9132,N_7749,N_8113);
nor U9133 (N_9133,N_8571,N_7931);
or U9134 (N_9134,N_8486,N_7933);
nand U9135 (N_9135,N_8914,N_8149);
nand U9136 (N_9136,N_8540,N_8849);
and U9137 (N_9137,N_8390,N_7829);
or U9138 (N_9138,N_8832,N_8376);
nand U9139 (N_9139,N_8557,N_7583);
nor U9140 (N_9140,N_8186,N_8012);
nand U9141 (N_9141,N_8662,N_8106);
and U9142 (N_9142,N_8136,N_8938);
nor U9143 (N_9143,N_8062,N_8823);
nor U9144 (N_9144,N_8111,N_8521);
or U9145 (N_9145,N_7617,N_8187);
nor U9146 (N_9146,N_8811,N_8437);
nor U9147 (N_9147,N_7908,N_7978);
nor U9148 (N_9148,N_7952,N_7868);
xnor U9149 (N_9149,N_8097,N_8033);
and U9150 (N_9150,N_7579,N_8580);
xor U9151 (N_9151,N_8758,N_8969);
or U9152 (N_9152,N_8676,N_8930);
xnor U9153 (N_9153,N_8325,N_7628);
xnor U9154 (N_9154,N_7577,N_7500);
nor U9155 (N_9155,N_8398,N_8055);
nor U9156 (N_9156,N_8897,N_8976);
nor U9157 (N_9157,N_8112,N_8845);
xor U9158 (N_9158,N_8794,N_8212);
nor U9159 (N_9159,N_7588,N_8079);
nand U9160 (N_9160,N_8844,N_7960);
nand U9161 (N_9161,N_8046,N_7973);
nor U9162 (N_9162,N_7666,N_8137);
or U9163 (N_9163,N_8005,N_8162);
nand U9164 (N_9164,N_8180,N_8236);
nand U9165 (N_9165,N_8337,N_7505);
nor U9166 (N_9166,N_7855,N_7640);
nor U9167 (N_9167,N_8006,N_7525);
nor U9168 (N_9168,N_8699,N_8902);
xnor U9169 (N_9169,N_8627,N_8851);
and U9170 (N_9170,N_8073,N_8392);
and U9171 (N_9171,N_8668,N_8864);
nor U9172 (N_9172,N_8585,N_7668);
xnor U9173 (N_9173,N_8089,N_8542);
nor U9174 (N_9174,N_7667,N_8629);
or U9175 (N_9175,N_8868,N_8335);
nor U9176 (N_9176,N_8063,N_8170);
or U9177 (N_9177,N_8956,N_8643);
nor U9178 (N_9178,N_8070,N_8242);
or U9179 (N_9179,N_7964,N_7806);
xor U9180 (N_9180,N_8035,N_7521);
nand U9181 (N_9181,N_8299,N_8462);
and U9182 (N_9182,N_8881,N_8760);
and U9183 (N_9183,N_8805,N_8182);
nand U9184 (N_9184,N_8174,N_8588);
and U9185 (N_9185,N_7547,N_8141);
xor U9186 (N_9186,N_8822,N_7916);
xnor U9187 (N_9187,N_8199,N_7650);
or U9188 (N_9188,N_7890,N_8021);
nor U9189 (N_9189,N_8603,N_8708);
xor U9190 (N_9190,N_7707,N_7675);
and U9191 (N_9191,N_8387,N_8691);
nor U9192 (N_9192,N_7852,N_8188);
and U9193 (N_9193,N_8227,N_8744);
nand U9194 (N_9194,N_8755,N_8565);
and U9195 (N_9195,N_8338,N_7985);
xor U9196 (N_9196,N_8013,N_7711);
and U9197 (N_9197,N_8034,N_8907);
nand U9198 (N_9198,N_7761,N_8025);
nand U9199 (N_9199,N_8840,N_8039);
nor U9200 (N_9200,N_8019,N_8467);
nor U9201 (N_9201,N_7814,N_8371);
and U9202 (N_9202,N_8808,N_8617);
xor U9203 (N_9203,N_8504,N_7607);
or U9204 (N_9204,N_8454,N_8067);
or U9205 (N_9205,N_8334,N_8752);
and U9206 (N_9206,N_8289,N_8987);
nor U9207 (N_9207,N_7512,N_7833);
nor U9208 (N_9208,N_8596,N_8587);
nand U9209 (N_9209,N_8795,N_7944);
and U9210 (N_9210,N_7764,N_8826);
and U9211 (N_9211,N_7563,N_8561);
or U9212 (N_9212,N_8377,N_8389);
nor U9213 (N_9213,N_8124,N_8931);
or U9214 (N_9214,N_7655,N_8804);
nor U9215 (N_9215,N_8634,N_8712);
and U9216 (N_9216,N_7631,N_8923);
xor U9217 (N_9217,N_7982,N_7835);
and U9218 (N_9218,N_7724,N_8044);
nand U9219 (N_9219,N_7979,N_8625);
xnor U9220 (N_9220,N_8302,N_8225);
nand U9221 (N_9221,N_8228,N_7606);
nand U9222 (N_9222,N_8489,N_7501);
nand U9223 (N_9223,N_8807,N_7981);
or U9224 (N_9224,N_8679,N_8511);
nor U9225 (N_9225,N_7927,N_7542);
and U9226 (N_9226,N_8446,N_7947);
and U9227 (N_9227,N_8562,N_8441);
nand U9228 (N_9228,N_8635,N_8224);
and U9229 (N_9229,N_8798,N_8862);
or U9230 (N_9230,N_8422,N_8748);
xnor U9231 (N_9231,N_7534,N_8474);
nor U9232 (N_9232,N_8445,N_8349);
and U9233 (N_9233,N_8925,N_8975);
and U9234 (N_9234,N_8284,N_8815);
nor U9235 (N_9235,N_8604,N_8496);
or U9236 (N_9236,N_8507,N_8219);
or U9237 (N_9237,N_7721,N_8264);
or U9238 (N_9238,N_8191,N_8593);
and U9239 (N_9239,N_8074,N_8366);
nor U9240 (N_9240,N_8121,N_8451);
nand U9241 (N_9241,N_7759,N_8480);
nor U9242 (N_9242,N_7587,N_8753);
xor U9243 (N_9243,N_8403,N_8316);
nand U9244 (N_9244,N_8301,N_8940);
nand U9245 (N_9245,N_7732,N_7691);
xnor U9246 (N_9246,N_8636,N_8837);
nor U9247 (N_9247,N_8517,N_7742);
xor U9248 (N_9248,N_7794,N_8500);
nor U9249 (N_9249,N_7688,N_8041);
xor U9250 (N_9250,N_8353,N_8910);
xnor U9251 (N_9251,N_7923,N_8711);
xor U9252 (N_9252,N_8501,N_7885);
or U9253 (N_9253,N_8383,N_8038);
and U9254 (N_9254,N_7950,N_7889);
and U9255 (N_9255,N_8597,N_7535);
or U9256 (N_9256,N_8205,N_8856);
and U9257 (N_9257,N_8379,N_7837);
and U9258 (N_9258,N_8829,N_8782);
xor U9259 (N_9259,N_7632,N_8973);
nand U9260 (N_9260,N_7863,N_8273);
nand U9261 (N_9261,N_7823,N_8416);
nand U9262 (N_9262,N_8911,N_8528);
or U9263 (N_9263,N_8692,N_7902);
nor U9264 (N_9264,N_7857,N_8978);
nand U9265 (N_9265,N_8698,N_8512);
xor U9266 (N_9266,N_8269,N_7574);
nand U9267 (N_9267,N_8994,N_7762);
xor U9268 (N_9268,N_7651,N_8548);
xor U9269 (N_9269,N_8381,N_8560);
xor U9270 (N_9270,N_7793,N_8298);
or U9271 (N_9271,N_8204,N_8029);
nor U9272 (N_9272,N_8615,N_8471);
or U9273 (N_9273,N_8495,N_7848);
or U9274 (N_9274,N_8424,N_8757);
and U9275 (N_9275,N_8955,N_8458);
nor U9276 (N_9276,N_8601,N_8003);
and U9277 (N_9277,N_8014,N_8015);
nor U9278 (N_9278,N_8139,N_8314);
and U9279 (N_9279,N_8425,N_7727);
xor U9280 (N_9280,N_8645,N_7530);
nand U9281 (N_9281,N_8527,N_7619);
and U9282 (N_9282,N_8666,N_7768);
or U9283 (N_9283,N_8646,N_8638);
and U9284 (N_9284,N_7911,N_7858);
nand U9285 (N_9285,N_7672,N_8385);
and U9286 (N_9286,N_8774,N_8330);
nand U9287 (N_9287,N_8754,N_8741);
and U9288 (N_9288,N_7781,N_8595);
or U9289 (N_9289,N_8202,N_8890);
nand U9290 (N_9290,N_7725,N_8828);
nor U9291 (N_9291,N_8056,N_8621);
or U9292 (N_9292,N_7503,N_8713);
xor U9293 (N_9293,N_8282,N_7613);
nand U9294 (N_9294,N_8026,N_8287);
xor U9295 (N_9295,N_7909,N_8350);
nand U9296 (N_9296,N_8196,N_8047);
xor U9297 (N_9297,N_8378,N_8663);
xor U9298 (N_9298,N_8594,N_8616);
and U9299 (N_9299,N_8088,N_8573);
nand U9300 (N_9300,N_7514,N_7896);
xor U9301 (N_9301,N_8268,N_8788);
nor U9302 (N_9302,N_8114,N_7661);
nand U9303 (N_9303,N_8746,N_7805);
or U9304 (N_9304,N_8086,N_8581);
or U9305 (N_9305,N_8414,N_7819);
and U9306 (N_9306,N_7552,N_7702);
or U9307 (N_9307,N_8415,N_8605);
or U9308 (N_9308,N_7936,N_8050);
nor U9309 (N_9309,N_8609,N_7996);
xnor U9310 (N_9310,N_8311,N_8671);
nor U9311 (N_9311,N_7673,N_8308);
nand U9312 (N_9312,N_8556,N_7610);
and U9313 (N_9313,N_7758,N_8696);
or U9314 (N_9314,N_8723,N_7629);
nand U9315 (N_9315,N_7698,N_7633);
xnor U9316 (N_9316,N_8098,N_8343);
and U9317 (N_9317,N_8555,N_8411);
nand U9318 (N_9318,N_7859,N_8818);
xor U9319 (N_9319,N_7748,N_8563);
nor U9320 (N_9320,N_7575,N_7737);
and U9321 (N_9321,N_7706,N_8599);
xor U9322 (N_9322,N_8535,N_8080);
xnor U9323 (N_9323,N_8409,N_7959);
nand U9324 (N_9324,N_7901,N_8749);
and U9325 (N_9325,N_8336,N_8990);
nor U9326 (N_9326,N_8656,N_8146);
nand U9327 (N_9327,N_7703,N_7830);
nor U9328 (N_9328,N_8924,N_8255);
xor U9329 (N_9329,N_8843,N_7519);
or U9330 (N_9330,N_8545,N_8886);
nor U9331 (N_9331,N_8650,N_7576);
nor U9332 (N_9332,N_8853,N_8457);
nor U9333 (N_9333,N_7941,N_8970);
xor U9334 (N_9334,N_7807,N_8611);
nand U9335 (N_9335,N_7573,N_7987);
or U9336 (N_9336,N_8215,N_7961);
nand U9337 (N_9337,N_8756,N_8879);
nand U9338 (N_9338,N_8172,N_7627);
nand U9339 (N_9339,N_8200,N_8168);
and U9340 (N_9340,N_8530,N_7821);
nand U9341 (N_9341,N_8048,N_8633);
or U9342 (N_9342,N_8968,N_8160);
and U9343 (N_9343,N_8244,N_8134);
xor U9344 (N_9344,N_8743,N_8678);
xnor U9345 (N_9345,N_8901,N_8100);
xnor U9346 (N_9346,N_7695,N_7728);
nand U9347 (N_9347,N_8893,N_8993);
and U9348 (N_9348,N_7599,N_7910);
and U9349 (N_9349,N_8427,N_7771);
and U9350 (N_9350,N_8444,N_8999);
or U9351 (N_9351,N_8251,N_8491);
nand U9352 (N_9352,N_8197,N_7790);
or U9353 (N_9353,N_8547,N_8610);
or U9354 (N_9354,N_7773,N_8860);
and U9355 (N_9355,N_7892,N_8290);
nand U9356 (N_9356,N_8092,N_7722);
nor U9357 (N_9357,N_7741,N_8008);
xor U9358 (N_9358,N_8320,N_7584);
and U9359 (N_9359,N_8173,N_8885);
or U9360 (N_9360,N_7740,N_7906);
xnor U9361 (N_9361,N_7810,N_7934);
or U9362 (N_9362,N_7815,N_7928);
xnor U9363 (N_9363,N_8476,N_8948);
xnor U9364 (N_9364,N_7962,N_8252);
nand U9365 (N_9365,N_7878,N_7772);
xor U9366 (N_9366,N_7638,N_8253);
nand U9367 (N_9367,N_8751,N_7879);
xnor U9368 (N_9368,N_7867,N_8838);
nand U9369 (N_9369,N_8525,N_8102);
xor U9370 (N_9370,N_8078,N_7699);
or U9371 (N_9371,N_8877,N_8396);
nor U9372 (N_9372,N_8846,N_8776);
nand U9373 (N_9373,N_8296,N_8553);
and U9374 (N_9374,N_7834,N_7518);
nand U9375 (N_9375,N_8291,N_8884);
nor U9376 (N_9376,N_7623,N_8644);
xor U9377 (N_9377,N_8060,N_7625);
nand U9378 (N_9378,N_8384,N_7602);
xnor U9379 (N_9379,N_8733,N_8612);
nor U9380 (N_9380,N_8002,N_7747);
xor U9381 (N_9381,N_7801,N_8129);
nor U9382 (N_9382,N_8222,N_8690);
and U9383 (N_9383,N_7508,N_8614);
xor U9384 (N_9384,N_8402,N_8406);
and U9385 (N_9385,N_7782,N_8768);
or U9386 (N_9386,N_8151,N_7887);
nor U9387 (N_9387,N_8772,N_8304);
nand U9388 (N_9388,N_8245,N_8463);
or U9389 (N_9389,N_8145,N_8742);
and U9390 (N_9390,N_8324,N_8216);
or U9391 (N_9391,N_7545,N_8355);
nor U9392 (N_9392,N_8028,N_8283);
and U9393 (N_9393,N_8790,N_8649);
nor U9394 (N_9394,N_7657,N_8237);
nand U9395 (N_9395,N_7832,N_7803);
and U9396 (N_9396,N_7888,N_8865);
nand U9397 (N_9397,N_7663,N_7862);
nand U9398 (N_9398,N_8201,N_8797);
and U9399 (N_9399,N_7926,N_7674);
nor U9400 (N_9400,N_8010,N_7622);
or U9401 (N_9401,N_8217,N_8726);
nor U9402 (N_9402,N_8867,N_8831);
and U9403 (N_9403,N_8131,N_8432);
or U9404 (N_9404,N_8766,N_8206);
nor U9405 (N_9405,N_8103,N_8423);
and U9406 (N_9406,N_8066,N_7942);
xnor U9407 (N_9407,N_8420,N_8584);
xnor U9408 (N_9408,N_8574,N_8051);
and U9409 (N_9409,N_8275,N_7565);
or U9410 (N_9410,N_8550,N_7968);
or U9411 (N_9411,N_7986,N_8771);
xnor U9412 (N_9412,N_7656,N_7874);
or U9413 (N_9413,N_8814,N_7643);
xor U9414 (N_9414,N_7684,N_8936);
xnor U9415 (N_9415,N_8863,N_8916);
or U9416 (N_9416,N_8391,N_7560);
nand U9417 (N_9417,N_8703,N_8531);
xnor U9418 (N_9418,N_7766,N_8208);
nor U9419 (N_9419,N_8786,N_7877);
or U9420 (N_9420,N_7999,N_8870);
or U9421 (N_9421,N_8436,N_7526);
and U9422 (N_9422,N_7904,N_7692);
and U9423 (N_9423,N_8989,N_7554);
nor U9424 (N_9424,N_8655,N_8767);
and U9425 (N_9425,N_8963,N_7533);
nor U9426 (N_9426,N_8158,N_8670);
nor U9427 (N_9427,N_8265,N_7522);
nor U9428 (N_9428,N_8813,N_8440);
and U9429 (N_9429,N_8306,N_7591);
nor U9430 (N_9430,N_7558,N_8660);
xor U9431 (N_9431,N_7891,N_8519);
nor U9432 (N_9432,N_8125,N_8977);
nand U9433 (N_9433,N_8270,N_7949);
nand U9434 (N_9434,N_8018,N_8982);
nor U9435 (N_9435,N_8127,N_8721);
nor U9436 (N_9436,N_7553,N_8470);
nor U9437 (N_9437,N_8568,N_8855);
nand U9438 (N_9438,N_7517,N_8118);
or U9439 (N_9439,N_8896,N_8842);
xnor U9440 (N_9440,N_8309,N_8971);
and U9441 (N_9441,N_8583,N_8647);
or U9442 (N_9442,N_7729,N_8153);
or U9443 (N_9443,N_8919,N_8827);
and U9444 (N_9444,N_7546,N_7568);
or U9445 (N_9445,N_8218,N_7683);
and U9446 (N_9446,N_8429,N_8904);
and U9447 (N_9447,N_8178,N_8140);
nor U9448 (N_9448,N_7516,N_8779);
or U9449 (N_9449,N_7994,N_8059);
nand U9450 (N_9450,N_8954,N_8665);
and U9451 (N_9451,N_8709,N_7824);
xnor U9452 (N_9452,N_7851,N_8834);
xor U9453 (N_9453,N_8175,N_7614);
and U9454 (N_9454,N_7513,N_7846);
nor U9455 (N_9455,N_8448,N_8966);
or U9456 (N_9456,N_7756,N_7548);
nor U9457 (N_9457,N_8559,N_7689);
or U9458 (N_9458,N_8848,N_8339);
nor U9459 (N_9459,N_8340,N_8672);
nand U9460 (N_9460,N_8116,N_7527);
nor U9461 (N_9461,N_8537,N_8220);
nor U9462 (N_9462,N_8541,N_8256);
nor U9463 (N_9463,N_7895,N_8362);
and U9464 (N_9464,N_8558,N_8825);
or U9465 (N_9465,N_8344,N_7734);
and U9466 (N_9466,N_8317,N_8763);
xnor U9467 (N_9467,N_8661,N_7849);
or U9468 (N_9468,N_7710,N_8329);
nor U9469 (N_9469,N_8906,N_8430);
xnor U9470 (N_9470,N_7929,N_8435);
xnor U9471 (N_9471,N_7757,N_8533);
nor U9472 (N_9472,N_8701,N_8181);
nand U9473 (N_9473,N_8986,N_8165);
and U9474 (N_9474,N_8586,N_7509);
nor U9475 (N_9475,N_7647,N_8957);
nor U9476 (N_9476,N_8933,N_7966);
nand U9477 (N_9477,N_8194,N_8307);
nor U9478 (N_9478,N_8761,N_8342);
nor U9479 (N_9479,N_8939,N_8293);
nand U9480 (N_9480,N_7789,N_8928);
nor U9481 (N_9481,N_8882,N_8143);
xor U9482 (N_9482,N_8697,N_8147);
or U9483 (N_9483,N_8397,N_7578);
and U9484 (N_9484,N_8577,N_7965);
or U9485 (N_9485,N_8258,N_8915);
nor U9486 (N_9486,N_8710,N_8368);
nor U9487 (N_9487,N_8810,N_7842);
nand U9488 (N_9488,N_7561,N_8543);
nand U9489 (N_9489,N_7639,N_8700);
nand U9490 (N_9490,N_8360,N_8899);
nor U9491 (N_9491,N_8618,N_8918);
nor U9492 (N_9492,N_7704,N_8438);
nor U9493 (N_9493,N_8027,N_8759);
nand U9494 (N_9494,N_8347,N_7984);
and U9495 (N_9495,N_8524,N_8460);
nand U9496 (N_9496,N_8061,N_7515);
xor U9497 (N_9497,N_8262,N_8833);
nor U9498 (N_9498,N_8498,N_8492);
nor U9499 (N_9499,N_8203,N_8266);
nand U9500 (N_9500,N_7714,N_7991);
xor U9501 (N_9501,N_8718,N_8210);
nor U9502 (N_9502,N_8613,N_8567);
xor U9503 (N_9503,N_7881,N_8777);
or U9504 (N_9504,N_7713,N_8589);
and U9505 (N_9505,N_7523,N_8632);
nor U9506 (N_9506,N_7844,N_8503);
and U9507 (N_9507,N_7678,N_8052);
xor U9508 (N_9508,N_7956,N_8045);
nor U9509 (N_9509,N_8926,N_8996);
nand U9510 (N_9510,N_8280,N_8793);
nor U9511 (N_9511,N_8468,N_8426);
or U9512 (N_9512,N_8431,N_8689);
nand U9513 (N_9513,N_7967,N_8421);
nor U9514 (N_9514,N_8142,N_8110);
nor U9515 (N_9515,N_8221,N_7843);
xor U9516 (N_9516,N_7976,N_8515);
xor U9517 (N_9517,N_8630,N_8326);
and U9518 (N_9518,N_8544,N_7618);
nand U9519 (N_9519,N_8356,N_8859);
nand U9520 (N_9520,N_7913,N_7528);
nand U9521 (N_9521,N_7787,N_8626);
nand U9522 (N_9522,N_8653,N_8485);
nand U9523 (N_9523,N_8606,N_8738);
nand U9524 (N_9524,N_8031,N_8238);
nor U9525 (N_9525,N_8648,N_8295);
nand U9526 (N_9526,N_8642,N_7977);
nor U9527 (N_9527,N_8739,N_8953);
and U9528 (N_9528,N_7752,N_8727);
nand U9529 (N_9529,N_7943,N_8546);
and U9530 (N_9530,N_8261,N_7779);
nor U9531 (N_9531,N_8857,N_8783);
xor U9532 (N_9532,N_7669,N_7664);
nand U9533 (N_9533,N_8058,N_8852);
nand U9534 (N_9534,N_8135,N_8297);
nor U9535 (N_9535,N_8891,N_8775);
nand U9536 (N_9536,N_8241,N_8475);
nand U9537 (N_9537,N_8835,N_8466);
nand U9538 (N_9538,N_8412,N_8714);
nor U9539 (N_9539,N_7544,N_8801);
xnor U9540 (N_9540,N_8927,N_8687);
xor U9541 (N_9541,N_8286,N_7652);
nor U9542 (N_9542,N_8974,N_7680);
nand U9543 (N_9543,N_8652,N_8043);
or U9544 (N_9544,N_7744,N_8323);
xnor U9545 (N_9545,N_8310,N_7671);
xnor U9546 (N_9546,N_8715,N_8958);
xor U9547 (N_9547,N_8382,N_7871);
or U9548 (N_9548,N_8464,N_7791);
and U9549 (N_9549,N_8821,N_7802);
and U9550 (N_9550,N_8413,N_8271);
xor U9551 (N_9551,N_8536,N_8816);
nand U9552 (N_9552,N_8624,N_8235);
or U9553 (N_9553,N_8598,N_8478);
nor U9554 (N_9554,N_8036,N_7605);
nand U9555 (N_9555,N_7595,N_8872);
xor U9556 (N_9556,N_8929,N_7626);
or U9557 (N_9557,N_7875,N_7555);
and U9558 (N_9558,N_7980,N_7736);
or U9559 (N_9559,N_7813,N_7955);
xor U9560 (N_9560,N_7676,N_8213);
xor U9561 (N_9561,N_8096,N_8449);
nor U9562 (N_9562,N_8892,N_8075);
xor U9563 (N_9563,N_7726,N_8231);
nand U9564 (N_9564,N_8150,N_7899);
or U9565 (N_9565,N_7665,N_8534);
xor U9566 (N_9566,N_8903,N_8288);
and U9567 (N_9567,N_8937,N_8641);
and U9568 (N_9568,N_8037,N_8998);
or U9569 (N_9569,N_8053,N_8683);
nand U9570 (N_9570,N_8895,N_7925);
nor U9571 (N_9571,N_8878,N_8248);
nand U9572 (N_9572,N_8364,N_8277);
or U9573 (N_9573,N_8765,N_8932);
and U9574 (N_9574,N_7694,N_7974);
and U9575 (N_9575,N_7648,N_8724);
nor U9576 (N_9576,N_7796,N_8099);
xor U9577 (N_9577,N_7739,N_7841);
nor U9578 (N_9578,N_7903,N_8133);
xor U9579 (N_9579,N_8967,N_7971);
nor U9580 (N_9580,N_8516,N_8572);
and U9581 (N_9581,N_8785,N_8211);
nor U9582 (N_9582,N_8722,N_8686);
xnor U9583 (N_9583,N_8817,N_7865);
or U9584 (N_9584,N_7780,N_8243);
xnor U9585 (N_9585,N_8177,N_8922);
nor U9586 (N_9586,N_7912,N_8367);
or U9587 (N_9587,N_7838,N_8303);
or U9588 (N_9588,N_8465,N_8640);
nor U9589 (N_9589,N_8494,N_8667);
xor U9590 (N_9590,N_8169,N_8680);
nor U9591 (N_9591,N_8365,N_8704);
or U9592 (N_9592,N_7784,N_8732);
nand U9593 (N_9593,N_7935,N_7659);
or U9594 (N_9594,N_8223,N_7827);
or U9595 (N_9595,N_7723,N_7532);
xnor U9596 (N_9596,N_7641,N_8207);
or U9597 (N_9597,N_8198,N_7873);
xnor U9598 (N_9598,N_8076,N_7541);
or U9599 (N_9599,N_7972,N_7776);
xnor U9600 (N_9600,N_8796,N_8456);
nor U9601 (N_9601,N_8991,N_7718);
nor U9602 (N_9602,N_8602,N_8888);
xnor U9603 (N_9603,N_8935,N_8866);
nor U9604 (N_9604,N_8836,N_8514);
or U9605 (N_9605,N_7570,N_7504);
nand U9606 (N_9606,N_8331,N_8566);
or U9607 (N_9607,N_8664,N_8688);
or U9608 (N_9608,N_8812,N_8327);
xnor U9609 (N_9609,N_8479,N_7597);
nor U9610 (N_9610,N_8623,N_8267);
or U9611 (N_9611,N_8322,N_7566);
nor U9612 (N_9612,N_8694,N_8960);
and U9613 (N_9613,N_8869,N_8189);
xnor U9614 (N_9614,N_7540,N_8762);
nand U9615 (N_9615,N_8104,N_8889);
nand U9616 (N_9616,N_8404,N_8230);
nand U9617 (N_9617,N_7562,N_7900);
and U9618 (N_9618,N_7630,N_8278);
or U9619 (N_9619,N_7884,N_8729);
or U9620 (N_9620,N_8109,N_8873);
nand U9621 (N_9621,N_7951,N_8773);
xnor U9622 (N_9622,N_8819,N_7611);
nor U9623 (N_9623,N_8784,N_8681);
nand U9624 (N_9624,N_8452,N_8247);
xor U9625 (N_9625,N_8250,N_8122);
and U9626 (N_9626,N_7882,N_8508);
or U9627 (N_9627,N_8523,N_8009);
nor U9628 (N_9628,N_7785,N_8450);
and U9629 (N_9629,N_7662,N_8731);
and U9630 (N_9630,N_8745,N_8164);
or U9631 (N_9631,N_8239,N_7876);
and U9632 (N_9632,N_7637,N_8375);
nor U9633 (N_9633,N_8016,N_8673);
or U9634 (N_9634,N_8483,N_7586);
nand U9635 (N_9635,N_8332,N_8292);
nand U9636 (N_9636,N_7709,N_8995);
nor U9637 (N_9637,N_7775,N_8952);
nor U9638 (N_9638,N_7918,N_7840);
nor U9639 (N_9639,N_7549,N_8706);
nand U9640 (N_9640,N_7993,N_8740);
or U9641 (N_9641,N_8030,N_7788);
xor U9642 (N_9642,N_8434,N_7529);
nand U9643 (N_9643,N_8386,N_8167);
and U9644 (N_9644,N_8085,N_7975);
and U9645 (N_9645,N_8407,N_8789);
nand U9646 (N_9646,N_7940,N_8357);
nor U9647 (N_9647,N_8984,N_7590);
and U9648 (N_9648,N_8874,N_8497);
nor U9649 (N_9649,N_8276,N_8764);
or U9650 (N_9650,N_8346,N_8908);
and U9651 (N_9651,N_8263,N_8946);
xnor U9652 (N_9652,N_7635,N_7658);
and U9653 (N_9653,N_8639,N_7919);
xnor U9654 (N_9654,N_8502,N_7589);
and U9655 (N_9655,N_8209,N_8373);
xor U9656 (N_9656,N_7864,N_7831);
nand U9657 (N_9657,N_7682,N_8600);
xor U9658 (N_9658,N_7701,N_8518);
or U9659 (N_9659,N_8510,N_8592);
xor U9660 (N_9660,N_8071,N_7804);
nand U9661 (N_9661,N_7811,N_8318);
xnor U9662 (N_9662,N_8628,N_8300);
nand U9663 (N_9663,N_7990,N_8734);
nand U9664 (N_9664,N_8949,N_8399);
or U9665 (N_9665,N_8564,N_8912);
nor U9666 (N_9666,N_7696,N_8233);
nand U9667 (N_9667,N_8920,N_8972);
xnor U9668 (N_9668,N_7847,N_8179);
or U9669 (N_9669,N_8249,N_7816);
and U9670 (N_9670,N_8447,N_8064);
xor U9671 (N_9671,N_8348,N_7634);
and U9672 (N_9672,N_8024,N_8393);
and U9673 (N_9673,N_8077,N_7559);
or U9674 (N_9674,N_8183,N_7917);
nor U9675 (N_9675,N_7642,N_8068);
and U9676 (N_9676,N_7567,N_8417);
nor U9677 (N_9677,N_8319,N_8453);
or U9678 (N_9678,N_8257,N_8780);
nor U9679 (N_9679,N_8341,N_7645);
nand U9680 (N_9680,N_8985,N_7883);
nand U9681 (N_9681,N_7880,N_8962);
xor U9682 (N_9682,N_7894,N_8637);
or U9683 (N_9683,N_8144,N_7854);
or U9684 (N_9684,N_7753,N_8747);
or U9685 (N_9685,N_8087,N_8934);
xnor U9686 (N_9686,N_7697,N_7616);
and U9687 (N_9687,N_7745,N_8192);
and U9688 (N_9688,N_8499,N_8352);
nand U9689 (N_9689,N_7624,N_8607);
and U9690 (N_9690,N_8130,N_7538);
xnor U9691 (N_9691,N_7953,N_8190);
and U9692 (N_9692,N_8105,N_8428);
nand U9693 (N_9693,N_8806,N_7992);
and U9694 (N_9694,N_8799,N_7800);
xnor U9695 (N_9695,N_8695,N_8108);
and U9696 (N_9696,N_7760,N_8579);
nor U9697 (N_9697,N_8229,N_7686);
or U9698 (N_9698,N_8898,N_8654);
nand U9699 (N_9699,N_7685,N_8090);
or U9700 (N_9700,N_8032,N_8022);
or U9701 (N_9701,N_7550,N_7812);
nand U9702 (N_9702,N_7850,N_7596);
nor U9703 (N_9703,N_7712,N_7922);
nand U9704 (N_9704,N_7636,N_8682);
xnor U9705 (N_9705,N_7797,N_8913);
xor U9706 (N_9706,N_8959,N_8400);
or U9707 (N_9707,N_8778,N_8120);
nor U9708 (N_9708,N_8281,N_8359);
nand U9709 (N_9709,N_8750,N_8997);
and U9710 (N_9710,N_7537,N_8582);
nor U9711 (N_9711,N_7531,N_8988);
nor U9712 (N_9712,N_8408,N_7719);
xnor U9713 (N_9713,N_7539,N_8315);
xor U9714 (N_9714,N_7612,N_7646);
nor U9715 (N_9715,N_8361,N_8128);
nand U9716 (N_9716,N_8735,N_7572);
and U9717 (N_9717,N_8354,N_8246);
nand U9718 (N_9718,N_8459,N_8980);
or U9719 (N_9719,N_7777,N_8802);
or U9720 (N_9720,N_8023,N_8482);
nor U9721 (N_9721,N_8065,N_8608);
nand U9722 (N_9722,N_7808,N_7938);
and U9723 (N_9723,N_8272,N_7705);
nor U9724 (N_9724,N_7569,N_8126);
nor U9725 (N_9725,N_7861,N_8983);
and U9726 (N_9726,N_8115,N_8861);
xnor U9727 (N_9727,N_7795,N_7681);
or U9728 (N_9728,N_7997,N_7946);
and U9729 (N_9729,N_7510,N_7557);
and U9730 (N_9730,N_8007,N_7822);
and U9731 (N_9731,N_8240,N_7825);
nor U9732 (N_9732,N_7836,N_8442);
or U9733 (N_9733,N_8964,N_7792);
and U9734 (N_9734,N_8880,N_8961);
nor U9735 (N_9735,N_8570,N_8401);
xor U9736 (N_9736,N_8054,N_8847);
xnor U9737 (N_9737,N_8154,N_8214);
and U9738 (N_9738,N_8781,N_7687);
nor U9739 (N_9739,N_8800,N_8769);
nor U9740 (N_9740,N_8693,N_8148);
and U9741 (N_9741,N_8285,N_7886);
or U9742 (N_9742,N_8171,N_8725);
xnor U9743 (N_9743,N_8313,N_7693);
nor U9744 (N_9744,N_7604,N_7932);
and U9745 (N_9745,N_7717,N_8132);
xor U9746 (N_9746,N_8770,N_7720);
xor U9747 (N_9747,N_8084,N_8004);
xor U9748 (N_9748,N_7649,N_8455);
nor U9749 (N_9749,N_8619,N_8921);
nand U9750 (N_9750,N_7837,N_8757);
and U9751 (N_9751,N_8376,N_7916);
or U9752 (N_9752,N_8074,N_8406);
nand U9753 (N_9753,N_7624,N_7772);
nand U9754 (N_9754,N_8663,N_8634);
nand U9755 (N_9755,N_7681,N_7671);
xor U9756 (N_9756,N_7761,N_8955);
nand U9757 (N_9757,N_8185,N_8724);
xor U9758 (N_9758,N_7784,N_8709);
nand U9759 (N_9759,N_7519,N_8074);
nor U9760 (N_9760,N_8113,N_7810);
nand U9761 (N_9761,N_8203,N_7682);
or U9762 (N_9762,N_8800,N_8403);
nand U9763 (N_9763,N_8550,N_8705);
xor U9764 (N_9764,N_8747,N_8478);
nand U9765 (N_9765,N_8448,N_7996);
nand U9766 (N_9766,N_8015,N_8895);
and U9767 (N_9767,N_8187,N_8909);
and U9768 (N_9768,N_8595,N_8894);
and U9769 (N_9769,N_7922,N_8930);
or U9770 (N_9770,N_8485,N_7724);
nor U9771 (N_9771,N_8012,N_8414);
nor U9772 (N_9772,N_8055,N_8289);
nor U9773 (N_9773,N_7980,N_7902);
nand U9774 (N_9774,N_7894,N_7629);
nand U9775 (N_9775,N_8872,N_8374);
and U9776 (N_9776,N_8456,N_8786);
and U9777 (N_9777,N_8910,N_8698);
nor U9778 (N_9778,N_8534,N_7891);
nor U9779 (N_9779,N_8521,N_8509);
nand U9780 (N_9780,N_8830,N_7793);
or U9781 (N_9781,N_8449,N_8131);
nor U9782 (N_9782,N_8131,N_8748);
or U9783 (N_9783,N_8850,N_8405);
nor U9784 (N_9784,N_8478,N_7926);
and U9785 (N_9785,N_8445,N_8307);
nand U9786 (N_9786,N_8569,N_8171);
or U9787 (N_9787,N_8287,N_8816);
and U9788 (N_9788,N_7850,N_8787);
and U9789 (N_9789,N_8146,N_8997);
or U9790 (N_9790,N_8591,N_8111);
xnor U9791 (N_9791,N_8333,N_7548);
and U9792 (N_9792,N_7843,N_7880);
or U9793 (N_9793,N_7725,N_7728);
xnor U9794 (N_9794,N_8341,N_8567);
nor U9795 (N_9795,N_8168,N_7787);
nor U9796 (N_9796,N_7646,N_8140);
or U9797 (N_9797,N_8444,N_8034);
and U9798 (N_9798,N_7963,N_8671);
nand U9799 (N_9799,N_7585,N_7863);
or U9800 (N_9800,N_7867,N_8801);
or U9801 (N_9801,N_8370,N_8309);
nand U9802 (N_9802,N_7892,N_8350);
or U9803 (N_9803,N_8644,N_7885);
xor U9804 (N_9804,N_7508,N_7615);
or U9805 (N_9805,N_8702,N_8619);
or U9806 (N_9806,N_7664,N_8125);
nand U9807 (N_9807,N_8775,N_8263);
and U9808 (N_9808,N_7531,N_7956);
nand U9809 (N_9809,N_7965,N_8372);
and U9810 (N_9810,N_8740,N_7576);
nand U9811 (N_9811,N_7613,N_7733);
nand U9812 (N_9812,N_7502,N_8990);
nor U9813 (N_9813,N_7598,N_8733);
nor U9814 (N_9814,N_8043,N_7560);
nand U9815 (N_9815,N_8955,N_8126);
nor U9816 (N_9816,N_8533,N_8876);
or U9817 (N_9817,N_8759,N_7957);
nand U9818 (N_9818,N_7948,N_8700);
and U9819 (N_9819,N_7710,N_7589);
and U9820 (N_9820,N_8080,N_8161);
and U9821 (N_9821,N_8398,N_7777);
nor U9822 (N_9822,N_8413,N_8715);
or U9823 (N_9823,N_7673,N_8691);
and U9824 (N_9824,N_7992,N_8079);
or U9825 (N_9825,N_8151,N_8022);
and U9826 (N_9826,N_8418,N_7544);
xnor U9827 (N_9827,N_8829,N_8225);
or U9828 (N_9828,N_7534,N_8317);
and U9829 (N_9829,N_8318,N_8776);
nand U9830 (N_9830,N_7613,N_7798);
nor U9831 (N_9831,N_8406,N_8631);
nand U9832 (N_9832,N_7566,N_8686);
and U9833 (N_9833,N_8887,N_8318);
or U9834 (N_9834,N_8893,N_7984);
or U9835 (N_9835,N_8474,N_8863);
nor U9836 (N_9836,N_8491,N_7986);
nor U9837 (N_9837,N_8576,N_8473);
nand U9838 (N_9838,N_7641,N_8141);
and U9839 (N_9839,N_8637,N_8846);
and U9840 (N_9840,N_7697,N_8066);
and U9841 (N_9841,N_8004,N_7989);
nor U9842 (N_9842,N_7841,N_8017);
and U9843 (N_9843,N_8943,N_7853);
nor U9844 (N_9844,N_8161,N_7871);
or U9845 (N_9845,N_7798,N_8781);
xor U9846 (N_9846,N_8962,N_7993);
xnor U9847 (N_9847,N_7555,N_8959);
xnor U9848 (N_9848,N_8784,N_7690);
and U9849 (N_9849,N_8069,N_8122);
xnor U9850 (N_9850,N_8544,N_7552);
nand U9851 (N_9851,N_7778,N_8925);
and U9852 (N_9852,N_8372,N_8941);
nand U9853 (N_9853,N_8751,N_8891);
xor U9854 (N_9854,N_8949,N_7692);
or U9855 (N_9855,N_8869,N_8508);
nor U9856 (N_9856,N_8942,N_7563);
or U9857 (N_9857,N_8878,N_7661);
nand U9858 (N_9858,N_7714,N_8431);
nor U9859 (N_9859,N_8055,N_8422);
nor U9860 (N_9860,N_7556,N_8153);
nand U9861 (N_9861,N_7569,N_8798);
and U9862 (N_9862,N_7660,N_8480);
nor U9863 (N_9863,N_7987,N_8357);
xor U9864 (N_9864,N_8927,N_8477);
nand U9865 (N_9865,N_8410,N_8077);
xnor U9866 (N_9866,N_8131,N_8033);
or U9867 (N_9867,N_8486,N_7728);
xor U9868 (N_9868,N_7729,N_7715);
xnor U9869 (N_9869,N_8039,N_8015);
or U9870 (N_9870,N_8889,N_7662);
or U9871 (N_9871,N_8804,N_8017);
xnor U9872 (N_9872,N_8011,N_7647);
xor U9873 (N_9873,N_7576,N_8619);
nor U9874 (N_9874,N_8223,N_8829);
nand U9875 (N_9875,N_8268,N_8733);
nand U9876 (N_9876,N_8216,N_8742);
and U9877 (N_9877,N_8070,N_8913);
nor U9878 (N_9878,N_7535,N_8269);
nand U9879 (N_9879,N_8989,N_8179);
and U9880 (N_9880,N_8139,N_7815);
and U9881 (N_9881,N_8543,N_8243);
and U9882 (N_9882,N_8565,N_7516);
nor U9883 (N_9883,N_7693,N_7630);
or U9884 (N_9884,N_8473,N_8140);
or U9885 (N_9885,N_7867,N_8845);
and U9886 (N_9886,N_8112,N_7969);
and U9887 (N_9887,N_8424,N_7810);
or U9888 (N_9888,N_8427,N_8465);
nand U9889 (N_9889,N_8269,N_8150);
nand U9890 (N_9890,N_8529,N_8318);
or U9891 (N_9891,N_8803,N_8152);
xor U9892 (N_9892,N_8247,N_7900);
nor U9893 (N_9893,N_7747,N_8498);
and U9894 (N_9894,N_7934,N_7660);
xor U9895 (N_9895,N_8583,N_8996);
xnor U9896 (N_9896,N_8815,N_7624);
xnor U9897 (N_9897,N_8886,N_8119);
and U9898 (N_9898,N_8551,N_7623);
nand U9899 (N_9899,N_8238,N_8107);
nor U9900 (N_9900,N_8882,N_7691);
or U9901 (N_9901,N_8976,N_7508);
nor U9902 (N_9902,N_8243,N_8541);
or U9903 (N_9903,N_7524,N_8804);
xnor U9904 (N_9904,N_8338,N_8981);
xor U9905 (N_9905,N_8389,N_7697);
or U9906 (N_9906,N_8408,N_8166);
nor U9907 (N_9907,N_8009,N_7512);
or U9908 (N_9908,N_7544,N_8199);
and U9909 (N_9909,N_7804,N_8854);
nand U9910 (N_9910,N_8572,N_8209);
nand U9911 (N_9911,N_8870,N_7625);
and U9912 (N_9912,N_7943,N_8107);
nor U9913 (N_9913,N_8779,N_7546);
and U9914 (N_9914,N_8116,N_8371);
nor U9915 (N_9915,N_8452,N_8832);
xor U9916 (N_9916,N_8905,N_8864);
nor U9917 (N_9917,N_8296,N_8617);
nand U9918 (N_9918,N_8700,N_8039);
or U9919 (N_9919,N_7543,N_7918);
xor U9920 (N_9920,N_8054,N_7655);
nand U9921 (N_9921,N_8667,N_7731);
or U9922 (N_9922,N_7796,N_7589);
nand U9923 (N_9923,N_8264,N_7579);
nand U9924 (N_9924,N_7639,N_8752);
nor U9925 (N_9925,N_8236,N_8389);
or U9926 (N_9926,N_8367,N_7868);
nand U9927 (N_9927,N_8358,N_8530);
nand U9928 (N_9928,N_8267,N_8105);
nor U9929 (N_9929,N_7740,N_7985);
xor U9930 (N_9930,N_8803,N_8895);
and U9931 (N_9931,N_8178,N_8686);
nand U9932 (N_9932,N_8744,N_8977);
or U9933 (N_9933,N_7825,N_8438);
or U9934 (N_9934,N_7716,N_8787);
xor U9935 (N_9935,N_8937,N_7559);
or U9936 (N_9936,N_8019,N_7768);
xnor U9937 (N_9937,N_8210,N_8380);
xnor U9938 (N_9938,N_8824,N_8277);
xor U9939 (N_9939,N_7569,N_8373);
or U9940 (N_9940,N_8366,N_7933);
xnor U9941 (N_9941,N_7858,N_8131);
xnor U9942 (N_9942,N_7569,N_8526);
nor U9943 (N_9943,N_8106,N_8204);
xor U9944 (N_9944,N_8294,N_8911);
or U9945 (N_9945,N_7625,N_8009);
or U9946 (N_9946,N_7731,N_8481);
xnor U9947 (N_9947,N_7842,N_8286);
and U9948 (N_9948,N_8952,N_8055);
nor U9949 (N_9949,N_7852,N_8919);
or U9950 (N_9950,N_8377,N_7584);
nor U9951 (N_9951,N_8893,N_8578);
nand U9952 (N_9952,N_7735,N_8447);
xnor U9953 (N_9953,N_7872,N_8156);
or U9954 (N_9954,N_8905,N_8976);
xor U9955 (N_9955,N_8926,N_8990);
nand U9956 (N_9956,N_8292,N_8804);
and U9957 (N_9957,N_7592,N_7624);
or U9958 (N_9958,N_8870,N_7873);
nor U9959 (N_9959,N_8357,N_8277);
nand U9960 (N_9960,N_7734,N_8096);
xnor U9961 (N_9961,N_7828,N_8748);
and U9962 (N_9962,N_7580,N_7718);
xnor U9963 (N_9963,N_8241,N_8098);
and U9964 (N_9964,N_8761,N_8817);
or U9965 (N_9965,N_8675,N_8636);
nand U9966 (N_9966,N_7935,N_8507);
and U9967 (N_9967,N_7534,N_8134);
or U9968 (N_9968,N_7910,N_8867);
xnor U9969 (N_9969,N_8417,N_8420);
and U9970 (N_9970,N_8889,N_8624);
and U9971 (N_9971,N_8191,N_8536);
nor U9972 (N_9972,N_8061,N_8710);
xor U9973 (N_9973,N_7954,N_8832);
and U9974 (N_9974,N_7647,N_8038);
nor U9975 (N_9975,N_8291,N_8076);
and U9976 (N_9976,N_8125,N_7676);
xor U9977 (N_9977,N_7650,N_7513);
nor U9978 (N_9978,N_7866,N_7660);
xnor U9979 (N_9979,N_8741,N_8871);
nor U9980 (N_9980,N_7614,N_8687);
nor U9981 (N_9981,N_8599,N_8932);
nand U9982 (N_9982,N_8637,N_8468);
nand U9983 (N_9983,N_8622,N_7730);
and U9984 (N_9984,N_8825,N_7803);
or U9985 (N_9985,N_8063,N_7892);
nand U9986 (N_9986,N_7964,N_7611);
xnor U9987 (N_9987,N_7889,N_8348);
and U9988 (N_9988,N_8735,N_7915);
nand U9989 (N_9989,N_8951,N_8261);
or U9990 (N_9990,N_7526,N_8675);
nor U9991 (N_9991,N_7560,N_7878);
or U9992 (N_9992,N_7728,N_8295);
nand U9993 (N_9993,N_8029,N_8068);
nand U9994 (N_9994,N_7878,N_7881);
or U9995 (N_9995,N_8475,N_8423);
or U9996 (N_9996,N_8746,N_7860);
nand U9997 (N_9997,N_8187,N_8301);
or U9998 (N_9998,N_7641,N_8025);
xnor U9999 (N_9999,N_8825,N_8412);
and U10000 (N_10000,N_8374,N_8430);
nand U10001 (N_10001,N_7982,N_7760);
or U10002 (N_10002,N_7919,N_7936);
nand U10003 (N_10003,N_8581,N_8344);
or U10004 (N_10004,N_8173,N_8077);
nand U10005 (N_10005,N_8984,N_8095);
nor U10006 (N_10006,N_7818,N_8707);
or U10007 (N_10007,N_8942,N_8085);
xnor U10008 (N_10008,N_7709,N_8155);
xnor U10009 (N_10009,N_8013,N_8629);
nor U10010 (N_10010,N_8802,N_7952);
nand U10011 (N_10011,N_8296,N_8534);
nor U10012 (N_10012,N_7879,N_8363);
or U10013 (N_10013,N_8383,N_8765);
and U10014 (N_10014,N_8182,N_8243);
xor U10015 (N_10015,N_8214,N_7722);
nor U10016 (N_10016,N_8159,N_8308);
or U10017 (N_10017,N_7753,N_7674);
nor U10018 (N_10018,N_8863,N_8897);
xnor U10019 (N_10019,N_8789,N_7977);
nor U10020 (N_10020,N_8886,N_8771);
nor U10021 (N_10021,N_8364,N_7989);
and U10022 (N_10022,N_8597,N_8097);
xnor U10023 (N_10023,N_7627,N_8412);
xor U10024 (N_10024,N_7511,N_7592);
and U10025 (N_10025,N_8812,N_8020);
or U10026 (N_10026,N_8411,N_7829);
or U10027 (N_10027,N_8211,N_8128);
xor U10028 (N_10028,N_8606,N_8035);
or U10029 (N_10029,N_7746,N_8064);
xor U10030 (N_10030,N_8338,N_8082);
xor U10031 (N_10031,N_8795,N_8490);
or U10032 (N_10032,N_7664,N_7985);
or U10033 (N_10033,N_8815,N_8821);
nand U10034 (N_10034,N_8611,N_8396);
xnor U10035 (N_10035,N_8523,N_8590);
xnor U10036 (N_10036,N_7653,N_8291);
xnor U10037 (N_10037,N_8652,N_8088);
nor U10038 (N_10038,N_8862,N_8963);
nor U10039 (N_10039,N_7595,N_7652);
and U10040 (N_10040,N_8829,N_7664);
or U10041 (N_10041,N_8580,N_7980);
and U10042 (N_10042,N_8731,N_8806);
or U10043 (N_10043,N_7512,N_8401);
or U10044 (N_10044,N_7895,N_8986);
and U10045 (N_10045,N_8200,N_8340);
nand U10046 (N_10046,N_7910,N_8472);
and U10047 (N_10047,N_8581,N_7570);
or U10048 (N_10048,N_7656,N_7564);
xnor U10049 (N_10049,N_8876,N_7698);
nand U10050 (N_10050,N_8733,N_8440);
and U10051 (N_10051,N_8638,N_8676);
nor U10052 (N_10052,N_8976,N_8865);
or U10053 (N_10053,N_8035,N_8488);
or U10054 (N_10054,N_8793,N_7608);
and U10055 (N_10055,N_7615,N_7855);
xor U10056 (N_10056,N_8133,N_7669);
and U10057 (N_10057,N_8831,N_7670);
nor U10058 (N_10058,N_8516,N_8065);
or U10059 (N_10059,N_8851,N_8481);
and U10060 (N_10060,N_7707,N_8640);
xnor U10061 (N_10061,N_8972,N_7944);
and U10062 (N_10062,N_7645,N_8505);
or U10063 (N_10063,N_7541,N_7997);
xor U10064 (N_10064,N_7904,N_7843);
xnor U10065 (N_10065,N_8014,N_7663);
nand U10066 (N_10066,N_8057,N_8970);
or U10067 (N_10067,N_8696,N_8337);
nor U10068 (N_10068,N_7939,N_8139);
nand U10069 (N_10069,N_8229,N_8128);
nor U10070 (N_10070,N_7814,N_8746);
xor U10071 (N_10071,N_7695,N_8750);
nor U10072 (N_10072,N_8960,N_8871);
xor U10073 (N_10073,N_7710,N_7667);
nor U10074 (N_10074,N_8989,N_8223);
xnor U10075 (N_10075,N_8803,N_8482);
nor U10076 (N_10076,N_8698,N_8153);
xnor U10077 (N_10077,N_8090,N_8405);
and U10078 (N_10078,N_7792,N_7917);
nand U10079 (N_10079,N_8740,N_7552);
and U10080 (N_10080,N_8343,N_8180);
nor U10081 (N_10081,N_8335,N_8305);
or U10082 (N_10082,N_8828,N_7726);
xnor U10083 (N_10083,N_7525,N_7845);
or U10084 (N_10084,N_8599,N_8344);
nand U10085 (N_10085,N_8368,N_7713);
xor U10086 (N_10086,N_7879,N_8073);
nor U10087 (N_10087,N_7630,N_8742);
nand U10088 (N_10088,N_8506,N_8418);
nor U10089 (N_10089,N_8221,N_7509);
xor U10090 (N_10090,N_7788,N_8534);
xnor U10091 (N_10091,N_8316,N_7936);
xor U10092 (N_10092,N_8410,N_8645);
nand U10093 (N_10093,N_7872,N_8573);
or U10094 (N_10094,N_7629,N_7509);
nand U10095 (N_10095,N_8522,N_8820);
nand U10096 (N_10096,N_8760,N_8485);
or U10097 (N_10097,N_8802,N_8303);
nand U10098 (N_10098,N_8972,N_8470);
nor U10099 (N_10099,N_7994,N_8185);
xor U10100 (N_10100,N_8117,N_8338);
nor U10101 (N_10101,N_7976,N_8152);
nand U10102 (N_10102,N_8915,N_7940);
nor U10103 (N_10103,N_8200,N_8705);
or U10104 (N_10104,N_7832,N_7796);
or U10105 (N_10105,N_8035,N_8927);
xor U10106 (N_10106,N_8019,N_7543);
and U10107 (N_10107,N_7580,N_8789);
nand U10108 (N_10108,N_8189,N_7643);
nand U10109 (N_10109,N_8686,N_8270);
or U10110 (N_10110,N_8292,N_8520);
nor U10111 (N_10111,N_8645,N_8605);
nor U10112 (N_10112,N_7563,N_8134);
nor U10113 (N_10113,N_8790,N_8328);
and U10114 (N_10114,N_8495,N_7729);
and U10115 (N_10115,N_8583,N_8144);
xnor U10116 (N_10116,N_7609,N_8321);
or U10117 (N_10117,N_8992,N_7926);
or U10118 (N_10118,N_8506,N_8098);
or U10119 (N_10119,N_7711,N_7509);
nand U10120 (N_10120,N_8474,N_7622);
and U10121 (N_10121,N_8964,N_8534);
xor U10122 (N_10122,N_7743,N_8805);
or U10123 (N_10123,N_8537,N_8797);
and U10124 (N_10124,N_7632,N_8702);
nor U10125 (N_10125,N_8486,N_8053);
or U10126 (N_10126,N_8040,N_7936);
or U10127 (N_10127,N_8326,N_7706);
and U10128 (N_10128,N_8605,N_8737);
nor U10129 (N_10129,N_8254,N_7665);
xnor U10130 (N_10130,N_7702,N_8517);
xor U10131 (N_10131,N_7931,N_7664);
nand U10132 (N_10132,N_7964,N_8372);
and U10133 (N_10133,N_8096,N_7562);
or U10134 (N_10134,N_8025,N_7606);
or U10135 (N_10135,N_8147,N_8058);
and U10136 (N_10136,N_7545,N_8846);
nand U10137 (N_10137,N_7598,N_8910);
nand U10138 (N_10138,N_8217,N_8107);
or U10139 (N_10139,N_7731,N_8389);
and U10140 (N_10140,N_8929,N_8675);
or U10141 (N_10141,N_8833,N_8803);
nor U10142 (N_10142,N_7929,N_8893);
nor U10143 (N_10143,N_8754,N_8404);
or U10144 (N_10144,N_8249,N_8368);
nor U10145 (N_10145,N_8992,N_8598);
and U10146 (N_10146,N_8050,N_8748);
nor U10147 (N_10147,N_8791,N_8503);
xor U10148 (N_10148,N_8223,N_8580);
xnor U10149 (N_10149,N_7722,N_7559);
xnor U10150 (N_10150,N_8065,N_8520);
xor U10151 (N_10151,N_8834,N_8978);
nand U10152 (N_10152,N_7789,N_8434);
nor U10153 (N_10153,N_7623,N_8454);
xnor U10154 (N_10154,N_7712,N_7900);
nand U10155 (N_10155,N_7528,N_7530);
nor U10156 (N_10156,N_7958,N_7777);
nor U10157 (N_10157,N_8628,N_7987);
nand U10158 (N_10158,N_8937,N_8169);
xnor U10159 (N_10159,N_8225,N_8059);
and U10160 (N_10160,N_8944,N_8108);
nor U10161 (N_10161,N_8770,N_8028);
nand U10162 (N_10162,N_8069,N_8040);
nand U10163 (N_10163,N_8139,N_8039);
or U10164 (N_10164,N_8097,N_8066);
and U10165 (N_10165,N_7523,N_7697);
nor U10166 (N_10166,N_7625,N_8937);
nand U10167 (N_10167,N_7549,N_7533);
nor U10168 (N_10168,N_8802,N_8525);
and U10169 (N_10169,N_8525,N_7776);
and U10170 (N_10170,N_7943,N_8259);
xor U10171 (N_10171,N_7786,N_8842);
and U10172 (N_10172,N_8663,N_8338);
and U10173 (N_10173,N_7918,N_8524);
or U10174 (N_10174,N_8973,N_8395);
xnor U10175 (N_10175,N_8962,N_7554);
or U10176 (N_10176,N_7978,N_8648);
xnor U10177 (N_10177,N_8551,N_8225);
nand U10178 (N_10178,N_8855,N_8606);
nand U10179 (N_10179,N_8181,N_8710);
nor U10180 (N_10180,N_8469,N_7902);
or U10181 (N_10181,N_8539,N_8049);
xor U10182 (N_10182,N_7882,N_7781);
or U10183 (N_10183,N_7618,N_7761);
or U10184 (N_10184,N_8471,N_8152);
or U10185 (N_10185,N_8916,N_8296);
xnor U10186 (N_10186,N_7548,N_8477);
or U10187 (N_10187,N_8396,N_8599);
nor U10188 (N_10188,N_8268,N_8361);
or U10189 (N_10189,N_8117,N_7567);
and U10190 (N_10190,N_8576,N_7634);
or U10191 (N_10191,N_8380,N_8575);
nand U10192 (N_10192,N_8373,N_8867);
nand U10193 (N_10193,N_7803,N_7936);
or U10194 (N_10194,N_8967,N_8757);
xnor U10195 (N_10195,N_8662,N_8679);
nor U10196 (N_10196,N_7512,N_8762);
nand U10197 (N_10197,N_8483,N_7679);
nor U10198 (N_10198,N_8416,N_7985);
nor U10199 (N_10199,N_8095,N_7744);
nor U10200 (N_10200,N_8234,N_7958);
xnor U10201 (N_10201,N_8419,N_7819);
or U10202 (N_10202,N_7866,N_8983);
nand U10203 (N_10203,N_8099,N_8575);
nor U10204 (N_10204,N_7949,N_8161);
xnor U10205 (N_10205,N_8610,N_7686);
or U10206 (N_10206,N_8247,N_7691);
nand U10207 (N_10207,N_8892,N_8845);
nand U10208 (N_10208,N_8475,N_8519);
or U10209 (N_10209,N_8888,N_8126);
xnor U10210 (N_10210,N_8369,N_8998);
or U10211 (N_10211,N_8675,N_8800);
nor U10212 (N_10212,N_7885,N_8053);
or U10213 (N_10213,N_8584,N_8449);
and U10214 (N_10214,N_8886,N_8211);
nand U10215 (N_10215,N_8211,N_8038);
nor U10216 (N_10216,N_8364,N_8960);
xnor U10217 (N_10217,N_8710,N_8337);
and U10218 (N_10218,N_8211,N_8745);
or U10219 (N_10219,N_7855,N_8224);
or U10220 (N_10220,N_8755,N_8435);
nand U10221 (N_10221,N_7893,N_7800);
and U10222 (N_10222,N_8118,N_8573);
and U10223 (N_10223,N_8137,N_8030);
nand U10224 (N_10224,N_8278,N_7971);
nor U10225 (N_10225,N_8045,N_8689);
and U10226 (N_10226,N_8624,N_8043);
xor U10227 (N_10227,N_8057,N_8849);
or U10228 (N_10228,N_7724,N_8406);
nand U10229 (N_10229,N_8913,N_8791);
nand U10230 (N_10230,N_8745,N_8560);
or U10231 (N_10231,N_8717,N_8869);
nand U10232 (N_10232,N_8955,N_8624);
or U10233 (N_10233,N_7703,N_8543);
or U10234 (N_10234,N_8373,N_8735);
xnor U10235 (N_10235,N_7631,N_8157);
nand U10236 (N_10236,N_7994,N_8634);
xnor U10237 (N_10237,N_7966,N_8952);
xor U10238 (N_10238,N_8008,N_8681);
xnor U10239 (N_10239,N_7525,N_7515);
or U10240 (N_10240,N_7504,N_8916);
or U10241 (N_10241,N_8345,N_8958);
nand U10242 (N_10242,N_8935,N_8904);
xnor U10243 (N_10243,N_7923,N_7903);
nand U10244 (N_10244,N_8435,N_8154);
or U10245 (N_10245,N_7634,N_8487);
xor U10246 (N_10246,N_8477,N_8280);
or U10247 (N_10247,N_8816,N_7606);
and U10248 (N_10248,N_7853,N_8308);
xor U10249 (N_10249,N_7671,N_8486);
and U10250 (N_10250,N_7701,N_8156);
and U10251 (N_10251,N_8039,N_8370);
nand U10252 (N_10252,N_8131,N_8820);
and U10253 (N_10253,N_8902,N_8440);
or U10254 (N_10254,N_8461,N_8378);
nor U10255 (N_10255,N_8625,N_8678);
or U10256 (N_10256,N_7635,N_8411);
or U10257 (N_10257,N_8891,N_8345);
nand U10258 (N_10258,N_8143,N_8467);
xor U10259 (N_10259,N_7571,N_8063);
nor U10260 (N_10260,N_7547,N_8809);
and U10261 (N_10261,N_7856,N_8114);
nor U10262 (N_10262,N_7652,N_7576);
and U10263 (N_10263,N_7600,N_8653);
nor U10264 (N_10264,N_7956,N_8937);
or U10265 (N_10265,N_8058,N_8025);
or U10266 (N_10266,N_7660,N_8820);
or U10267 (N_10267,N_8682,N_8242);
or U10268 (N_10268,N_8789,N_8177);
and U10269 (N_10269,N_7544,N_7597);
or U10270 (N_10270,N_8565,N_8843);
nand U10271 (N_10271,N_8918,N_8649);
and U10272 (N_10272,N_8439,N_8239);
xnor U10273 (N_10273,N_8446,N_8494);
nor U10274 (N_10274,N_8662,N_8828);
or U10275 (N_10275,N_8311,N_7603);
nand U10276 (N_10276,N_7980,N_7920);
or U10277 (N_10277,N_7517,N_7938);
nor U10278 (N_10278,N_8741,N_7831);
and U10279 (N_10279,N_8525,N_8929);
or U10280 (N_10280,N_8645,N_7643);
xor U10281 (N_10281,N_8106,N_8327);
nor U10282 (N_10282,N_8132,N_8624);
xor U10283 (N_10283,N_8128,N_8796);
nor U10284 (N_10284,N_8267,N_8566);
and U10285 (N_10285,N_8909,N_8867);
nand U10286 (N_10286,N_8031,N_8329);
nand U10287 (N_10287,N_8590,N_8176);
or U10288 (N_10288,N_7873,N_8114);
nand U10289 (N_10289,N_8344,N_7597);
or U10290 (N_10290,N_8631,N_8069);
nor U10291 (N_10291,N_8870,N_8120);
nor U10292 (N_10292,N_8632,N_8177);
xor U10293 (N_10293,N_8543,N_8477);
and U10294 (N_10294,N_8255,N_7696);
nor U10295 (N_10295,N_7701,N_8439);
nand U10296 (N_10296,N_7913,N_8056);
and U10297 (N_10297,N_8537,N_7510);
nor U10298 (N_10298,N_8733,N_7930);
or U10299 (N_10299,N_7617,N_8023);
or U10300 (N_10300,N_7617,N_7533);
xor U10301 (N_10301,N_7959,N_8365);
or U10302 (N_10302,N_7901,N_8864);
or U10303 (N_10303,N_8019,N_8173);
and U10304 (N_10304,N_8318,N_7917);
or U10305 (N_10305,N_7747,N_8463);
nor U10306 (N_10306,N_7764,N_7925);
xor U10307 (N_10307,N_7783,N_8984);
or U10308 (N_10308,N_7718,N_8014);
nand U10309 (N_10309,N_8294,N_8336);
or U10310 (N_10310,N_7797,N_7706);
xor U10311 (N_10311,N_8100,N_8742);
nand U10312 (N_10312,N_7682,N_7910);
xor U10313 (N_10313,N_8703,N_7747);
and U10314 (N_10314,N_8963,N_8324);
nor U10315 (N_10315,N_8868,N_7852);
nor U10316 (N_10316,N_8821,N_8707);
and U10317 (N_10317,N_8648,N_7841);
or U10318 (N_10318,N_8740,N_8830);
nor U10319 (N_10319,N_8628,N_7838);
nor U10320 (N_10320,N_7504,N_8591);
nand U10321 (N_10321,N_8760,N_8351);
nor U10322 (N_10322,N_8998,N_7658);
nor U10323 (N_10323,N_8767,N_8174);
and U10324 (N_10324,N_8419,N_7873);
nand U10325 (N_10325,N_7843,N_8163);
xnor U10326 (N_10326,N_8989,N_7979);
or U10327 (N_10327,N_8558,N_8570);
xor U10328 (N_10328,N_7552,N_8304);
xor U10329 (N_10329,N_7634,N_8126);
nor U10330 (N_10330,N_8774,N_7670);
nor U10331 (N_10331,N_8624,N_8159);
nand U10332 (N_10332,N_7745,N_8695);
or U10333 (N_10333,N_8201,N_8413);
or U10334 (N_10334,N_8274,N_8385);
xnor U10335 (N_10335,N_8698,N_8879);
nand U10336 (N_10336,N_7850,N_8728);
or U10337 (N_10337,N_7867,N_8710);
xnor U10338 (N_10338,N_8719,N_7895);
and U10339 (N_10339,N_8149,N_8857);
and U10340 (N_10340,N_8215,N_8979);
nor U10341 (N_10341,N_7529,N_7827);
nand U10342 (N_10342,N_8429,N_8466);
xor U10343 (N_10343,N_7659,N_8098);
nor U10344 (N_10344,N_8036,N_8956);
nor U10345 (N_10345,N_8176,N_7664);
nor U10346 (N_10346,N_7604,N_8874);
xnor U10347 (N_10347,N_7657,N_8927);
nor U10348 (N_10348,N_7808,N_8971);
nand U10349 (N_10349,N_8628,N_8830);
and U10350 (N_10350,N_8667,N_8893);
or U10351 (N_10351,N_8061,N_8327);
or U10352 (N_10352,N_8825,N_8880);
nand U10353 (N_10353,N_7699,N_7865);
nor U10354 (N_10354,N_8832,N_8570);
and U10355 (N_10355,N_8110,N_8467);
xor U10356 (N_10356,N_7641,N_8063);
or U10357 (N_10357,N_7959,N_8681);
nand U10358 (N_10358,N_8591,N_8856);
nand U10359 (N_10359,N_8751,N_7688);
nor U10360 (N_10360,N_8247,N_8655);
nand U10361 (N_10361,N_8768,N_8353);
or U10362 (N_10362,N_7815,N_8459);
nor U10363 (N_10363,N_7614,N_7949);
and U10364 (N_10364,N_7778,N_8640);
nand U10365 (N_10365,N_7738,N_8757);
nor U10366 (N_10366,N_7576,N_7765);
nor U10367 (N_10367,N_8693,N_8452);
nor U10368 (N_10368,N_8636,N_7611);
xnor U10369 (N_10369,N_7754,N_8222);
nor U10370 (N_10370,N_8677,N_7792);
nor U10371 (N_10371,N_7938,N_7803);
and U10372 (N_10372,N_8227,N_8900);
xor U10373 (N_10373,N_8749,N_8209);
or U10374 (N_10374,N_8748,N_7760);
nor U10375 (N_10375,N_7598,N_8978);
or U10376 (N_10376,N_7982,N_8667);
and U10377 (N_10377,N_8888,N_8577);
nor U10378 (N_10378,N_8521,N_7647);
xor U10379 (N_10379,N_7703,N_7717);
and U10380 (N_10380,N_8485,N_8098);
xor U10381 (N_10381,N_8474,N_7553);
nor U10382 (N_10382,N_8520,N_7910);
and U10383 (N_10383,N_7990,N_7978);
and U10384 (N_10384,N_8769,N_8676);
or U10385 (N_10385,N_8183,N_8131);
or U10386 (N_10386,N_8989,N_8649);
and U10387 (N_10387,N_7981,N_7608);
xor U10388 (N_10388,N_8685,N_8503);
nor U10389 (N_10389,N_8788,N_8036);
nor U10390 (N_10390,N_8697,N_8641);
nand U10391 (N_10391,N_8667,N_7540);
nand U10392 (N_10392,N_7699,N_8994);
nor U10393 (N_10393,N_8054,N_8383);
xnor U10394 (N_10394,N_7587,N_7610);
xor U10395 (N_10395,N_8001,N_8354);
xnor U10396 (N_10396,N_8696,N_7705);
nand U10397 (N_10397,N_7774,N_8196);
nor U10398 (N_10398,N_8898,N_7742);
nor U10399 (N_10399,N_7575,N_8218);
and U10400 (N_10400,N_7664,N_7845);
or U10401 (N_10401,N_7911,N_7765);
or U10402 (N_10402,N_7995,N_8788);
xor U10403 (N_10403,N_8215,N_7718);
xor U10404 (N_10404,N_8787,N_7973);
or U10405 (N_10405,N_8191,N_8154);
xnor U10406 (N_10406,N_8382,N_8978);
nor U10407 (N_10407,N_8645,N_7812);
xnor U10408 (N_10408,N_7588,N_8363);
xnor U10409 (N_10409,N_8062,N_8570);
xor U10410 (N_10410,N_7524,N_7784);
and U10411 (N_10411,N_7666,N_8986);
and U10412 (N_10412,N_8570,N_8629);
nand U10413 (N_10413,N_8237,N_8623);
nor U10414 (N_10414,N_8763,N_8930);
nor U10415 (N_10415,N_8770,N_7985);
nand U10416 (N_10416,N_8289,N_8942);
xnor U10417 (N_10417,N_7798,N_8553);
and U10418 (N_10418,N_8643,N_8687);
and U10419 (N_10419,N_8181,N_8029);
or U10420 (N_10420,N_8905,N_8559);
nor U10421 (N_10421,N_7513,N_7802);
xor U10422 (N_10422,N_8555,N_7604);
nor U10423 (N_10423,N_8027,N_8662);
or U10424 (N_10424,N_7615,N_8866);
xnor U10425 (N_10425,N_7606,N_8108);
xnor U10426 (N_10426,N_8400,N_7856);
or U10427 (N_10427,N_8303,N_8809);
nor U10428 (N_10428,N_8777,N_8697);
xor U10429 (N_10429,N_8306,N_8676);
or U10430 (N_10430,N_7846,N_8674);
xor U10431 (N_10431,N_8021,N_8562);
xnor U10432 (N_10432,N_8103,N_8215);
nand U10433 (N_10433,N_8130,N_8841);
or U10434 (N_10434,N_7632,N_8595);
or U10435 (N_10435,N_8650,N_8780);
xnor U10436 (N_10436,N_8041,N_7892);
or U10437 (N_10437,N_8324,N_8689);
and U10438 (N_10438,N_7858,N_8832);
xnor U10439 (N_10439,N_8618,N_8808);
xnor U10440 (N_10440,N_7938,N_7518);
or U10441 (N_10441,N_8680,N_8576);
nor U10442 (N_10442,N_7732,N_8829);
xnor U10443 (N_10443,N_8818,N_7979);
xnor U10444 (N_10444,N_8751,N_8735);
xnor U10445 (N_10445,N_8518,N_8929);
or U10446 (N_10446,N_8057,N_7738);
nand U10447 (N_10447,N_8110,N_7904);
nor U10448 (N_10448,N_8937,N_8754);
or U10449 (N_10449,N_8163,N_8431);
nor U10450 (N_10450,N_8358,N_8058);
nor U10451 (N_10451,N_7743,N_8432);
and U10452 (N_10452,N_8118,N_8246);
or U10453 (N_10453,N_8687,N_7505);
or U10454 (N_10454,N_8051,N_7867);
or U10455 (N_10455,N_8053,N_7553);
xor U10456 (N_10456,N_8548,N_8827);
or U10457 (N_10457,N_8348,N_8063);
and U10458 (N_10458,N_8100,N_7610);
and U10459 (N_10459,N_8258,N_7829);
xnor U10460 (N_10460,N_7614,N_8985);
xnor U10461 (N_10461,N_7868,N_8117);
nor U10462 (N_10462,N_7803,N_7808);
and U10463 (N_10463,N_8745,N_8302);
nand U10464 (N_10464,N_8553,N_8083);
and U10465 (N_10465,N_7577,N_8209);
or U10466 (N_10466,N_8741,N_7590);
and U10467 (N_10467,N_8899,N_7948);
nand U10468 (N_10468,N_8162,N_8336);
nor U10469 (N_10469,N_8005,N_8861);
xnor U10470 (N_10470,N_7908,N_7721);
xor U10471 (N_10471,N_8839,N_8859);
and U10472 (N_10472,N_8495,N_8100);
nor U10473 (N_10473,N_8669,N_7560);
nand U10474 (N_10474,N_8714,N_8038);
nand U10475 (N_10475,N_8351,N_8673);
or U10476 (N_10476,N_7764,N_8707);
xnor U10477 (N_10477,N_8138,N_7515);
and U10478 (N_10478,N_7906,N_7578);
nor U10479 (N_10479,N_7562,N_7800);
xnor U10480 (N_10480,N_7975,N_8264);
or U10481 (N_10481,N_7567,N_8833);
xnor U10482 (N_10482,N_8350,N_8599);
nor U10483 (N_10483,N_8664,N_8152);
and U10484 (N_10484,N_8511,N_7692);
nand U10485 (N_10485,N_8429,N_8911);
or U10486 (N_10486,N_8540,N_8899);
or U10487 (N_10487,N_8844,N_7661);
and U10488 (N_10488,N_8387,N_7911);
and U10489 (N_10489,N_8864,N_8950);
and U10490 (N_10490,N_8435,N_8560);
or U10491 (N_10491,N_8186,N_8593);
and U10492 (N_10492,N_7575,N_8460);
nand U10493 (N_10493,N_7870,N_8162);
nor U10494 (N_10494,N_7726,N_8961);
and U10495 (N_10495,N_8080,N_7977);
nor U10496 (N_10496,N_8252,N_8873);
xnor U10497 (N_10497,N_8040,N_7851);
and U10498 (N_10498,N_8220,N_8458);
and U10499 (N_10499,N_8575,N_7702);
or U10500 (N_10500,N_10178,N_9136);
xnor U10501 (N_10501,N_9936,N_9831);
xnor U10502 (N_10502,N_9685,N_10054);
xor U10503 (N_10503,N_10356,N_10166);
nor U10504 (N_10504,N_9354,N_9609);
xnor U10505 (N_10505,N_10499,N_10319);
nand U10506 (N_10506,N_10049,N_9603);
nand U10507 (N_10507,N_9122,N_9601);
or U10508 (N_10508,N_9907,N_9184);
xnor U10509 (N_10509,N_9116,N_10142);
or U10510 (N_10510,N_10068,N_9864);
nor U10511 (N_10511,N_10280,N_10351);
nor U10512 (N_10512,N_9489,N_9349);
and U10513 (N_10513,N_10424,N_10087);
or U10514 (N_10514,N_10435,N_9911);
nor U10515 (N_10515,N_10271,N_9219);
xor U10516 (N_10516,N_10228,N_10485);
or U10517 (N_10517,N_10400,N_9398);
or U10518 (N_10518,N_9072,N_9187);
nand U10519 (N_10519,N_9730,N_9148);
nor U10520 (N_10520,N_9445,N_9215);
nand U10521 (N_10521,N_10312,N_9559);
nor U10522 (N_10522,N_10127,N_9826);
nand U10523 (N_10523,N_9278,N_9202);
or U10524 (N_10524,N_10223,N_9425);
nand U10525 (N_10525,N_9413,N_9423);
nor U10526 (N_10526,N_10182,N_9650);
xnor U10527 (N_10527,N_9690,N_10406);
nand U10528 (N_10528,N_9721,N_10484);
nand U10529 (N_10529,N_9162,N_9263);
nor U10530 (N_10530,N_9056,N_10396);
and U10531 (N_10531,N_9078,N_9541);
xor U10532 (N_10532,N_10222,N_9086);
nor U10533 (N_10533,N_9450,N_9150);
or U10534 (N_10534,N_9369,N_9688);
or U10535 (N_10535,N_10468,N_9572);
nand U10536 (N_10536,N_10027,N_9241);
or U10537 (N_10537,N_9870,N_9446);
or U10538 (N_10538,N_9871,N_10200);
nand U10539 (N_10539,N_9363,N_9507);
or U10540 (N_10540,N_9329,N_10327);
nand U10541 (N_10541,N_10452,N_9291);
nand U10542 (N_10542,N_9647,N_9678);
xor U10543 (N_10543,N_10118,N_9383);
nor U10544 (N_10544,N_10414,N_9320);
or U10545 (N_10545,N_9523,N_9075);
and U10546 (N_10546,N_10162,N_9807);
nor U10547 (N_10547,N_9391,N_9280);
nor U10548 (N_10548,N_9612,N_9798);
or U10549 (N_10549,N_9128,N_9805);
or U10550 (N_10550,N_10195,N_9697);
and U10551 (N_10551,N_9502,N_9331);
xor U10552 (N_10552,N_9927,N_9324);
or U10553 (N_10553,N_9550,N_9754);
or U10554 (N_10554,N_10139,N_10364);
nand U10555 (N_10555,N_10269,N_9412);
xor U10556 (N_10556,N_10264,N_10196);
nor U10557 (N_10557,N_10279,N_9856);
xor U10558 (N_10558,N_10447,N_9036);
and U10559 (N_10559,N_9583,N_9475);
nand U10560 (N_10560,N_9582,N_9282);
xnor U10561 (N_10561,N_9220,N_10020);
or U10562 (N_10562,N_9943,N_10132);
nor U10563 (N_10563,N_9654,N_10354);
or U10564 (N_10564,N_9537,N_10079);
and U10565 (N_10565,N_9766,N_9186);
and U10566 (N_10566,N_9135,N_9313);
xor U10567 (N_10567,N_9683,N_9246);
nand U10568 (N_10568,N_10011,N_10183);
or U10569 (N_10569,N_10022,N_9935);
nand U10570 (N_10570,N_10475,N_10425);
or U10571 (N_10571,N_9906,N_9046);
nor U10572 (N_10572,N_10140,N_10403);
or U10573 (N_10573,N_10117,N_9535);
or U10574 (N_10574,N_10301,N_9012);
xnor U10575 (N_10575,N_9640,N_9053);
and U10576 (N_10576,N_9659,N_9615);
nand U10577 (N_10577,N_9231,N_9065);
nor U10578 (N_10578,N_10263,N_10032);
nor U10579 (N_10579,N_9720,N_9226);
or U10580 (N_10580,N_10275,N_9813);
and U10581 (N_10581,N_9029,N_10202);
nand U10582 (N_10582,N_9620,N_10066);
or U10583 (N_10583,N_9516,N_10433);
nor U10584 (N_10584,N_10226,N_9458);
and U10585 (N_10585,N_9768,N_10455);
nor U10586 (N_10586,N_9443,N_9913);
nor U10587 (N_10587,N_9140,N_9747);
nor U10588 (N_10588,N_9984,N_9777);
nor U10589 (N_10589,N_9314,N_9157);
or U10590 (N_10590,N_9763,N_9748);
nand U10591 (N_10591,N_9515,N_9019);
and U10592 (N_10592,N_9343,N_10276);
nand U10593 (N_10593,N_9170,N_9481);
nor U10594 (N_10594,N_9463,N_10394);
nor U10595 (N_10595,N_10262,N_9933);
nand U10596 (N_10596,N_9464,N_9909);
and U10597 (N_10597,N_10229,N_10482);
nand U10598 (N_10598,N_9045,N_9209);
and U10599 (N_10599,N_9492,N_9899);
nand U10600 (N_10600,N_9477,N_10445);
nor U10601 (N_10601,N_9451,N_9179);
or U10602 (N_10602,N_9607,N_10401);
nor U10603 (N_10603,N_9994,N_9691);
and U10604 (N_10604,N_9119,N_9670);
and U10605 (N_10605,N_9321,N_9457);
nor U10606 (N_10606,N_9123,N_9786);
nor U10607 (N_10607,N_9661,N_9904);
nor U10608 (N_10608,N_10465,N_9410);
nand U10609 (N_10609,N_10036,N_10135);
nand U10610 (N_10610,N_10207,N_9945);
nor U10611 (N_10611,N_9762,N_10480);
and U10612 (N_10612,N_9037,N_10421);
nor U10613 (N_10613,N_10398,N_10431);
xnor U10614 (N_10614,N_10357,N_10080);
and U10615 (N_10615,N_9663,N_10487);
or U10616 (N_10616,N_9438,N_10383);
and U10617 (N_10617,N_10008,N_10405);
and U10618 (N_10618,N_9804,N_10417);
nand U10619 (N_10619,N_10215,N_9573);
nand U10620 (N_10620,N_9919,N_10044);
and U10621 (N_10621,N_9701,N_9962);
and U10622 (N_10622,N_10091,N_9323);
and U10623 (N_10623,N_10246,N_9111);
and U10624 (N_10624,N_9695,N_9352);
nand U10625 (N_10625,N_9333,N_9792);
xor U10626 (N_10626,N_9047,N_10442);
or U10627 (N_10627,N_10368,N_10112);
and U10628 (N_10628,N_9420,N_9724);
nand U10629 (N_10629,N_9161,N_10429);
nand U10630 (N_10630,N_9195,N_9755);
or U10631 (N_10631,N_9881,N_9093);
or U10632 (N_10632,N_9501,N_10441);
nand U10633 (N_10633,N_9461,N_10411);
and U10634 (N_10634,N_10393,N_10052);
nor U10635 (N_10635,N_9561,N_10165);
or U10636 (N_10636,N_9764,N_9783);
or U10637 (N_10637,N_9505,N_10326);
nand U10638 (N_10638,N_9417,N_10169);
or U10639 (N_10639,N_9375,N_9370);
nand U10640 (N_10640,N_9656,N_9338);
or U10641 (N_10641,N_9570,N_10230);
xor U10642 (N_10642,N_9480,N_9668);
or U10643 (N_10643,N_9266,N_9828);
and U10644 (N_10644,N_10185,N_10151);
and U10645 (N_10645,N_10110,N_9429);
xor U10646 (N_10646,N_9660,N_10496);
or U10647 (N_10647,N_9509,N_9932);
nand U10648 (N_10648,N_9360,N_9041);
nor U10649 (N_10649,N_9127,N_9000);
xnor U10650 (N_10650,N_10095,N_9013);
nand U10651 (N_10651,N_9348,N_9776);
or U10652 (N_10652,N_9073,N_9026);
and U10653 (N_10653,N_10476,N_9257);
xnor U10654 (N_10654,N_9512,N_10259);
nor U10655 (N_10655,N_9990,N_10416);
nand U10656 (N_10656,N_9518,N_10121);
nand U10657 (N_10657,N_10258,N_9532);
and U10658 (N_10658,N_9880,N_9811);
and U10659 (N_10659,N_9163,N_9846);
xnor U10660 (N_10660,N_9181,N_9414);
nor U10661 (N_10661,N_10244,N_9062);
and U10662 (N_10662,N_9283,N_9729);
xor U10663 (N_10663,N_10302,N_9571);
nor U10664 (N_10664,N_10371,N_10028);
nor U10665 (N_10665,N_9569,N_9589);
xnor U10666 (N_10666,N_9767,N_10076);
or U10667 (N_10667,N_9844,N_10104);
nand U10668 (N_10668,N_10314,N_9963);
xnor U10669 (N_10669,N_10218,N_10133);
nand U10670 (N_10670,N_10489,N_9672);
xor U10671 (N_10671,N_9273,N_10242);
and U10672 (N_10672,N_10106,N_9960);
and U10673 (N_10673,N_10131,N_9334);
and U10674 (N_10674,N_9210,N_10192);
nand U10675 (N_10675,N_9397,N_9519);
nand U10676 (N_10676,N_9938,N_9097);
and U10677 (N_10677,N_10333,N_10399);
nand U10678 (N_10678,N_9230,N_10119);
or U10679 (N_10679,N_10346,N_10341);
or U10680 (N_10680,N_10248,N_9934);
nor U10681 (N_10681,N_10213,N_10078);
or U10682 (N_10682,N_9415,N_9905);
or U10683 (N_10683,N_10220,N_10331);
nand U10684 (N_10684,N_10187,N_10126);
nor U10685 (N_10685,N_9598,N_9973);
or U10686 (N_10686,N_10464,N_9091);
nand U10687 (N_10687,N_9981,N_10330);
or U10688 (N_10688,N_10461,N_10491);
xor U10689 (N_10689,N_9568,N_9703);
nand U10690 (N_10690,N_10077,N_9172);
nor U10691 (N_10691,N_10313,N_10474);
nor U10692 (N_10692,N_10245,N_9218);
nor U10693 (N_10693,N_9787,N_9453);
xnor U10694 (N_10694,N_9867,N_9432);
or U10695 (N_10695,N_9590,N_9107);
nor U10696 (N_10696,N_9789,N_9920);
nand U10697 (N_10697,N_10157,N_9437);
and U10698 (N_10698,N_10369,N_10296);
nand U10699 (N_10699,N_10039,N_10316);
xor U10700 (N_10700,N_9821,N_9782);
xnor U10701 (N_10701,N_10349,N_9449);
nor U10702 (N_10702,N_9617,N_9486);
or U10703 (N_10703,N_10025,N_10328);
and U10704 (N_10704,N_10385,N_10168);
xor U10705 (N_10705,N_9033,N_9587);
or U10706 (N_10706,N_9325,N_9109);
nor U10707 (N_10707,N_9365,N_10317);
nor U10708 (N_10708,N_9832,N_10146);
or U10709 (N_10709,N_9336,N_9521);
nor U10710 (N_10710,N_10448,N_10409);
nand U10711 (N_10711,N_9245,N_9009);
and U10712 (N_10712,N_9709,N_9513);
nor U10713 (N_10713,N_9493,N_9728);
or U10714 (N_10714,N_9866,N_9017);
nand U10715 (N_10715,N_9433,N_10209);
or U10716 (N_10716,N_9232,N_10380);
or U10717 (N_10717,N_9628,N_9547);
xnor U10718 (N_10718,N_10239,N_9542);
or U10719 (N_10719,N_9916,N_9969);
and U10720 (N_10720,N_10324,N_10029);
nand U10721 (N_10721,N_9626,N_9667);
nand U10722 (N_10722,N_10234,N_10379);
nand U10723 (N_10723,N_10407,N_9576);
nand U10724 (N_10724,N_9233,N_9490);
nor U10725 (N_10725,N_10083,N_9727);
nand U10726 (N_10726,N_9982,N_10096);
nor U10727 (N_10727,N_9169,N_9514);
nor U10728 (N_10728,N_10221,N_10120);
xnor U10729 (N_10729,N_10339,N_9436);
xnor U10730 (N_10730,N_10188,N_10268);
nor U10731 (N_10731,N_9105,N_9791);
nand U10732 (N_10732,N_9838,N_9040);
xnor U10733 (N_10733,N_10211,N_9752);
xor U10734 (N_10734,N_10412,N_9106);
xnor U10735 (N_10735,N_10235,N_10298);
and U10736 (N_10736,N_9305,N_9546);
nand U10737 (N_10737,N_9194,N_9407);
and U10738 (N_10738,N_9669,N_10426);
and U10739 (N_10739,N_9657,N_9694);
xnor U10740 (N_10740,N_9430,N_10374);
xnor U10741 (N_10741,N_9753,N_9188);
nor U10742 (N_10742,N_9971,N_9070);
nor U10743 (N_10743,N_10446,N_9539);
or U10744 (N_10744,N_9137,N_9902);
nor U10745 (N_10745,N_9424,N_9942);
or U10746 (N_10746,N_9854,N_9869);
nor U10747 (N_10747,N_9643,N_9886);
nor U10748 (N_10748,N_9228,N_9406);
xor U10749 (N_10749,N_9771,N_9998);
xnor U10750 (N_10750,N_9800,N_10019);
or U10751 (N_10751,N_9774,N_10274);
nand U10752 (N_10752,N_9303,N_10055);
xor U10753 (N_10753,N_10261,N_10031);
and U10754 (N_10754,N_9985,N_9810);
and U10755 (N_10755,N_9722,N_9680);
nor U10756 (N_10756,N_9085,N_9606);
xor U10757 (N_10757,N_9893,N_9779);
and U10758 (N_10758,N_10361,N_9892);
and U10759 (N_10759,N_9081,N_9742);
or U10760 (N_10760,N_10457,N_9819);
nor U10761 (N_10761,N_9165,N_9176);
or U10762 (N_10762,N_10343,N_9859);
xor U10763 (N_10763,N_9051,N_9098);
xnor U10764 (N_10764,N_9925,N_9421);
or U10765 (N_10765,N_10430,N_9635);
and U10766 (N_10766,N_9958,N_9847);
nor U10767 (N_10767,N_9396,N_10255);
xor U10768 (N_10768,N_10353,N_9623);
xnor U10769 (N_10769,N_9957,N_9031);
and U10770 (N_10770,N_10041,N_9297);
nor U10771 (N_10771,N_10288,N_10490);
and U10772 (N_10772,N_9473,N_9770);
nor U10773 (N_10773,N_9716,N_10267);
xnor U10774 (N_10774,N_10320,N_9714);
xnor U10775 (N_10775,N_9835,N_10241);
nand U10776 (N_10776,N_9740,N_10065);
and U10777 (N_10777,N_10062,N_9482);
nand U10778 (N_10778,N_9564,N_9624);
nand U10779 (N_10779,N_10309,N_9316);
nor U10780 (N_10780,N_9600,N_9256);
nor U10781 (N_10781,N_10030,N_10105);
xnor U10782 (N_10782,N_9462,N_9860);
xnor U10783 (N_10783,N_9682,N_10086);
nand U10784 (N_10784,N_10124,N_10250);
and U10785 (N_10785,N_10170,N_10073);
and U10786 (N_10786,N_9353,N_9112);
nand U10787 (N_10787,N_10212,N_9686);
and U10788 (N_10788,N_10048,N_10365);
nand U10789 (N_10789,N_10056,N_9426);
xor U10790 (N_10790,N_9185,N_9487);
or U10791 (N_10791,N_10350,N_9164);
xnor U10792 (N_10792,N_9113,N_9853);
or U10793 (N_10793,N_9288,N_9760);
and U10794 (N_10794,N_10175,N_9021);
xor U10795 (N_10795,N_10059,N_9198);
and U10796 (N_10796,N_9393,N_9706);
or U10797 (N_10797,N_10172,N_10377);
or U10798 (N_10798,N_10224,N_10470);
and U10799 (N_10799,N_10141,N_9708);
and U10800 (N_10800,N_9063,N_9843);
or U10801 (N_10801,N_10286,N_9646);
and U10802 (N_10802,N_9260,N_9978);
xor U10803 (N_10803,N_10103,N_10006);
xnor U10804 (N_10804,N_9967,N_9567);
or U10805 (N_10805,N_9772,N_9794);
nor U10806 (N_10806,N_9824,N_10034);
nor U10807 (N_10807,N_9633,N_9553);
xnor U10808 (N_10808,N_10043,N_9315);
and U10809 (N_10809,N_10021,N_9739);
nor U10810 (N_10810,N_10089,N_9637);
nor U10811 (N_10811,N_10444,N_9498);
or U10812 (N_10812,N_9955,N_9379);
nand U10813 (N_10813,N_9634,N_9168);
or U10814 (N_10814,N_9117,N_9224);
xnor U10815 (N_10815,N_10463,N_9830);
and U10816 (N_10816,N_9290,N_9213);
or U10817 (N_10817,N_9861,N_9236);
nor U10818 (N_10818,N_10097,N_9736);
nor U10819 (N_10819,N_10432,N_9883);
xnor U10820 (N_10820,N_9508,N_9608);
nor U10821 (N_10821,N_9503,N_10260);
and U10822 (N_10822,N_9868,N_9745);
or U10823 (N_10823,N_9848,N_9775);
nor U10824 (N_10824,N_9946,N_9803);
xnor U10825 (N_10825,N_9983,N_9255);
or U10826 (N_10826,N_10300,N_9010);
xor U10827 (N_10827,N_9055,N_9818);
and U10828 (N_10828,N_10018,N_9014);
and U10829 (N_10829,N_9298,N_10359);
and U10830 (N_10830,N_9071,N_9545);
nand U10831 (N_10831,N_10014,N_9235);
xnor U10832 (N_10832,N_9193,N_9217);
and U10833 (N_10833,N_9725,N_9008);
xnor U10834 (N_10834,N_9738,N_10240);
xnor U10835 (N_10835,N_9988,N_9941);
nand U10836 (N_10836,N_9227,N_10307);
nor U10837 (N_10837,N_10384,N_10004);
nor U10838 (N_10838,N_10382,N_10428);
nor U10839 (N_10839,N_9929,N_10469);
xnor U10840 (N_10840,N_10415,N_9917);
nor U10841 (N_10841,N_9952,N_9799);
or U10842 (N_10842,N_9915,N_10373);
and U10843 (N_10843,N_9469,N_9833);
or U10844 (N_10844,N_10238,N_9271);
nand U10845 (N_10845,N_10051,N_9671);
xor U10846 (N_10846,N_9476,N_10386);
xor U10847 (N_10847,N_9816,N_9743);
nor U10848 (N_10848,N_10254,N_9281);
or U10849 (N_10849,N_9715,N_10342);
nand U10850 (N_10850,N_9448,N_9319);
and U10851 (N_10851,N_9852,N_9318);
and U10852 (N_10852,N_9673,N_10345);
nor U10853 (N_10853,N_10375,N_9820);
and U10854 (N_10854,N_9342,N_9049);
nor U10855 (N_10855,N_10367,N_9035);
nor U10856 (N_10856,N_9928,N_9525);
nor U10857 (N_10857,N_9103,N_9857);
or U10858 (N_10858,N_9447,N_10094);
xnor U10859 (N_10859,N_9858,N_9675);
and U10860 (N_10860,N_9189,N_9894);
and U10861 (N_10861,N_9837,N_9454);
nand U10862 (N_10862,N_9471,N_9999);
nand U10863 (N_10863,N_9956,N_9616);
xnor U10864 (N_10864,N_10017,N_9597);
nor U10865 (N_10865,N_9110,N_9399);
and U10866 (N_10866,N_9154,N_9344);
or U10867 (N_10867,N_10438,N_10325);
or U10868 (N_10868,N_9274,N_10100);
or U10869 (N_10869,N_9238,N_10453);
nor U10870 (N_10870,N_9054,N_9889);
xor U10871 (N_10871,N_10191,N_9629);
nor U10872 (N_10872,N_10123,N_9264);
nand U10873 (N_10873,N_9947,N_9627);
xnor U10874 (N_10874,N_9265,N_10072);
nor U10875 (N_10875,N_10085,N_9653);
xnor U10876 (N_10876,N_9006,N_9276);
and U10877 (N_10877,N_9310,N_9300);
or U10878 (N_10878,N_10016,N_9152);
and U10879 (N_10879,N_9850,N_9586);
and U10880 (N_10880,N_10233,N_9485);
and U10881 (N_10881,N_9196,N_9699);
xor U10882 (N_10882,N_9155,N_10033);
xor U10883 (N_10883,N_10381,N_9139);
xnor U10884 (N_10884,N_9347,N_9050);
or U10885 (N_10885,N_9216,N_10205);
nand U10886 (N_10886,N_10413,N_10451);
or U10887 (N_10887,N_9307,N_9757);
nand U10888 (N_10888,N_9872,N_9479);
or U10889 (N_10889,N_9292,N_9386);
xnor U10890 (N_10890,N_10201,N_9689);
and U10891 (N_10891,N_10256,N_9631);
xnor U10892 (N_10892,N_10303,N_9442);
xor U10893 (N_10893,N_9944,N_9733);
nand U10894 (N_10894,N_9077,N_9707);
xor U10895 (N_10895,N_9178,N_9244);
xor U10896 (N_10896,N_9710,N_10387);
nand U10897 (N_10897,N_9577,N_10498);
nand U10898 (N_10898,N_9897,N_9039);
xnor U10899 (N_10899,N_9996,N_9506);
xor U10900 (N_10900,N_9912,N_9534);
nor U10901 (N_10901,N_10299,N_9666);
nand U10902 (N_10902,N_10290,N_9851);
nor U10903 (N_10903,N_9080,N_9878);
or U10904 (N_10904,N_9769,N_9328);
nor U10905 (N_10905,N_9930,N_9524);
and U10906 (N_10906,N_9403,N_9903);
and U10907 (N_10907,N_9484,N_9434);
and U10908 (N_10908,N_9149,N_10336);
or U10909 (N_10909,N_10360,N_10292);
xor U10910 (N_10910,N_10176,N_9024);
and U10911 (N_10911,N_9409,N_10098);
xor U10912 (N_10912,N_9102,N_9279);
and U10913 (N_10913,N_9520,N_9240);
nor U10914 (N_10914,N_9560,N_9834);
nand U10915 (N_10915,N_9326,N_9989);
and U10916 (N_10916,N_10366,N_10363);
or U10917 (N_10917,N_9530,N_9581);
nand U10918 (N_10918,N_9142,N_9395);
or U10919 (N_10919,N_9585,N_9225);
and U10920 (N_10920,N_9190,N_9977);
xnor U10921 (N_10921,N_9679,N_9337);
or U10922 (N_10922,N_9364,N_9793);
and U10923 (N_10923,N_10347,N_9997);
nor U10924 (N_10924,N_9043,N_9836);
or U10925 (N_10925,N_10253,N_9839);
nor U10926 (N_10926,N_10156,N_9644);
nand U10927 (N_10927,N_10338,N_9378);
xnor U10928 (N_10928,N_9367,N_10322);
and U10929 (N_10929,N_9500,N_9986);
and U10930 (N_10930,N_9079,N_9118);
and U10931 (N_10931,N_9084,N_9808);
and U10932 (N_10932,N_9011,N_10372);
nand U10933 (N_10933,N_9735,N_10071);
or U10934 (N_10934,N_10236,N_10291);
xnor U10935 (N_10935,N_9717,N_9048);
nor U10936 (N_10936,N_9992,N_10152);
xnor U10937 (N_10937,N_9970,N_9829);
nand U10938 (N_10938,N_9533,N_9677);
xnor U10939 (N_10939,N_9759,N_10277);
xor U10940 (N_10940,N_9052,N_9548);
or U10941 (N_10941,N_9293,N_10422);
xnor U10942 (N_10942,N_10177,N_9350);
nor U10943 (N_10943,N_9191,N_10180);
xnor U10944 (N_10944,N_9734,N_9483);
and U10945 (N_10945,N_9173,N_9890);
and U10946 (N_10946,N_10047,N_9918);
or U10947 (N_10947,N_9574,N_9208);
nor U10948 (N_10948,N_9435,N_9596);
nor U10949 (N_10949,N_9115,N_9884);
nand U10950 (N_10950,N_9020,N_9180);
and U10951 (N_10951,N_9993,N_10148);
or U10952 (N_10952,N_9340,N_9849);
nand U10953 (N_10953,N_10147,N_9972);
nand U10954 (N_10954,N_9611,N_9797);
and U10955 (N_10955,N_9538,N_9089);
nor U10956 (N_10956,N_9555,N_9802);
nor U10957 (N_10957,N_10003,N_9704);
or U10958 (N_10958,N_9460,N_9382);
nor U10959 (N_10959,N_9222,N_10294);
nand U10960 (N_10960,N_10467,N_9206);
nand U10961 (N_10961,N_10488,N_9773);
and U10962 (N_10962,N_10362,N_9028);
or U10963 (N_10963,N_9939,N_10000);
nand U10964 (N_10964,N_9199,N_9719);
or U10965 (N_10965,N_10450,N_9285);
nand U10966 (N_10966,N_9277,N_9101);
nand U10967 (N_10967,N_9174,N_9723);
nor U10968 (N_10968,N_10249,N_9427);
and U10969 (N_10969,N_9253,N_10344);
or U10970 (N_10970,N_10186,N_9076);
and U10971 (N_10971,N_9175,N_9376);
nand U10972 (N_10972,N_10060,N_9674);
and U10973 (N_10973,N_9599,N_10084);
or U10974 (N_10974,N_9964,N_9243);
and U10975 (N_10975,N_9845,N_9444);
nand U10976 (N_10976,N_9953,N_9692);
and U10977 (N_10977,N_9067,N_10462);
or U10978 (N_10978,N_9234,N_9681);
xor U10979 (N_10979,N_9749,N_9068);
xnor U10980 (N_10980,N_9004,N_9355);
xnor U10981 (N_10981,N_9422,N_9287);
nand U10982 (N_10982,N_10460,N_10067);
and U10983 (N_10983,N_9951,N_10323);
xnor U10984 (N_10984,N_9156,N_10289);
xnor U10985 (N_10985,N_10005,N_9258);
xor U10986 (N_10986,N_9252,N_10311);
nand U10987 (N_10987,N_10392,N_9995);
nand U10988 (N_10988,N_9562,N_10437);
or U10989 (N_10989,N_9875,N_9531);
or U10990 (N_10990,N_9212,N_10308);
xor U10991 (N_10991,N_10497,N_9827);
or U10992 (N_10992,N_9478,N_9924);
nand U10993 (N_10993,N_10037,N_9472);
or U10994 (N_10994,N_10332,N_9384);
xnor U10995 (N_10995,N_9419,N_10473);
nand U10996 (N_10996,N_9261,N_9402);
nand U10997 (N_10997,N_9183,N_10443);
or U10998 (N_10998,N_10418,N_9380);
or U10999 (N_10999,N_9275,N_9027);
nor U11000 (N_11000,N_9979,N_10122);
and U11001 (N_11001,N_9959,N_9649);
nand U11002 (N_11002,N_9579,N_9251);
xnor U11003 (N_11003,N_9751,N_10082);
nand U11004 (N_11004,N_10459,N_10419);
and U11005 (N_11005,N_9455,N_10109);
or U11006 (N_11006,N_9491,N_9312);
nand U11007 (N_11007,N_9641,N_9923);
nand U11008 (N_11008,N_10063,N_10150);
xnor U11009 (N_11009,N_9823,N_9544);
or U11010 (N_11010,N_9044,N_9160);
nand U11011 (N_11011,N_10102,N_9229);
nor U11012 (N_11012,N_9898,N_9638);
or U11013 (N_11013,N_10171,N_9474);
xor U11014 (N_11014,N_10203,N_10007);
nand U11015 (N_11015,N_9002,N_10138);
and U11016 (N_11016,N_9790,N_9138);
and U11017 (N_11017,N_9921,N_9007);
xnor U11018 (N_11018,N_10227,N_9621);
nand U11019 (N_11019,N_10310,N_9980);
xnor U11020 (N_11020,N_9302,N_10283);
or U11021 (N_11021,N_9104,N_9591);
nor U11022 (N_11022,N_9094,N_9750);
or U11023 (N_11023,N_9015,N_10391);
and U11024 (N_11024,N_9066,N_9301);
and U11025 (N_11025,N_9200,N_10483);
and U11026 (N_11026,N_9171,N_10410);
nand U11027 (N_11027,N_9182,N_9387);
or U11028 (N_11028,N_10088,N_9781);
nor U11029 (N_11029,N_10295,N_9095);
or U11030 (N_11030,N_9239,N_9948);
xnor U11031 (N_11031,N_9025,N_9120);
nor U11032 (N_11032,N_9642,N_9284);
or U11033 (N_11033,N_9726,N_9940);
nand U11034 (N_11034,N_9146,N_9558);
nand U11035 (N_11035,N_10237,N_9130);
nand U11036 (N_11036,N_9204,N_9249);
nand U11037 (N_11037,N_9459,N_9741);
xnor U11038 (N_11038,N_10111,N_9732);
and U11039 (N_11039,N_9510,N_9134);
xnor U11040 (N_11040,N_9910,N_9566);
and U11041 (N_11041,N_10305,N_10404);
nor U11042 (N_11042,N_10061,N_9267);
and U11043 (N_11043,N_10315,N_9632);
or U11044 (N_11044,N_9322,N_9737);
nand U11045 (N_11045,N_10108,N_9499);
nand U11046 (N_11046,N_9408,N_10335);
nand U11047 (N_11047,N_9205,N_10454);
xor U11048 (N_11048,N_9511,N_9900);
xnor U11049 (N_11049,N_9765,N_9488);
nor U11050 (N_11050,N_9652,N_9470);
nor U11051 (N_11051,N_9394,N_9896);
and U11052 (N_11052,N_9330,N_9557);
nand U11053 (N_11053,N_9362,N_10252);
or U11054 (N_11054,N_9526,N_10427);
or U11055 (N_11055,N_10378,N_9242);
and U11056 (N_11056,N_9361,N_9731);
and U11057 (N_11057,N_10293,N_9676);
nand U11058 (N_11058,N_9373,N_9390);
nand U11059 (N_11059,N_10045,N_10272);
nor U11060 (N_11060,N_9418,N_9456);
nand U11061 (N_11061,N_9372,N_9294);
xor U11062 (N_11062,N_9718,N_10439);
and U11063 (N_11063,N_10284,N_10478);
nand U11064 (N_11064,N_9099,N_9032);
xor U11065 (N_11065,N_9237,N_9817);
nand U11066 (N_11066,N_9431,N_9578);
xor U11067 (N_11067,N_9584,N_10214);
nor U11068 (N_11068,N_9891,N_10081);
or U11069 (N_11069,N_9144,N_10128);
nand U11070 (N_11070,N_10494,N_10174);
and U11071 (N_11071,N_10206,N_9003);
xnor U11072 (N_11072,N_10390,N_9439);
and U11073 (N_11073,N_9796,N_9061);
and U11074 (N_11074,N_10270,N_9556);
or U11075 (N_11075,N_10466,N_10167);
nand U11076 (N_11076,N_10273,N_10340);
and U11077 (N_11077,N_9901,N_10208);
or U11078 (N_11078,N_9696,N_9374);
and U11079 (N_11079,N_9648,N_9575);
xnor U11080 (N_11080,N_9863,N_9822);
xor U11081 (N_11081,N_9341,N_10134);
xnor U11082 (N_11082,N_9922,N_10440);
nor U11083 (N_11083,N_9428,N_9873);
or U11084 (N_11084,N_10472,N_10074);
xnor U11085 (N_11085,N_10477,N_10197);
nand U11086 (N_11086,N_9877,N_9166);
xor U11087 (N_11087,N_9440,N_9167);
nor U11088 (N_11088,N_10064,N_9636);
nor U11089 (N_11089,N_9131,N_9339);
nor U11090 (N_11090,N_9987,N_9452);
xor U11091 (N_11091,N_9038,N_9788);
nor U11092 (N_11092,N_9018,N_9074);
and U11093 (N_11093,N_9693,N_9494);
or U11094 (N_11094,N_9416,N_9270);
nand U11095 (N_11095,N_9346,N_10115);
or U11096 (N_11096,N_10058,N_10024);
nand U11097 (N_11097,N_10154,N_10481);
and U11098 (N_11098,N_9664,N_9058);
and U11099 (N_11099,N_9064,N_10458);
nor U11100 (N_11100,N_9658,N_9124);
nand U11101 (N_11101,N_10337,N_10423);
xnor U11102 (N_11102,N_9159,N_10143);
xor U11103 (N_11103,N_9778,N_10189);
or U11104 (N_11104,N_9595,N_10471);
nor U11105 (N_11105,N_9388,N_10251);
nor U11106 (N_11106,N_9974,N_10160);
nand U11107 (N_11107,N_9060,N_10190);
and U11108 (N_11108,N_10090,N_9088);
nand U11109 (N_11109,N_9966,N_9304);
or U11110 (N_11110,N_10436,N_10318);
and U11111 (N_11111,N_9780,N_10012);
and U11112 (N_11112,N_9528,N_9876);
or U11113 (N_11113,N_10002,N_9214);
nor U11114 (N_11114,N_9625,N_10395);
xnor U11115 (N_11115,N_10070,N_10113);
or U11116 (N_11116,N_9069,N_9529);
nor U11117 (N_11117,N_9259,N_9949);
xor U11118 (N_11118,N_10001,N_9268);
nand U11119 (N_11119,N_9565,N_10199);
or U11120 (N_11120,N_10219,N_9543);
nand U11121 (N_11121,N_10163,N_9042);
or U11122 (N_11122,N_9645,N_9914);
or U11123 (N_11123,N_9308,N_9975);
and U11124 (N_11124,N_9814,N_9713);
nor U11125 (N_11125,N_9712,N_9005);
nor U11126 (N_11126,N_9400,N_9466);
or U11127 (N_11127,N_9812,N_10125);
xnor U11128 (N_11128,N_9357,N_10265);
or U11129 (N_11129,N_9926,N_9517);
nor U11130 (N_11130,N_9201,N_10130);
and U11131 (N_11131,N_9385,N_9795);
nand U11132 (N_11132,N_10304,N_9662);
nor U11133 (N_11133,N_9248,N_9392);
nand U11134 (N_11134,N_9855,N_9630);
nor U11135 (N_11135,N_10247,N_9552);
nand U11136 (N_11136,N_10159,N_9153);
and U11137 (N_11137,N_10184,N_10035);
or U11138 (N_11138,N_10144,N_9700);
nand U11139 (N_11139,N_9758,N_9207);
xor U11140 (N_11140,N_9311,N_10158);
or U11141 (N_11141,N_10420,N_9815);
nor U11142 (N_11142,N_10389,N_9030);
nor U11143 (N_11143,N_9497,N_9651);
xor U11144 (N_11144,N_9887,N_9937);
xor U11145 (N_11145,N_10492,N_9862);
nand U11146 (N_11146,N_10402,N_9619);
and U11147 (N_11147,N_9092,N_9684);
and U11148 (N_11148,N_9613,N_9295);
xnor U11149 (N_11149,N_9888,N_9622);
or U11150 (N_11150,N_10231,N_10334);
and U11151 (N_11151,N_9540,N_10321);
xnor U11152 (N_11152,N_10129,N_9874);
nand U11153 (N_11153,N_9711,N_9991);
and U11154 (N_11154,N_9158,N_10216);
nor U11155 (N_11155,N_10173,N_9801);
or U11156 (N_11156,N_9145,N_10137);
or U11157 (N_11157,N_9133,N_9806);
nand U11158 (N_11158,N_10329,N_10053);
xnor U11159 (N_11159,N_9687,N_9841);
xor U11160 (N_11160,N_9885,N_9592);
xor U11161 (N_11161,N_10153,N_10348);
xor U11162 (N_11162,N_9931,N_10013);
xor U11163 (N_11163,N_10075,N_9588);
and U11164 (N_11164,N_9404,N_9057);
and U11165 (N_11165,N_9272,N_9665);
nand U11166 (N_11166,N_9147,N_9702);
nand U11167 (N_11167,N_9551,N_9604);
and U11168 (N_11168,N_9618,N_10297);
nor U11169 (N_11169,N_10204,N_9034);
or U11170 (N_11170,N_9954,N_9223);
and U11171 (N_11171,N_9203,N_9610);
or U11172 (N_11172,N_10449,N_10023);
xnor U11173 (N_11173,N_9825,N_10306);
and U11174 (N_11174,N_9262,N_9381);
or U11175 (N_11175,N_10266,N_9468);
nand U11176 (N_11176,N_9332,N_10408);
nand U11177 (N_11177,N_10010,N_10434);
nand U11178 (N_11178,N_10038,N_9950);
and U11179 (N_11179,N_9879,N_9377);
nor U11180 (N_11180,N_10009,N_9192);
or U11181 (N_11181,N_9096,N_10194);
or U11182 (N_11182,N_9366,N_9976);
nor U11183 (N_11183,N_9809,N_10287);
or U11184 (N_11184,N_9001,N_9023);
or U11185 (N_11185,N_9132,N_9389);
nand U11186 (N_11186,N_10210,N_9605);
or U11187 (N_11187,N_10114,N_10198);
xnor U11188 (N_11188,N_9177,N_9536);
nor U11189 (N_11189,N_10217,N_10161);
or U11190 (N_11190,N_9908,N_9882);
xnor U11191 (N_11191,N_10352,N_10193);
and U11192 (N_11192,N_9563,N_9504);
nor U11193 (N_11193,N_9465,N_9129);
nor U11194 (N_11194,N_9309,N_10282);
xnor U11195 (N_11195,N_9197,N_10181);
nor U11196 (N_11196,N_9121,N_9016);
xor U11197 (N_11197,N_9593,N_10376);
nor U11198 (N_11198,N_9411,N_9059);
nand U11199 (N_11199,N_9356,N_9840);
or U11200 (N_11200,N_10145,N_9371);
and U11201 (N_11201,N_10232,N_9317);
or U11202 (N_11202,N_9125,N_9865);
and U11203 (N_11203,N_10495,N_10486);
nand U11204 (N_11204,N_9254,N_10050);
and U11205 (N_11205,N_9358,N_10093);
and U11206 (N_11206,N_10281,N_9114);
xor U11207 (N_11207,N_9602,N_10155);
and U11208 (N_11208,N_9141,N_9090);
and U11209 (N_11209,N_9495,N_10179);
xnor U11210 (N_11210,N_9580,N_9549);
nor U11211 (N_11211,N_9842,N_10015);
xnor U11212 (N_11212,N_10042,N_9655);
nor U11213 (N_11213,N_9756,N_9895);
nor U11214 (N_11214,N_10057,N_9286);
nand U11215 (N_11215,N_9269,N_10257);
or U11216 (N_11216,N_9151,N_9744);
nor U11217 (N_11217,N_9784,N_9761);
nand U11218 (N_11218,N_9022,N_9705);
xor U11219 (N_11219,N_9126,N_9639);
nor U11220 (N_11220,N_10355,N_9289);
and U11221 (N_11221,N_9965,N_10026);
nand U11222 (N_11222,N_10164,N_9250);
nand U11223 (N_11223,N_10069,N_9496);
xor U11224 (N_11224,N_9100,N_9327);
and U11225 (N_11225,N_9335,N_10397);
nor U11226 (N_11226,N_10493,N_10107);
or U11227 (N_11227,N_9108,N_10243);
and U11228 (N_11228,N_10225,N_10046);
and U11229 (N_11229,N_9441,N_9083);
or U11230 (N_11230,N_9351,N_9359);
nand U11231 (N_11231,N_9522,N_10092);
or U11232 (N_11232,N_9527,N_10099);
xor U11233 (N_11233,N_10370,N_10116);
nand U11234 (N_11234,N_9299,N_10149);
and U11235 (N_11235,N_10278,N_10456);
nor U11236 (N_11236,N_9368,N_9698);
xor U11237 (N_11237,N_9401,N_10285);
nor U11238 (N_11238,N_9296,N_10101);
and U11239 (N_11239,N_9961,N_9746);
nand U11240 (N_11240,N_9614,N_9554);
nand U11241 (N_11241,N_9405,N_10136);
nor U11242 (N_11242,N_9087,N_10358);
and U11243 (N_11243,N_9594,N_9467);
and U11244 (N_11244,N_10040,N_9345);
or U11245 (N_11245,N_9306,N_10388);
nor U11246 (N_11246,N_9968,N_9247);
nand U11247 (N_11247,N_9082,N_9785);
nand U11248 (N_11248,N_9211,N_9143);
nor U11249 (N_11249,N_10479,N_9221);
nor U11250 (N_11250,N_9750,N_9438);
nand U11251 (N_11251,N_10218,N_9473);
xnor U11252 (N_11252,N_9420,N_9535);
nand U11253 (N_11253,N_10400,N_9341);
and U11254 (N_11254,N_9911,N_9226);
and U11255 (N_11255,N_9744,N_10373);
and U11256 (N_11256,N_9245,N_9771);
nand U11257 (N_11257,N_9569,N_10127);
or U11258 (N_11258,N_9145,N_9194);
nor U11259 (N_11259,N_9428,N_9389);
or U11260 (N_11260,N_9638,N_10230);
xnor U11261 (N_11261,N_9264,N_10313);
nand U11262 (N_11262,N_10167,N_9119);
nor U11263 (N_11263,N_10426,N_9297);
or U11264 (N_11264,N_9934,N_9003);
nand U11265 (N_11265,N_10269,N_9074);
nand U11266 (N_11266,N_10136,N_9958);
xor U11267 (N_11267,N_9867,N_9759);
xnor U11268 (N_11268,N_9792,N_9303);
nor U11269 (N_11269,N_9171,N_9591);
nand U11270 (N_11270,N_9411,N_9732);
or U11271 (N_11271,N_10391,N_10482);
nor U11272 (N_11272,N_10441,N_9907);
nor U11273 (N_11273,N_10092,N_9303);
nand U11274 (N_11274,N_9475,N_9085);
xor U11275 (N_11275,N_10400,N_9444);
and U11276 (N_11276,N_10306,N_9733);
or U11277 (N_11277,N_10487,N_9170);
xnor U11278 (N_11278,N_9701,N_10270);
or U11279 (N_11279,N_10279,N_10094);
nor U11280 (N_11280,N_9402,N_9471);
nor U11281 (N_11281,N_9114,N_9985);
nand U11282 (N_11282,N_9125,N_9193);
nand U11283 (N_11283,N_9314,N_9043);
and U11284 (N_11284,N_9289,N_10313);
or U11285 (N_11285,N_9974,N_9797);
nand U11286 (N_11286,N_9249,N_10358);
or U11287 (N_11287,N_9887,N_9636);
xnor U11288 (N_11288,N_10158,N_10296);
nor U11289 (N_11289,N_9758,N_9660);
or U11290 (N_11290,N_9890,N_10327);
nor U11291 (N_11291,N_9924,N_10426);
or U11292 (N_11292,N_9815,N_9395);
nand U11293 (N_11293,N_9409,N_9267);
or U11294 (N_11294,N_10394,N_9964);
nor U11295 (N_11295,N_9782,N_10317);
xnor U11296 (N_11296,N_9887,N_9833);
nor U11297 (N_11297,N_9409,N_10100);
nor U11298 (N_11298,N_9604,N_9866);
and U11299 (N_11299,N_10411,N_10056);
and U11300 (N_11300,N_9419,N_10138);
or U11301 (N_11301,N_9686,N_10390);
or U11302 (N_11302,N_9522,N_9176);
xor U11303 (N_11303,N_10448,N_9950);
or U11304 (N_11304,N_10096,N_10306);
or U11305 (N_11305,N_9992,N_9394);
or U11306 (N_11306,N_9586,N_9879);
xor U11307 (N_11307,N_10372,N_10469);
nand U11308 (N_11308,N_10395,N_9027);
or U11309 (N_11309,N_9064,N_9822);
and U11310 (N_11310,N_9873,N_10247);
or U11311 (N_11311,N_9877,N_9775);
xor U11312 (N_11312,N_9698,N_9407);
nor U11313 (N_11313,N_9805,N_9500);
and U11314 (N_11314,N_10105,N_9781);
or U11315 (N_11315,N_9490,N_10099);
nand U11316 (N_11316,N_10261,N_9015);
or U11317 (N_11317,N_10009,N_9758);
nor U11318 (N_11318,N_9993,N_10354);
or U11319 (N_11319,N_10132,N_9750);
and U11320 (N_11320,N_10137,N_10245);
or U11321 (N_11321,N_9734,N_9954);
nand U11322 (N_11322,N_10055,N_10194);
nand U11323 (N_11323,N_9535,N_9817);
nand U11324 (N_11324,N_10059,N_9217);
and U11325 (N_11325,N_9428,N_9003);
and U11326 (N_11326,N_10167,N_9649);
nand U11327 (N_11327,N_9700,N_9776);
xnor U11328 (N_11328,N_9319,N_9810);
nand U11329 (N_11329,N_10453,N_10478);
nor U11330 (N_11330,N_9730,N_9820);
nor U11331 (N_11331,N_9196,N_9322);
or U11332 (N_11332,N_9313,N_9629);
and U11333 (N_11333,N_9417,N_10124);
nand U11334 (N_11334,N_10236,N_9981);
xor U11335 (N_11335,N_10001,N_9830);
or U11336 (N_11336,N_9836,N_9320);
nor U11337 (N_11337,N_9418,N_9219);
or U11338 (N_11338,N_9341,N_9400);
nor U11339 (N_11339,N_9158,N_10289);
nand U11340 (N_11340,N_9021,N_9619);
nand U11341 (N_11341,N_9877,N_10092);
xor U11342 (N_11342,N_10419,N_9702);
and U11343 (N_11343,N_10261,N_9349);
or U11344 (N_11344,N_9457,N_9856);
xnor U11345 (N_11345,N_9402,N_9177);
xor U11346 (N_11346,N_9347,N_9036);
xor U11347 (N_11347,N_9146,N_10375);
xnor U11348 (N_11348,N_10080,N_9466);
and U11349 (N_11349,N_10160,N_9854);
and U11350 (N_11350,N_9724,N_9308);
xnor U11351 (N_11351,N_9499,N_9594);
and U11352 (N_11352,N_9098,N_9705);
xnor U11353 (N_11353,N_9410,N_9002);
nand U11354 (N_11354,N_9032,N_10392);
xor U11355 (N_11355,N_9816,N_10430);
or U11356 (N_11356,N_9422,N_9340);
nor U11357 (N_11357,N_10389,N_9303);
nor U11358 (N_11358,N_9222,N_10119);
xor U11359 (N_11359,N_9431,N_9831);
and U11360 (N_11360,N_9960,N_9861);
nor U11361 (N_11361,N_9975,N_10155);
or U11362 (N_11362,N_9281,N_9194);
xnor U11363 (N_11363,N_10257,N_10041);
or U11364 (N_11364,N_9016,N_9772);
or U11365 (N_11365,N_9704,N_10373);
nor U11366 (N_11366,N_10311,N_9163);
nand U11367 (N_11367,N_9873,N_9565);
and U11368 (N_11368,N_9992,N_10430);
and U11369 (N_11369,N_9164,N_10474);
nor U11370 (N_11370,N_9507,N_10488);
nor U11371 (N_11371,N_9078,N_9747);
xnor U11372 (N_11372,N_9481,N_9415);
or U11373 (N_11373,N_9532,N_9949);
and U11374 (N_11374,N_9320,N_9087);
nand U11375 (N_11375,N_9169,N_9786);
nand U11376 (N_11376,N_9541,N_10195);
nand U11377 (N_11377,N_9009,N_10050);
or U11378 (N_11378,N_9019,N_10010);
or U11379 (N_11379,N_9136,N_10155);
and U11380 (N_11380,N_9379,N_9350);
nand U11381 (N_11381,N_9285,N_9026);
xnor U11382 (N_11382,N_10251,N_9330);
or U11383 (N_11383,N_10128,N_10465);
xnor U11384 (N_11384,N_9524,N_9943);
and U11385 (N_11385,N_9552,N_9153);
xnor U11386 (N_11386,N_10310,N_9072);
xor U11387 (N_11387,N_9463,N_9625);
xnor U11388 (N_11388,N_9835,N_9220);
xnor U11389 (N_11389,N_10032,N_10456);
xnor U11390 (N_11390,N_9920,N_10139);
nand U11391 (N_11391,N_9661,N_9047);
and U11392 (N_11392,N_9199,N_10212);
xor U11393 (N_11393,N_9595,N_9216);
nand U11394 (N_11394,N_10284,N_10170);
nand U11395 (N_11395,N_10487,N_9800);
and U11396 (N_11396,N_9865,N_9204);
and U11397 (N_11397,N_10006,N_9313);
and U11398 (N_11398,N_9861,N_10355);
and U11399 (N_11399,N_9500,N_9816);
or U11400 (N_11400,N_9811,N_9300);
xnor U11401 (N_11401,N_9586,N_9002);
nor U11402 (N_11402,N_9244,N_10486);
xor U11403 (N_11403,N_10156,N_10472);
nor U11404 (N_11404,N_9909,N_9499);
nand U11405 (N_11405,N_9678,N_10040);
nand U11406 (N_11406,N_10473,N_10072);
xnor U11407 (N_11407,N_9026,N_9483);
nand U11408 (N_11408,N_10132,N_9564);
and U11409 (N_11409,N_9218,N_9050);
and U11410 (N_11410,N_10362,N_9330);
nor U11411 (N_11411,N_9946,N_9565);
nor U11412 (N_11412,N_10260,N_9106);
nand U11413 (N_11413,N_9842,N_9161);
nand U11414 (N_11414,N_9853,N_9878);
or U11415 (N_11415,N_9894,N_10185);
and U11416 (N_11416,N_9492,N_9692);
nor U11417 (N_11417,N_9703,N_9997);
and U11418 (N_11418,N_9390,N_10355);
and U11419 (N_11419,N_9439,N_9269);
xor U11420 (N_11420,N_9119,N_9695);
and U11421 (N_11421,N_10180,N_9332);
xnor U11422 (N_11422,N_9395,N_9655);
xor U11423 (N_11423,N_10230,N_10036);
nor U11424 (N_11424,N_9781,N_9509);
and U11425 (N_11425,N_10176,N_9440);
nand U11426 (N_11426,N_9559,N_10495);
nor U11427 (N_11427,N_9537,N_9381);
nand U11428 (N_11428,N_9586,N_10472);
xnor U11429 (N_11429,N_9807,N_10091);
nor U11430 (N_11430,N_9749,N_10197);
and U11431 (N_11431,N_9370,N_9349);
nor U11432 (N_11432,N_9758,N_9124);
xor U11433 (N_11433,N_9347,N_9231);
xor U11434 (N_11434,N_9189,N_10225);
nand U11435 (N_11435,N_10467,N_10402);
nand U11436 (N_11436,N_9508,N_9075);
or U11437 (N_11437,N_10314,N_10390);
or U11438 (N_11438,N_9425,N_10249);
and U11439 (N_11439,N_10234,N_10138);
nand U11440 (N_11440,N_10280,N_9429);
xor U11441 (N_11441,N_9617,N_9201);
nand U11442 (N_11442,N_9247,N_9582);
xor U11443 (N_11443,N_9687,N_9184);
and U11444 (N_11444,N_9326,N_10275);
nand U11445 (N_11445,N_9454,N_10431);
and U11446 (N_11446,N_9747,N_10466);
nand U11447 (N_11447,N_10164,N_9078);
or U11448 (N_11448,N_9010,N_9822);
and U11449 (N_11449,N_9191,N_9803);
nor U11450 (N_11450,N_9167,N_9040);
xor U11451 (N_11451,N_10402,N_9959);
nand U11452 (N_11452,N_9573,N_9047);
xor U11453 (N_11453,N_9165,N_10135);
and U11454 (N_11454,N_9643,N_10258);
or U11455 (N_11455,N_9274,N_9298);
nor U11456 (N_11456,N_10190,N_9238);
and U11457 (N_11457,N_9379,N_10279);
nor U11458 (N_11458,N_9906,N_10138);
or U11459 (N_11459,N_9175,N_10252);
nand U11460 (N_11460,N_9914,N_9121);
xnor U11461 (N_11461,N_9627,N_10309);
or U11462 (N_11462,N_9935,N_9626);
and U11463 (N_11463,N_9974,N_9951);
and U11464 (N_11464,N_9223,N_10266);
nand U11465 (N_11465,N_10082,N_10498);
nor U11466 (N_11466,N_9137,N_10126);
or U11467 (N_11467,N_9629,N_9953);
or U11468 (N_11468,N_9582,N_10010);
nor U11469 (N_11469,N_9715,N_10099);
xor U11470 (N_11470,N_10295,N_10441);
or U11471 (N_11471,N_10309,N_9258);
nand U11472 (N_11472,N_9475,N_9136);
or U11473 (N_11473,N_10268,N_9433);
and U11474 (N_11474,N_9435,N_9494);
xnor U11475 (N_11475,N_10160,N_9679);
nand U11476 (N_11476,N_10415,N_9309);
nand U11477 (N_11477,N_9396,N_9976);
or U11478 (N_11478,N_9005,N_9914);
xnor U11479 (N_11479,N_9194,N_9344);
xor U11480 (N_11480,N_9472,N_9958);
or U11481 (N_11481,N_10239,N_9933);
nand U11482 (N_11482,N_9042,N_9316);
or U11483 (N_11483,N_9622,N_9864);
and U11484 (N_11484,N_9901,N_9630);
nand U11485 (N_11485,N_10372,N_10383);
nor U11486 (N_11486,N_9508,N_10354);
and U11487 (N_11487,N_9971,N_9287);
xor U11488 (N_11488,N_9680,N_10327);
xnor U11489 (N_11489,N_9764,N_9353);
xnor U11490 (N_11490,N_10153,N_10170);
nor U11491 (N_11491,N_9413,N_9393);
nand U11492 (N_11492,N_9702,N_9927);
xor U11493 (N_11493,N_10320,N_9974);
xor U11494 (N_11494,N_9388,N_9893);
xor U11495 (N_11495,N_10185,N_10492);
and U11496 (N_11496,N_10173,N_9067);
nor U11497 (N_11497,N_9525,N_10093);
or U11498 (N_11498,N_9346,N_9183);
nand U11499 (N_11499,N_9087,N_9639);
nor U11500 (N_11500,N_9245,N_9435);
xor U11501 (N_11501,N_9775,N_9125);
xnor U11502 (N_11502,N_9129,N_10113);
xnor U11503 (N_11503,N_9192,N_10387);
nand U11504 (N_11504,N_9241,N_9999);
nor U11505 (N_11505,N_9881,N_9923);
nor U11506 (N_11506,N_9041,N_9372);
and U11507 (N_11507,N_10109,N_9823);
nor U11508 (N_11508,N_10295,N_9797);
xnor U11509 (N_11509,N_9420,N_9332);
nand U11510 (N_11510,N_9902,N_9514);
nor U11511 (N_11511,N_10210,N_9519);
nor U11512 (N_11512,N_10408,N_9211);
nand U11513 (N_11513,N_9674,N_9124);
or U11514 (N_11514,N_9118,N_9944);
nand U11515 (N_11515,N_10007,N_9738);
and U11516 (N_11516,N_9621,N_9151);
nand U11517 (N_11517,N_9111,N_9906);
xor U11518 (N_11518,N_9146,N_9549);
and U11519 (N_11519,N_10330,N_10497);
nor U11520 (N_11520,N_10299,N_9984);
nor U11521 (N_11521,N_9502,N_9475);
xor U11522 (N_11522,N_9772,N_9007);
and U11523 (N_11523,N_9835,N_10127);
nand U11524 (N_11524,N_9440,N_9808);
and U11525 (N_11525,N_9112,N_10069);
xnor U11526 (N_11526,N_10342,N_9928);
and U11527 (N_11527,N_10022,N_9249);
or U11528 (N_11528,N_9518,N_9807);
nor U11529 (N_11529,N_10254,N_10293);
nand U11530 (N_11530,N_9384,N_9560);
xnor U11531 (N_11531,N_9287,N_9721);
xor U11532 (N_11532,N_9415,N_10263);
nand U11533 (N_11533,N_10462,N_10144);
and U11534 (N_11534,N_10253,N_10402);
or U11535 (N_11535,N_9448,N_9758);
or U11536 (N_11536,N_10182,N_10199);
xnor U11537 (N_11537,N_10369,N_10364);
or U11538 (N_11538,N_10209,N_9796);
nand U11539 (N_11539,N_9472,N_10115);
and U11540 (N_11540,N_9853,N_10107);
and U11541 (N_11541,N_9851,N_9121);
nand U11542 (N_11542,N_9930,N_9974);
nor U11543 (N_11543,N_9299,N_9885);
or U11544 (N_11544,N_9506,N_9924);
nor U11545 (N_11545,N_10296,N_9292);
and U11546 (N_11546,N_10253,N_9660);
xnor U11547 (N_11547,N_9885,N_9778);
and U11548 (N_11548,N_10045,N_9353);
xnor U11549 (N_11549,N_10322,N_9241);
xor U11550 (N_11550,N_10432,N_9744);
and U11551 (N_11551,N_9470,N_9572);
xor U11552 (N_11552,N_10097,N_9301);
nand U11553 (N_11553,N_9958,N_9554);
or U11554 (N_11554,N_10247,N_9183);
nor U11555 (N_11555,N_9667,N_9531);
nand U11556 (N_11556,N_10402,N_10173);
or U11557 (N_11557,N_9941,N_9722);
nor U11558 (N_11558,N_9674,N_9265);
nor U11559 (N_11559,N_9092,N_9514);
nand U11560 (N_11560,N_9572,N_10066);
nand U11561 (N_11561,N_9571,N_9109);
nor U11562 (N_11562,N_10246,N_9083);
and U11563 (N_11563,N_9671,N_10287);
xnor U11564 (N_11564,N_9935,N_9602);
nor U11565 (N_11565,N_9590,N_10389);
nor U11566 (N_11566,N_9815,N_10310);
nor U11567 (N_11567,N_9223,N_9216);
and U11568 (N_11568,N_10337,N_10035);
or U11569 (N_11569,N_10474,N_10464);
nor U11570 (N_11570,N_9585,N_9061);
and U11571 (N_11571,N_9510,N_9182);
nand U11572 (N_11572,N_10221,N_9961);
nand U11573 (N_11573,N_9979,N_10301);
or U11574 (N_11574,N_9004,N_9673);
or U11575 (N_11575,N_9922,N_9291);
nand U11576 (N_11576,N_9145,N_9439);
xnor U11577 (N_11577,N_10120,N_9565);
nor U11578 (N_11578,N_10365,N_10212);
or U11579 (N_11579,N_9816,N_10306);
and U11580 (N_11580,N_10244,N_9191);
xor U11581 (N_11581,N_9022,N_10002);
and U11582 (N_11582,N_10434,N_10213);
xnor U11583 (N_11583,N_9635,N_9968);
or U11584 (N_11584,N_9106,N_10140);
or U11585 (N_11585,N_10321,N_9916);
nor U11586 (N_11586,N_10144,N_9098);
xor U11587 (N_11587,N_9150,N_9201);
nand U11588 (N_11588,N_10016,N_9326);
xnor U11589 (N_11589,N_10111,N_10060);
xor U11590 (N_11590,N_9114,N_9483);
xor U11591 (N_11591,N_9569,N_9999);
nand U11592 (N_11592,N_9527,N_10199);
and U11593 (N_11593,N_9043,N_9894);
and U11594 (N_11594,N_10313,N_9442);
or U11595 (N_11595,N_9263,N_9959);
and U11596 (N_11596,N_9038,N_10349);
nor U11597 (N_11597,N_10409,N_10312);
and U11598 (N_11598,N_9150,N_9071);
xnor U11599 (N_11599,N_9381,N_9292);
xnor U11600 (N_11600,N_10121,N_10007);
and U11601 (N_11601,N_9471,N_10329);
xnor U11602 (N_11602,N_10275,N_9233);
nor U11603 (N_11603,N_9536,N_10156);
nor U11604 (N_11604,N_9748,N_9325);
nand U11605 (N_11605,N_10409,N_9103);
or U11606 (N_11606,N_9514,N_9297);
nand U11607 (N_11607,N_10133,N_9288);
nand U11608 (N_11608,N_10169,N_10309);
and U11609 (N_11609,N_9158,N_10494);
and U11610 (N_11610,N_9824,N_10349);
and U11611 (N_11611,N_9270,N_9352);
nor U11612 (N_11612,N_9550,N_9561);
xor U11613 (N_11613,N_9722,N_9413);
xor U11614 (N_11614,N_9746,N_9339);
xnor U11615 (N_11615,N_10143,N_10198);
or U11616 (N_11616,N_9045,N_9915);
xnor U11617 (N_11617,N_10472,N_9059);
nand U11618 (N_11618,N_10058,N_9226);
nor U11619 (N_11619,N_10228,N_9689);
or U11620 (N_11620,N_9140,N_10246);
or U11621 (N_11621,N_10328,N_9711);
nand U11622 (N_11622,N_9942,N_9267);
nand U11623 (N_11623,N_10499,N_10092);
and U11624 (N_11624,N_9704,N_10011);
nand U11625 (N_11625,N_10210,N_10208);
xnor U11626 (N_11626,N_10494,N_9777);
nor U11627 (N_11627,N_10403,N_9576);
nand U11628 (N_11628,N_9074,N_9524);
and U11629 (N_11629,N_10135,N_9122);
nand U11630 (N_11630,N_10339,N_10330);
or U11631 (N_11631,N_9844,N_9853);
nor U11632 (N_11632,N_9236,N_9652);
nand U11633 (N_11633,N_9428,N_9417);
and U11634 (N_11634,N_9006,N_9200);
nor U11635 (N_11635,N_9826,N_10035);
nand U11636 (N_11636,N_9344,N_10399);
and U11637 (N_11637,N_9274,N_10004);
or U11638 (N_11638,N_10193,N_10494);
xor U11639 (N_11639,N_9781,N_9443);
and U11640 (N_11640,N_9100,N_9425);
nor U11641 (N_11641,N_9623,N_9756);
nor U11642 (N_11642,N_9131,N_10007);
nor U11643 (N_11643,N_10163,N_9431);
or U11644 (N_11644,N_9465,N_9551);
xnor U11645 (N_11645,N_10111,N_10252);
or U11646 (N_11646,N_9243,N_9038);
xor U11647 (N_11647,N_9492,N_10431);
or U11648 (N_11648,N_9010,N_9343);
nor U11649 (N_11649,N_9788,N_9531);
xnor U11650 (N_11650,N_9384,N_9036);
nor U11651 (N_11651,N_10109,N_9909);
or U11652 (N_11652,N_9124,N_9782);
xnor U11653 (N_11653,N_9421,N_9391);
and U11654 (N_11654,N_9701,N_9879);
or U11655 (N_11655,N_9619,N_10147);
nand U11656 (N_11656,N_10167,N_10278);
or U11657 (N_11657,N_10478,N_9460);
nand U11658 (N_11658,N_10464,N_10277);
nor U11659 (N_11659,N_10493,N_9168);
nand U11660 (N_11660,N_9521,N_9228);
xor U11661 (N_11661,N_9686,N_9811);
nand U11662 (N_11662,N_9763,N_10412);
nor U11663 (N_11663,N_10228,N_9128);
and U11664 (N_11664,N_10393,N_9018);
xor U11665 (N_11665,N_9057,N_9380);
xnor U11666 (N_11666,N_9694,N_9582);
nor U11667 (N_11667,N_9006,N_9460);
nand U11668 (N_11668,N_9910,N_10129);
nand U11669 (N_11669,N_9069,N_9424);
or U11670 (N_11670,N_9260,N_9837);
or U11671 (N_11671,N_9496,N_10204);
nor U11672 (N_11672,N_10022,N_10373);
nor U11673 (N_11673,N_9498,N_9137);
or U11674 (N_11674,N_10369,N_9732);
or U11675 (N_11675,N_9287,N_10253);
nor U11676 (N_11676,N_10318,N_9752);
xnor U11677 (N_11677,N_9096,N_10381);
nand U11678 (N_11678,N_9132,N_9883);
nor U11679 (N_11679,N_9608,N_10340);
nand U11680 (N_11680,N_10386,N_9981);
xor U11681 (N_11681,N_9869,N_9971);
xor U11682 (N_11682,N_9930,N_10236);
xnor U11683 (N_11683,N_10165,N_10182);
nor U11684 (N_11684,N_9350,N_10144);
nor U11685 (N_11685,N_10458,N_9875);
or U11686 (N_11686,N_9354,N_9753);
nand U11687 (N_11687,N_10473,N_10483);
nor U11688 (N_11688,N_10147,N_9145);
nor U11689 (N_11689,N_9228,N_9981);
or U11690 (N_11690,N_9116,N_10274);
xor U11691 (N_11691,N_9113,N_9437);
and U11692 (N_11692,N_9667,N_9783);
nor U11693 (N_11693,N_9339,N_9879);
xnor U11694 (N_11694,N_9766,N_9198);
and U11695 (N_11695,N_9516,N_9386);
nand U11696 (N_11696,N_9127,N_9625);
nand U11697 (N_11697,N_9076,N_9989);
xnor U11698 (N_11698,N_10367,N_10294);
xnor U11699 (N_11699,N_9430,N_9935);
xor U11700 (N_11700,N_10477,N_10029);
nand U11701 (N_11701,N_9610,N_10358);
and U11702 (N_11702,N_10482,N_10006);
nand U11703 (N_11703,N_9927,N_9145);
nand U11704 (N_11704,N_9567,N_10414);
nand U11705 (N_11705,N_9082,N_10416);
or U11706 (N_11706,N_9383,N_9584);
nand U11707 (N_11707,N_10345,N_9282);
xor U11708 (N_11708,N_10457,N_9144);
and U11709 (N_11709,N_9150,N_10079);
nand U11710 (N_11710,N_10147,N_9558);
xnor U11711 (N_11711,N_9366,N_9074);
xnor U11712 (N_11712,N_10189,N_9098);
and U11713 (N_11713,N_9449,N_9041);
or U11714 (N_11714,N_10324,N_9549);
and U11715 (N_11715,N_10423,N_10340);
nand U11716 (N_11716,N_9235,N_10254);
or U11717 (N_11717,N_10427,N_10104);
nor U11718 (N_11718,N_9029,N_9792);
xnor U11719 (N_11719,N_9082,N_9577);
and U11720 (N_11720,N_10398,N_9100);
nand U11721 (N_11721,N_10315,N_9045);
nand U11722 (N_11722,N_9580,N_10276);
and U11723 (N_11723,N_9490,N_10436);
nand U11724 (N_11724,N_9019,N_9470);
xnor U11725 (N_11725,N_10182,N_10432);
or U11726 (N_11726,N_10254,N_10338);
nand U11727 (N_11727,N_9707,N_10472);
and U11728 (N_11728,N_9088,N_9976);
nand U11729 (N_11729,N_10082,N_9586);
nor U11730 (N_11730,N_9778,N_9985);
or U11731 (N_11731,N_10133,N_10120);
nor U11732 (N_11732,N_10123,N_10194);
nand U11733 (N_11733,N_9516,N_10264);
and U11734 (N_11734,N_9300,N_9720);
xor U11735 (N_11735,N_9482,N_9091);
xor U11736 (N_11736,N_9612,N_9935);
nand U11737 (N_11737,N_9069,N_9213);
xor U11738 (N_11738,N_10226,N_10002);
xnor U11739 (N_11739,N_9572,N_9612);
nor U11740 (N_11740,N_9379,N_10360);
nor U11741 (N_11741,N_9836,N_9977);
and U11742 (N_11742,N_10051,N_9468);
and U11743 (N_11743,N_9626,N_9397);
and U11744 (N_11744,N_9730,N_10306);
or U11745 (N_11745,N_9554,N_9921);
nor U11746 (N_11746,N_9812,N_9035);
or U11747 (N_11747,N_9125,N_9369);
nand U11748 (N_11748,N_10146,N_9139);
and U11749 (N_11749,N_9697,N_9849);
or U11750 (N_11750,N_10001,N_9637);
nor U11751 (N_11751,N_9708,N_10119);
or U11752 (N_11752,N_10095,N_9310);
xnor U11753 (N_11753,N_9935,N_9860);
or U11754 (N_11754,N_9186,N_10486);
or U11755 (N_11755,N_9600,N_10287);
or U11756 (N_11756,N_10258,N_9383);
and U11757 (N_11757,N_9722,N_10307);
xor U11758 (N_11758,N_9797,N_9794);
nand U11759 (N_11759,N_9773,N_9227);
xnor U11760 (N_11760,N_9153,N_9802);
xor U11761 (N_11761,N_9643,N_10126);
xor U11762 (N_11762,N_9765,N_9072);
or U11763 (N_11763,N_10205,N_10312);
nand U11764 (N_11764,N_9976,N_9760);
and U11765 (N_11765,N_9350,N_9896);
xnor U11766 (N_11766,N_10328,N_9321);
xnor U11767 (N_11767,N_9097,N_9801);
xnor U11768 (N_11768,N_9621,N_10202);
nand U11769 (N_11769,N_9844,N_9729);
or U11770 (N_11770,N_10405,N_9461);
xor U11771 (N_11771,N_9959,N_9655);
nor U11772 (N_11772,N_10086,N_10429);
nand U11773 (N_11773,N_9751,N_9525);
and U11774 (N_11774,N_9964,N_9952);
and U11775 (N_11775,N_9247,N_9844);
xor U11776 (N_11776,N_9878,N_9004);
nor U11777 (N_11777,N_10306,N_9346);
or U11778 (N_11778,N_10391,N_9848);
nor U11779 (N_11779,N_9069,N_9647);
or U11780 (N_11780,N_10288,N_10425);
nor U11781 (N_11781,N_9300,N_9157);
nor U11782 (N_11782,N_10118,N_9471);
nand U11783 (N_11783,N_10445,N_10161);
xor U11784 (N_11784,N_9202,N_10423);
and U11785 (N_11785,N_10479,N_9266);
xnor U11786 (N_11786,N_9550,N_9016);
and U11787 (N_11787,N_9845,N_9336);
xor U11788 (N_11788,N_10169,N_10099);
and U11789 (N_11789,N_9712,N_9016);
nor U11790 (N_11790,N_10424,N_10306);
nand U11791 (N_11791,N_10270,N_9643);
xnor U11792 (N_11792,N_9784,N_9305);
nand U11793 (N_11793,N_10008,N_10282);
nor U11794 (N_11794,N_9432,N_9671);
nor U11795 (N_11795,N_9732,N_10247);
nand U11796 (N_11796,N_9515,N_9671);
nor U11797 (N_11797,N_9157,N_9395);
nand U11798 (N_11798,N_9280,N_9370);
or U11799 (N_11799,N_10209,N_10199);
xnor U11800 (N_11800,N_9919,N_10234);
and U11801 (N_11801,N_10196,N_10470);
nand U11802 (N_11802,N_10008,N_9823);
xnor U11803 (N_11803,N_9406,N_10287);
and U11804 (N_11804,N_10001,N_9741);
and U11805 (N_11805,N_9019,N_9032);
nor U11806 (N_11806,N_9489,N_10333);
nand U11807 (N_11807,N_9926,N_10327);
nor U11808 (N_11808,N_10228,N_10247);
nand U11809 (N_11809,N_10086,N_9544);
nor U11810 (N_11810,N_9565,N_9385);
or U11811 (N_11811,N_10122,N_9321);
or U11812 (N_11812,N_10430,N_9461);
nor U11813 (N_11813,N_9102,N_10149);
nor U11814 (N_11814,N_9883,N_9330);
xnor U11815 (N_11815,N_9661,N_9954);
or U11816 (N_11816,N_9029,N_10394);
xor U11817 (N_11817,N_9464,N_10312);
or U11818 (N_11818,N_10041,N_9369);
nor U11819 (N_11819,N_10178,N_9824);
or U11820 (N_11820,N_9711,N_10180);
and U11821 (N_11821,N_10217,N_9111);
nand U11822 (N_11822,N_9000,N_9182);
nand U11823 (N_11823,N_10048,N_9643);
nand U11824 (N_11824,N_9849,N_9315);
xor U11825 (N_11825,N_9739,N_9158);
xnor U11826 (N_11826,N_9144,N_9597);
xor U11827 (N_11827,N_9391,N_9409);
or U11828 (N_11828,N_9450,N_9132);
nor U11829 (N_11829,N_9115,N_10318);
and U11830 (N_11830,N_10236,N_9092);
xnor U11831 (N_11831,N_9131,N_9253);
nand U11832 (N_11832,N_9014,N_9732);
or U11833 (N_11833,N_9542,N_10395);
xor U11834 (N_11834,N_9404,N_9145);
nand U11835 (N_11835,N_10432,N_9353);
or U11836 (N_11836,N_9187,N_9614);
or U11837 (N_11837,N_9894,N_9579);
or U11838 (N_11838,N_9941,N_9009);
nand U11839 (N_11839,N_9651,N_9813);
xnor U11840 (N_11840,N_9160,N_9118);
or U11841 (N_11841,N_9124,N_9702);
xor U11842 (N_11842,N_9678,N_10265);
and U11843 (N_11843,N_10448,N_9327);
or U11844 (N_11844,N_9451,N_9141);
or U11845 (N_11845,N_9666,N_10308);
and U11846 (N_11846,N_9111,N_9453);
and U11847 (N_11847,N_9432,N_10050);
or U11848 (N_11848,N_9386,N_9816);
xnor U11849 (N_11849,N_10116,N_9961);
nand U11850 (N_11850,N_10212,N_9838);
nor U11851 (N_11851,N_9653,N_9383);
nor U11852 (N_11852,N_9222,N_9150);
xnor U11853 (N_11853,N_9541,N_9513);
xnor U11854 (N_11854,N_9186,N_10187);
or U11855 (N_11855,N_10312,N_9346);
nor U11856 (N_11856,N_10168,N_10154);
or U11857 (N_11857,N_9766,N_10243);
xor U11858 (N_11858,N_9657,N_9619);
nand U11859 (N_11859,N_9931,N_9061);
and U11860 (N_11860,N_10476,N_9989);
and U11861 (N_11861,N_9783,N_10020);
nor U11862 (N_11862,N_10263,N_9741);
nand U11863 (N_11863,N_10049,N_9528);
nor U11864 (N_11864,N_9405,N_9033);
nor U11865 (N_11865,N_10418,N_9770);
nand U11866 (N_11866,N_10496,N_9199);
xor U11867 (N_11867,N_9329,N_9013);
nor U11868 (N_11868,N_9663,N_9847);
nor U11869 (N_11869,N_9049,N_10051);
and U11870 (N_11870,N_9166,N_9172);
xnor U11871 (N_11871,N_9913,N_10081);
nor U11872 (N_11872,N_9432,N_9569);
or U11873 (N_11873,N_9323,N_9485);
or U11874 (N_11874,N_9236,N_9101);
nor U11875 (N_11875,N_9394,N_10435);
and U11876 (N_11876,N_9587,N_9878);
nor U11877 (N_11877,N_9446,N_10427);
and U11878 (N_11878,N_10302,N_10047);
and U11879 (N_11879,N_9430,N_9901);
nand U11880 (N_11880,N_9084,N_9289);
xnor U11881 (N_11881,N_9950,N_10222);
or U11882 (N_11882,N_9142,N_9495);
nor U11883 (N_11883,N_10181,N_9026);
or U11884 (N_11884,N_9582,N_9328);
xor U11885 (N_11885,N_9739,N_10078);
or U11886 (N_11886,N_9826,N_10231);
xnor U11887 (N_11887,N_9099,N_9612);
nand U11888 (N_11888,N_9649,N_9565);
nand U11889 (N_11889,N_10042,N_10236);
and U11890 (N_11890,N_9184,N_10291);
xnor U11891 (N_11891,N_9586,N_10449);
nand U11892 (N_11892,N_10354,N_10269);
nor U11893 (N_11893,N_9288,N_9325);
and U11894 (N_11894,N_10124,N_9406);
or U11895 (N_11895,N_9188,N_9985);
and U11896 (N_11896,N_9182,N_9469);
nor U11897 (N_11897,N_9705,N_9453);
nor U11898 (N_11898,N_9401,N_9939);
nand U11899 (N_11899,N_10202,N_9365);
nand U11900 (N_11900,N_10006,N_10040);
nand U11901 (N_11901,N_9271,N_9648);
nor U11902 (N_11902,N_10078,N_9196);
and U11903 (N_11903,N_9650,N_9200);
and U11904 (N_11904,N_9671,N_9739);
xnor U11905 (N_11905,N_10298,N_10416);
and U11906 (N_11906,N_9744,N_9556);
nand U11907 (N_11907,N_9228,N_9482);
nor U11908 (N_11908,N_9978,N_10462);
nor U11909 (N_11909,N_9433,N_10179);
xnor U11910 (N_11910,N_10360,N_9954);
nor U11911 (N_11911,N_9901,N_10446);
or U11912 (N_11912,N_9333,N_9016);
and U11913 (N_11913,N_9226,N_10490);
nand U11914 (N_11914,N_9325,N_9752);
and U11915 (N_11915,N_9604,N_10169);
xor U11916 (N_11916,N_9286,N_9670);
and U11917 (N_11917,N_9834,N_10106);
xor U11918 (N_11918,N_9037,N_9962);
nor U11919 (N_11919,N_9115,N_9761);
nand U11920 (N_11920,N_10409,N_10185);
nor U11921 (N_11921,N_9808,N_10356);
xor U11922 (N_11922,N_9399,N_9239);
xor U11923 (N_11923,N_10177,N_10406);
nand U11924 (N_11924,N_9251,N_9887);
nor U11925 (N_11925,N_9146,N_9863);
nor U11926 (N_11926,N_10315,N_9154);
nand U11927 (N_11927,N_9844,N_9286);
nor U11928 (N_11928,N_9448,N_9593);
and U11929 (N_11929,N_9959,N_10071);
and U11930 (N_11930,N_9831,N_10403);
nand U11931 (N_11931,N_9494,N_10199);
nand U11932 (N_11932,N_10336,N_9472);
xor U11933 (N_11933,N_10477,N_10104);
nand U11934 (N_11934,N_9475,N_9799);
xor U11935 (N_11935,N_9072,N_9715);
nand U11936 (N_11936,N_9439,N_10029);
nand U11937 (N_11937,N_9845,N_9669);
nand U11938 (N_11938,N_9110,N_10284);
nor U11939 (N_11939,N_9515,N_9582);
nand U11940 (N_11940,N_9498,N_9403);
nor U11941 (N_11941,N_10340,N_10374);
nand U11942 (N_11942,N_9680,N_9270);
nand U11943 (N_11943,N_9704,N_9510);
nor U11944 (N_11944,N_9341,N_9593);
nor U11945 (N_11945,N_10343,N_9533);
nand U11946 (N_11946,N_10067,N_10294);
and U11947 (N_11947,N_10018,N_9305);
and U11948 (N_11948,N_9334,N_9009);
xor U11949 (N_11949,N_9190,N_10385);
xnor U11950 (N_11950,N_9810,N_10399);
nor U11951 (N_11951,N_9769,N_9907);
nand U11952 (N_11952,N_9879,N_9845);
and U11953 (N_11953,N_9503,N_9557);
and U11954 (N_11954,N_9144,N_10377);
or U11955 (N_11955,N_9070,N_9678);
xor U11956 (N_11956,N_9792,N_9351);
xor U11957 (N_11957,N_9765,N_10132);
and U11958 (N_11958,N_10389,N_9142);
nand U11959 (N_11959,N_9769,N_9645);
xor U11960 (N_11960,N_10422,N_10055);
nand U11961 (N_11961,N_9135,N_10165);
and U11962 (N_11962,N_10178,N_10482);
nand U11963 (N_11963,N_9074,N_10111);
and U11964 (N_11964,N_9622,N_9110);
or U11965 (N_11965,N_9945,N_9751);
xnor U11966 (N_11966,N_9858,N_9013);
or U11967 (N_11967,N_9121,N_10079);
and U11968 (N_11968,N_10267,N_9504);
and U11969 (N_11969,N_10417,N_9481);
xnor U11970 (N_11970,N_9060,N_10450);
xnor U11971 (N_11971,N_10352,N_9828);
and U11972 (N_11972,N_9233,N_9833);
xnor U11973 (N_11973,N_9555,N_10116);
or U11974 (N_11974,N_9822,N_10304);
or U11975 (N_11975,N_10011,N_9560);
nand U11976 (N_11976,N_9422,N_10214);
nand U11977 (N_11977,N_9812,N_9217);
or U11978 (N_11978,N_9633,N_10054);
nand U11979 (N_11979,N_9428,N_10168);
xnor U11980 (N_11980,N_9049,N_9607);
or U11981 (N_11981,N_9750,N_10378);
and U11982 (N_11982,N_9176,N_10117);
xnor U11983 (N_11983,N_9582,N_10323);
or U11984 (N_11984,N_9356,N_10239);
and U11985 (N_11985,N_9119,N_9495);
or U11986 (N_11986,N_10373,N_10446);
and U11987 (N_11987,N_9956,N_10060);
or U11988 (N_11988,N_9755,N_9504);
and U11989 (N_11989,N_9652,N_9946);
xnor U11990 (N_11990,N_9604,N_9059);
nand U11991 (N_11991,N_9824,N_10209);
nand U11992 (N_11992,N_10442,N_10063);
nor U11993 (N_11993,N_10139,N_10260);
or U11994 (N_11994,N_9459,N_10458);
xor U11995 (N_11995,N_10131,N_10171);
and U11996 (N_11996,N_9120,N_9329);
xor U11997 (N_11997,N_10126,N_10180);
nand U11998 (N_11998,N_10231,N_10216);
nor U11999 (N_11999,N_10319,N_9721);
xnor U12000 (N_12000,N_10711,N_10944);
nor U12001 (N_12001,N_10745,N_11310);
or U12002 (N_12002,N_11870,N_11545);
nor U12003 (N_12003,N_11512,N_11719);
nor U12004 (N_12004,N_11750,N_11786);
nand U12005 (N_12005,N_11099,N_11768);
or U12006 (N_12006,N_11200,N_11450);
or U12007 (N_12007,N_11509,N_10630);
xnor U12008 (N_12008,N_10727,N_11673);
or U12009 (N_12009,N_11015,N_10951);
nand U12010 (N_12010,N_11458,N_11248);
nand U12011 (N_12011,N_11635,N_11687);
xnor U12012 (N_12012,N_11594,N_11033);
xor U12013 (N_12013,N_10642,N_10996);
or U12014 (N_12014,N_11517,N_11929);
nor U12015 (N_12015,N_10509,N_10969);
xor U12016 (N_12016,N_11727,N_11653);
xnor U12017 (N_12017,N_11550,N_10999);
nor U12018 (N_12018,N_11948,N_11215);
nand U12019 (N_12019,N_11159,N_10656);
and U12020 (N_12020,N_11365,N_11868);
xnor U12021 (N_12021,N_11129,N_11337);
nor U12022 (N_12022,N_11655,N_11206);
nand U12023 (N_12023,N_11490,N_11505);
or U12024 (N_12024,N_11158,N_11493);
nand U12025 (N_12025,N_10571,N_10804);
and U12026 (N_12026,N_11724,N_11104);
or U12027 (N_12027,N_11026,N_11187);
nand U12028 (N_12028,N_11809,N_11559);
xnor U12029 (N_12029,N_11895,N_10643);
or U12030 (N_12030,N_10654,N_10907);
nor U12031 (N_12031,N_10742,N_11257);
nor U12032 (N_12032,N_11642,N_10629);
nand U12033 (N_12033,N_11621,N_11848);
nand U12034 (N_12034,N_11637,N_10635);
xor U12035 (N_12035,N_11538,N_11306);
nor U12036 (N_12036,N_11580,N_11228);
nand U12037 (N_12037,N_11772,N_11836);
and U12038 (N_12038,N_11562,N_11424);
nand U12039 (N_12039,N_11074,N_11363);
nor U12040 (N_12040,N_10661,N_10522);
nand U12041 (N_12041,N_11987,N_11284);
or U12042 (N_12042,N_11759,N_11318);
xnor U12043 (N_12043,N_11633,N_10750);
nor U12044 (N_12044,N_11057,N_11077);
nor U12045 (N_12045,N_11526,N_11276);
nand U12046 (N_12046,N_10720,N_11646);
and U12047 (N_12047,N_10834,N_11247);
nand U12048 (N_12048,N_11991,N_11064);
and U12049 (N_12049,N_11027,N_10556);
and U12050 (N_12050,N_11155,N_11445);
or U12051 (N_12051,N_11919,N_11875);
xnor U12052 (N_12052,N_11934,N_10774);
or U12053 (N_12053,N_11502,N_11908);
and U12054 (N_12054,N_11715,N_11983);
and U12055 (N_12055,N_10660,N_10922);
xor U12056 (N_12056,N_11397,N_11881);
nand U12057 (N_12057,N_11349,N_10825);
xor U12058 (N_12058,N_11704,N_11495);
nor U12059 (N_12059,N_11938,N_11196);
or U12060 (N_12060,N_11024,N_10505);
or U12061 (N_12061,N_11234,N_11554);
and U12062 (N_12062,N_10705,N_10702);
xnor U12063 (N_12063,N_10559,N_11326);
or U12064 (N_12064,N_11792,N_10506);
nand U12065 (N_12065,N_11080,N_11877);
or U12066 (N_12066,N_10903,N_10770);
and U12067 (N_12067,N_11328,N_11553);
nand U12068 (N_12068,N_11639,N_11497);
and U12069 (N_12069,N_10688,N_11858);
xor U12070 (N_12070,N_10896,N_11720);
or U12071 (N_12071,N_11455,N_11590);
nand U12072 (N_12072,N_11360,N_11779);
nor U12073 (N_12073,N_10726,N_11543);
xor U12074 (N_12074,N_11971,N_11616);
xnor U12075 (N_12075,N_11128,N_11043);
nand U12076 (N_12076,N_11804,N_10572);
nor U12077 (N_12077,N_10843,N_10703);
and U12078 (N_12078,N_11636,N_11912);
nor U12079 (N_12079,N_11066,N_11652);
nand U12080 (N_12080,N_11463,N_11243);
nor U12081 (N_12081,N_10611,N_11816);
and U12082 (N_12082,N_10956,N_11709);
nand U12083 (N_12083,N_11974,N_10963);
and U12084 (N_12084,N_10827,N_11609);
xor U12085 (N_12085,N_11765,N_11420);
or U12086 (N_12086,N_11489,N_11299);
xor U12087 (N_12087,N_11356,N_11939);
xnor U12088 (N_12088,N_10916,N_11574);
or U12089 (N_12089,N_11465,N_11408);
nand U12090 (N_12090,N_11712,N_11675);
nand U12091 (N_12091,N_10771,N_10679);
and U12092 (N_12092,N_11643,N_10796);
nor U12093 (N_12093,N_11028,N_10980);
nor U12094 (N_12094,N_10680,N_11118);
nand U12095 (N_12095,N_11253,N_11492);
and U12096 (N_12096,N_11857,N_11901);
and U12097 (N_12097,N_11905,N_10676);
or U12098 (N_12098,N_10718,N_11321);
and U12099 (N_12099,N_11604,N_11979);
and U12100 (N_12100,N_11418,N_11127);
nand U12101 (N_12101,N_10936,N_11893);
nand U12102 (N_12102,N_11319,N_10909);
xor U12103 (N_12103,N_11100,N_11823);
or U12104 (N_12104,N_11138,N_11866);
and U12105 (N_12105,N_11072,N_11903);
nor U12106 (N_12106,N_11936,N_11101);
nand U12107 (N_12107,N_10613,N_11812);
nor U12108 (N_12108,N_11476,N_10520);
and U12109 (N_12109,N_10507,N_10952);
xnor U12110 (N_12110,N_11746,N_11725);
and U12111 (N_12111,N_11392,N_10684);
nor U12112 (N_12112,N_11157,N_10723);
or U12113 (N_12113,N_10518,N_10886);
xnor U12114 (N_12114,N_11953,N_10816);
nand U12115 (N_12115,N_11928,N_10538);
and U12116 (N_12116,N_11203,N_11946);
xor U12117 (N_12117,N_11689,N_11568);
xor U12118 (N_12118,N_11073,N_11593);
or U12119 (N_12119,N_11051,N_11210);
nor U12120 (N_12120,N_11666,N_11479);
nor U12121 (N_12121,N_11718,N_11930);
and U12122 (N_12122,N_11638,N_11193);
xnor U12123 (N_12123,N_11199,N_11841);
xnor U12124 (N_12124,N_11025,N_11041);
and U12125 (N_12125,N_10540,N_11143);
xor U12126 (N_12126,N_11068,N_10740);
nand U12127 (N_12127,N_11592,N_11737);
and U12128 (N_12128,N_11270,N_10695);
nand U12129 (N_12129,N_10650,N_11327);
and U12130 (N_12130,N_11464,N_11373);
xor U12131 (N_12131,N_11021,N_11045);
nor U12132 (N_12132,N_10889,N_11470);
xor U12133 (N_12133,N_11958,N_10512);
nand U12134 (N_12134,N_10555,N_11396);
nand U12135 (N_12135,N_10706,N_11165);
nand U12136 (N_12136,N_10819,N_10839);
nand U12137 (N_12137,N_11314,N_10970);
xnor U12138 (N_12138,N_10582,N_11387);
nand U12139 (N_12139,N_11589,N_11743);
and U12140 (N_12140,N_10817,N_10754);
or U12141 (N_12141,N_10966,N_10531);
nand U12142 (N_12142,N_11347,N_10870);
nor U12143 (N_12143,N_10850,N_11218);
xor U12144 (N_12144,N_11226,N_11240);
nand U12145 (N_12145,N_11130,N_11126);
and U12146 (N_12146,N_10788,N_11726);
nor U12147 (N_12147,N_10655,N_11307);
and U12148 (N_12148,N_11947,N_10781);
nand U12149 (N_12149,N_11566,N_10514);
nand U12150 (N_12150,N_11849,N_10618);
nand U12151 (N_12151,N_11195,N_11255);
and U12152 (N_12152,N_11410,N_11703);
nand U12153 (N_12153,N_11518,N_10561);
nand U12154 (N_12154,N_11522,N_11379);
xor U12155 (N_12155,N_11585,N_11829);
nor U12156 (N_12156,N_11790,N_10810);
nand U12157 (N_12157,N_11457,N_10529);
or U12158 (N_12158,N_11006,N_10837);
nor U12159 (N_12159,N_10586,N_11851);
and U12160 (N_12160,N_11884,N_11002);
or U12161 (N_12161,N_10647,N_10793);
xnor U12162 (N_12162,N_11969,N_11472);
xor U12163 (N_12163,N_10717,N_11362);
and U12164 (N_12164,N_11565,N_11915);
and U12165 (N_12165,N_11649,N_11173);
and U12166 (N_12166,N_11007,N_11521);
or U12167 (N_12167,N_11582,N_11401);
and U12168 (N_12168,N_11607,N_10607);
nor U12169 (N_12169,N_11448,N_10517);
xor U12170 (N_12170,N_11169,N_10857);
or U12171 (N_12171,N_11442,N_11180);
and U12172 (N_12172,N_11966,N_11177);
or U12173 (N_12173,N_11113,N_11413);
nand U12174 (N_12174,N_10867,N_10585);
and U12175 (N_12175,N_10734,N_10544);
xor U12176 (N_12176,N_11437,N_11668);
nor U12177 (N_12177,N_11811,N_11439);
nor U12178 (N_12178,N_10880,N_11899);
xnor U12179 (N_12179,N_10962,N_11451);
nor U12180 (N_12180,N_11188,N_11935);
and U12181 (N_12181,N_11814,N_10534);
xor U12182 (N_12182,N_11046,N_10609);
or U12183 (N_12183,N_10764,N_11667);
or U12184 (N_12184,N_11535,N_11569);
or U12185 (N_12185,N_11528,N_11432);
nor U12186 (N_12186,N_10532,N_10605);
xor U12187 (N_12187,N_10649,N_11350);
nand U12188 (N_12188,N_10574,N_11163);
or U12189 (N_12189,N_10998,N_10710);
xor U12190 (N_12190,N_11778,N_11441);
and U12191 (N_12191,N_11296,N_10504);
and U12192 (N_12192,N_11632,N_11133);
nor U12193 (N_12193,N_10692,N_10523);
and U12194 (N_12194,N_11047,N_10694);
nor U12195 (N_12195,N_11523,N_10537);
and U12196 (N_12196,N_11008,N_10614);
or U12197 (N_12197,N_10873,N_10871);
and U12198 (N_12198,N_10791,N_11467);
and U12199 (N_12199,N_11287,N_10566);
or U12200 (N_12200,N_10636,N_10878);
nand U12201 (N_12201,N_11970,N_11229);
nor U12202 (N_12202,N_11277,N_11009);
and U12203 (N_12203,N_11692,N_11909);
or U12204 (N_12204,N_10578,N_11600);
or U12205 (N_12205,N_11605,N_10964);
nor U12206 (N_12206,N_11601,N_11300);
xnor U12207 (N_12207,N_10883,N_10704);
or U12208 (N_12208,N_11878,N_11656);
nand U12209 (N_12209,N_11411,N_11407);
xnor U12210 (N_12210,N_11861,N_10939);
nor U12211 (N_12211,N_10855,N_11531);
or U12212 (N_12212,N_10906,N_11251);
and U12213 (N_12213,N_11902,N_11052);
nand U12214 (N_12214,N_10776,N_11941);
nor U12215 (N_12215,N_11452,N_11537);
xnor U12216 (N_12216,N_11579,N_10800);
and U12217 (N_12217,N_11124,N_11670);
nor U12218 (N_12218,N_11886,N_10846);
nor U12219 (N_12219,N_11406,N_11209);
xnor U12220 (N_12220,N_11520,N_10553);
or U12221 (N_12221,N_11087,N_11748);
and U12222 (N_12222,N_11576,N_11863);
xor U12223 (N_12223,N_10844,N_10608);
nor U12224 (N_12224,N_10925,N_10890);
nor U12225 (N_12225,N_10866,N_10603);
or U12226 (N_12226,N_11791,N_11181);
xnor U12227 (N_12227,N_10851,N_10623);
or U12228 (N_12228,N_11611,N_11053);
nor U12229 (N_12229,N_11612,N_11063);
nor U12230 (N_12230,N_11696,N_11835);
or U12231 (N_12231,N_11731,N_10881);
nand U12232 (N_12232,N_11211,N_10780);
xnor U12233 (N_12233,N_11894,N_11144);
or U12234 (N_12234,N_11162,N_11586);
or U12235 (N_12235,N_11910,N_11681);
and U12236 (N_12236,N_11984,N_11595);
nand U12237 (N_12237,N_10511,N_11446);
or U12238 (N_12238,N_10539,N_10550);
xnor U12239 (N_12239,N_11044,N_11572);
nor U12240 (N_12240,N_10986,N_11182);
xor U12241 (N_12241,N_11274,N_11444);
nor U12242 (N_12242,N_11993,N_11891);
xor U12243 (N_12243,N_11892,N_11977);
and U12244 (N_12244,N_11515,N_11659);
nand U12245 (N_12245,N_11065,N_11781);
xor U12246 (N_12246,N_10591,N_11887);
nor U12247 (N_12247,N_11660,N_11419);
nand U12248 (N_12248,N_11753,N_10905);
or U12249 (N_12249,N_11599,N_11664);
nand U12250 (N_12250,N_11943,N_10516);
nor U12251 (N_12251,N_11510,N_10786);
xnor U12252 (N_12252,N_11810,N_11959);
nand U12253 (N_12253,N_10610,N_11242);
nor U12254 (N_12254,N_10564,N_11558);
and U12255 (N_12255,N_10849,N_11888);
and U12256 (N_12256,N_11376,N_10845);
or U12257 (N_12257,N_11076,N_11844);
nor U12258 (N_12258,N_11271,N_11440);
xor U12259 (N_12259,N_11091,N_11346);
or U12260 (N_12260,N_10882,N_10784);
xor U12261 (N_12261,N_11377,N_11294);
and U12262 (N_12262,N_11949,N_11466);
or U12263 (N_12263,N_11691,N_10648);
xnor U12264 (N_12264,N_11353,N_10926);
nor U12265 (N_12265,N_11685,N_11175);
nor U12266 (N_12266,N_11096,N_10666);
and U12267 (N_12267,N_10693,N_11343);
nor U12268 (N_12268,N_11429,N_10665);
nor U12269 (N_12269,N_10722,N_11216);
xnor U12270 (N_12270,N_10747,N_11000);
xor U12271 (N_12271,N_11031,N_11864);
xnor U12272 (N_12272,N_11333,N_11796);
or U12273 (N_12273,N_10616,N_11312);
and U12274 (N_12274,N_11749,N_11005);
xnor U12275 (N_12275,N_11264,N_10859);
or U12276 (N_12276,N_10949,N_10502);
nand U12277 (N_12277,N_10932,N_10976);
and U12278 (N_12278,N_11771,N_11239);
and U12279 (N_12279,N_11230,N_11086);
xnor U12280 (N_12280,N_10592,N_10779);
xnor U12281 (N_12281,N_10904,N_11067);
or U12282 (N_12282,N_11571,N_11539);
or U12283 (N_12283,N_10674,N_10872);
nand U12284 (N_12284,N_11303,N_10961);
xor U12285 (N_12285,N_10785,N_11821);
and U12286 (N_12286,N_11733,N_11161);
or U12287 (N_12287,N_11603,N_10596);
nand U12288 (N_12288,N_11121,N_11975);
nor U12289 (N_12289,N_10624,N_11116);
xnor U12290 (N_12290,N_10792,N_11190);
or U12291 (N_12291,N_11221,N_11862);
or U12292 (N_12292,N_10831,N_11534);
nor U12293 (N_12293,N_10766,N_10746);
nand U12294 (N_12294,N_11281,N_10991);
nor U12295 (N_12295,N_11679,N_10924);
and U12296 (N_12296,N_11735,N_11202);
and U12297 (N_12297,N_11815,N_11354);
nand U12298 (N_12298,N_11485,N_10668);
or U12299 (N_12299,N_10639,N_11705);
and U12300 (N_12300,N_11702,N_10876);
nand U12301 (N_12301,N_11361,N_11828);
xnor U12302 (N_12302,N_10777,N_11114);
nand U12303 (N_12303,N_11334,N_11784);
xnor U12304 (N_12304,N_11856,N_11707);
and U12305 (N_12305,N_10653,N_10590);
xor U12306 (N_12306,N_11629,N_11978);
nand U12307 (N_12307,N_10937,N_11508);
and U12308 (N_12308,N_10802,N_11069);
xnor U12309 (N_12309,N_11070,N_10958);
nor U12310 (N_12310,N_10978,N_11140);
nor U12311 (N_12311,N_11739,N_10945);
nand U12312 (N_12312,N_11246,N_10858);
and U12313 (N_12313,N_11491,N_10874);
nand U12314 (N_12314,N_11054,N_11785);
or U12315 (N_12315,N_11488,N_11674);
and U12316 (N_12316,N_10911,N_10893);
nand U12317 (N_12317,N_11817,N_11220);
nor U12318 (N_12318,N_11701,N_10569);
or U12319 (N_12319,N_10736,N_10875);
and U12320 (N_12320,N_11222,N_10664);
or U12321 (N_12321,N_11142,N_10887);
xnor U12322 (N_12322,N_11298,N_11961);
nand U12323 (N_12323,N_10767,N_11560);
xnor U12324 (N_12324,N_10775,N_10806);
and U12325 (N_12325,N_11166,N_10987);
and U12326 (N_12326,N_11677,N_11214);
nor U12327 (N_12327,N_11436,N_10808);
or U12328 (N_12328,N_10910,N_10852);
and U12329 (N_12329,N_11430,N_11381);
nor U12330 (N_12330,N_10955,N_10812);
nand U12331 (N_12331,N_11117,N_11747);
or U12332 (N_12332,N_11108,N_10601);
or U12333 (N_12333,N_10801,N_11095);
nor U12334 (N_12334,N_10933,N_11793);
xor U12335 (N_12335,N_11774,N_10739);
or U12336 (N_12336,N_11478,N_10860);
nand U12337 (N_12337,N_11414,N_11336);
or U12338 (N_12338,N_10515,N_11665);
nor U12339 (N_12339,N_11014,N_11624);
and U12340 (N_12340,N_11194,N_11316);
xnor U12341 (N_12341,N_11711,N_11083);
or U12342 (N_12342,N_11507,N_10580);
nand U12343 (N_12343,N_10683,N_10892);
nor U12344 (N_12344,N_11797,N_10640);
nor U12345 (N_12345,N_11807,N_11514);
or U12346 (N_12346,N_10715,N_11421);
xor U12347 (N_12347,N_10545,N_11504);
nor U12348 (N_12348,N_11198,N_10573);
and U12349 (N_12349,N_11004,N_11358);
and U12350 (N_12350,N_10584,N_11345);
nand U12351 (N_12351,N_11871,N_11662);
nand U12352 (N_12352,N_11153,N_11952);
or U12353 (N_12353,N_11205,N_11237);
xor U12354 (N_12354,N_11106,N_11141);
and U12355 (N_12355,N_11967,N_10923);
and U12356 (N_12356,N_11090,N_10954);
xor U12357 (N_12357,N_11266,N_11956);
nor U12358 (N_12358,N_11272,N_11911);
nor U12359 (N_12359,N_10563,N_11304);
nand U12360 (N_12360,N_10644,N_11992);
and U12361 (N_12361,N_11957,N_11650);
and U12362 (N_12362,N_11453,N_11780);
and U12363 (N_12363,N_11275,N_11179);
nor U12364 (N_12364,N_11530,N_11093);
or U12365 (N_12365,N_10928,N_11285);
nand U12366 (N_12366,N_11907,N_10697);
nor U12367 (N_12367,N_10678,N_11315);
nor U12368 (N_12368,N_11317,N_11940);
xnor U12369 (N_12369,N_10841,N_10913);
and U12370 (N_12370,N_11532,N_10967);
or U12371 (N_12371,N_11965,N_10513);
nand U12372 (N_12372,N_11762,N_10814);
and U12373 (N_12373,N_10576,N_11519);
and U12374 (N_12374,N_10988,N_10990);
nor U12375 (N_12375,N_11787,N_11925);
xnor U12376 (N_12376,N_10594,N_10617);
nand U12377 (N_12377,N_10918,N_10593);
xor U12378 (N_12378,N_11798,N_11852);
nand U12379 (N_12379,N_11741,N_11680);
xor U12380 (N_12380,N_11035,N_11029);
and U12381 (N_12381,N_10914,N_11769);
and U12382 (N_12382,N_11156,N_11032);
or U12383 (N_12383,N_11955,N_10753);
and U12384 (N_12384,N_10769,N_11999);
xor U12385 (N_12385,N_11588,N_11754);
or U12386 (N_12386,N_10546,N_11475);
and U12387 (N_12387,N_11827,N_11308);
xnor U12388 (N_12388,N_11001,N_11695);
nand U12389 (N_12389,N_11351,N_10543);
nand U12390 (N_12390,N_11320,N_11980);
or U12391 (N_12391,N_11846,N_11972);
or U12392 (N_12392,N_11596,N_10599);
and U12393 (N_12393,N_10638,N_11217);
or U12394 (N_12394,N_11698,N_10789);
xor U12395 (N_12395,N_10815,N_11613);
or U12396 (N_12396,N_11567,N_10588);
nor U12397 (N_12397,N_11191,N_10912);
and U12398 (N_12398,N_11721,N_11012);
xnor U12399 (N_12399,N_10687,N_10549);
or U12400 (N_12400,N_11832,N_10861);
xnor U12401 (N_12401,N_10847,N_10899);
or U12402 (N_12402,N_11716,N_11071);
xnor U12403 (N_12403,N_10853,N_11942);
nand U12404 (N_12404,N_11438,N_11498);
xnor U12405 (N_12405,N_10790,N_11167);
nor U12406 (N_12406,N_11988,N_11135);
nand U12407 (N_12407,N_11736,N_11602);
or U12408 (N_12408,N_11147,N_11697);
nor U12409 (N_12409,N_11795,N_11295);
xnor U12410 (N_12410,N_11079,N_11500);
nand U12411 (N_12411,N_10983,N_11088);
nor U12412 (N_12412,N_11366,N_11869);
xor U12413 (N_12413,N_10552,N_11710);
xnor U12414 (N_12414,N_10631,N_11766);
nor U12415 (N_12415,N_10778,N_11648);
nand U12416 (N_12416,N_11591,N_11060);
nor U12417 (N_12417,N_10671,N_11149);
and U12418 (N_12418,N_10921,N_11192);
and U12419 (N_12419,N_11575,N_11482);
nand U12420 (N_12420,N_11728,N_11986);
and U12421 (N_12421,N_11564,N_10818);
or U12422 (N_12422,N_11803,N_11996);
nor U12423 (N_12423,N_11922,N_10824);
nand U12424 (N_12424,N_10995,N_11431);
or U12425 (N_12425,N_10669,N_11368);
or U12426 (N_12426,N_11380,N_11962);
xor U12427 (N_12427,N_11486,N_11644);
or U12428 (N_12428,N_11404,N_11018);
nand U12429 (N_12429,N_11085,N_10562);
xor U12430 (N_12430,N_11402,N_11740);
nand U12431 (N_12431,N_10807,N_10673);
nand U12432 (N_12432,N_11831,N_11865);
or U12433 (N_12433,N_11122,N_10690);
or U12434 (N_12434,N_11061,N_11838);
or U12435 (N_12435,N_11174,N_11617);
or U12436 (N_12436,N_11917,N_11839);
xnor U12437 (N_12437,N_11391,N_11082);
nor U12438 (N_12438,N_11089,N_10637);
xnor U12439 (N_12439,N_10752,N_11322);
or U12440 (N_12440,N_11422,N_11120);
nor U12441 (N_12441,N_11729,N_10565);
or U12442 (N_12442,N_11706,N_11717);
or U12443 (N_12443,N_11168,N_10536);
and U12444 (N_12444,N_11081,N_10598);
xnor U12445 (N_12445,N_11761,N_11950);
xor U12446 (N_12446,N_10842,N_11541);
xor U12447 (N_12447,N_11540,N_11324);
nor U12448 (N_12448,N_11584,N_11669);
and U12449 (N_12449,N_11259,N_10943);
nand U12450 (N_12450,N_11049,N_11389);
xor U12451 (N_12451,N_10689,N_11577);
nand U12452 (N_12452,N_10768,N_11906);
xnor U12453 (N_12453,N_11386,N_11760);
xnor U12454 (N_12454,N_11244,N_10732);
xnor U12455 (N_12455,N_11151,N_11011);
and U12456 (N_12456,N_10898,N_11896);
xnor U12457 (N_12457,N_11631,N_10959);
and U12458 (N_12458,N_11723,N_10743);
nor U12459 (N_12459,N_11783,N_11494);
nand U12460 (N_12460,N_11103,N_10838);
or U12461 (N_12461,N_10579,N_11506);
and U12462 (N_12462,N_11503,N_11964);
or U12463 (N_12463,N_11425,N_11527);
or U12464 (N_12464,N_11806,N_10530);
or U12465 (N_12465,N_11820,N_11039);
nand U12466 (N_12466,N_10685,N_11037);
and U12467 (N_12467,N_11139,N_10942);
xnor U12468 (N_12468,N_11914,N_11678);
and U12469 (N_12469,N_11265,N_10548);
nand U12470 (N_12470,N_11843,N_10950);
nand U12471 (N_12471,N_11433,N_10641);
nor U12472 (N_12472,N_10938,N_11890);
and U12473 (N_12473,N_11808,N_11375);
xnor U12474 (N_12474,N_10981,N_11184);
xor U12475 (N_12475,N_10863,N_11824);
or U12476 (N_12476,N_11235,N_11344);
nor U12477 (N_12477,N_11826,N_11767);
nor U12478 (N_12478,N_10568,N_11456);
or U12479 (N_12479,N_11618,N_11227);
xor U12480 (N_12480,N_11098,N_11551);
xor U12481 (N_12481,N_11867,N_11288);
nor U12482 (N_12482,N_10560,N_11136);
or U12483 (N_12483,N_10587,N_11305);
xor U12484 (N_12484,N_11763,N_10542);
and U12485 (N_12485,N_11152,N_11250);
nand U12486 (N_12486,N_11933,N_11186);
and U12487 (N_12487,N_10934,N_11889);
and U12488 (N_12488,N_11020,N_10628);
nand U12489 (N_12489,N_11547,N_10888);
nor U12490 (N_12490,N_10541,N_10953);
or U12491 (N_12491,N_11799,N_10833);
xnor U12492 (N_12492,N_10662,N_11078);
nor U12493 (N_12493,N_11770,N_11383);
and U12494 (N_12494,N_11399,N_11332);
nor U12495 (N_12495,N_10760,N_11758);
or U12496 (N_12496,N_10652,N_11654);
and U12497 (N_12497,N_11625,N_11058);
nor U12498 (N_12498,N_10900,N_11622);
or U12499 (N_12499,N_10691,N_11570);
nor U12500 (N_12500,N_11742,N_11297);
or U12501 (N_12501,N_11985,N_10524);
and U12502 (N_12502,N_10634,N_11170);
and U12503 (N_12503,N_11850,N_11447);
or U12504 (N_12504,N_11403,N_11378);
and U12505 (N_12505,N_11262,N_10994);
or U12506 (N_12506,N_10567,N_11496);
xor U12507 (N_12507,N_11405,N_11134);
xnor U12508 (N_12508,N_11462,N_10948);
or U12509 (N_12509,N_11471,N_11651);
nand U12510 (N_12510,N_11830,N_10535);
and U12511 (N_12511,N_11511,N_11897);
and U12512 (N_12512,N_11212,N_10595);
xor U12513 (N_12513,N_11676,N_11150);
nand U12514 (N_12514,N_10619,N_10947);
nor U12515 (N_12515,N_11097,N_11944);
xnor U12516 (N_12516,N_11207,N_10583);
and U12517 (N_12517,N_11623,N_10772);
nor U12518 (N_12518,N_10716,N_11722);
nand U12519 (N_12519,N_11435,N_11876);
nor U12520 (N_12520,N_11647,N_11423);
nor U12521 (N_12521,N_11688,N_11777);
nor U12522 (N_12522,N_11487,N_11918);
or U12523 (N_12523,N_10960,N_11578);
and U12524 (N_12524,N_10667,N_11880);
nand U12525 (N_12525,N_11714,N_11546);
nor U12526 (N_12526,N_11428,N_11094);
or U12527 (N_12527,N_11374,N_11443);
nor U12528 (N_12528,N_11700,N_10798);
and U12529 (N_12529,N_11672,N_11657);
and U12530 (N_12530,N_11708,N_11394);
nor U12531 (N_12531,N_11178,N_11788);
xnor U12532 (N_12532,N_11256,N_11882);
nand U12533 (N_12533,N_10713,N_10701);
xnor U12534 (N_12534,N_11010,N_11335);
nand U12535 (N_12535,N_10620,N_11279);
nand U12536 (N_12536,N_11110,N_11183);
xor U12537 (N_12537,N_10759,N_10749);
nand U12538 (N_12538,N_11348,N_11663);
xor U12539 (N_12539,N_10737,N_11055);
xnor U12540 (N_12540,N_11197,N_11610);
nor U12541 (N_12541,N_11084,N_11059);
and U12542 (N_12542,N_11125,N_10622);
or U12543 (N_12543,N_11208,N_10989);
xor U12544 (N_12544,N_11822,N_11751);
and U12545 (N_12545,N_11968,N_10526);
nand U12546 (N_12546,N_11819,N_10621);
nor U12547 (N_12547,N_10920,N_11286);
or U12548 (N_12548,N_11292,N_10557);
xnor U12549 (N_12549,N_10698,N_10977);
or U12550 (N_12550,N_11241,N_11615);
and U12551 (N_12551,N_10659,N_10554);
xor U12552 (N_12552,N_10974,N_11415);
nand U12553 (N_12553,N_11395,N_10709);
and U12554 (N_12554,N_11734,N_10729);
or U12555 (N_12555,N_10795,N_11920);
nor U12556 (N_12556,N_11682,N_10809);
nor U12557 (N_12557,N_11801,N_11854);
xnor U12558 (N_12558,N_10927,N_11367);
nor U12559 (N_12559,N_11499,N_10547);
or U12560 (N_12560,N_11645,N_10525);
nand U12561 (N_12561,N_10696,N_11879);
xor U12562 (N_12562,N_11641,N_11238);
nand U12563 (N_12563,N_11185,N_11626);
or U12564 (N_12564,N_11544,N_10820);
xor U12565 (N_12565,N_11369,N_11075);
or U12566 (N_12566,N_11323,N_11923);
nand U12567 (N_12567,N_11782,N_10829);
xnor U12568 (N_12568,N_11834,N_11459);
nand U12569 (N_12569,N_10708,N_11254);
and U12570 (N_12570,N_11548,N_10930);
or U12571 (N_12571,N_10738,N_11873);
and U12572 (N_12572,N_10589,N_10551);
or U12573 (N_12573,N_11837,N_11261);
nand U12574 (N_12574,N_11105,N_10803);
nand U12575 (N_12575,N_10675,N_11524);
xor U12576 (N_12576,N_10500,N_11267);
nand U12577 (N_12577,N_10681,N_10570);
nor U12578 (N_12578,N_11699,N_10811);
nand U12579 (N_12579,N_10645,N_10558);
and U12580 (N_12580,N_11628,N_11164);
and U12581 (N_12581,N_11536,N_11683);
xor U12582 (N_12582,N_11982,N_10794);
xor U12583 (N_12583,N_11400,N_11690);
and U12584 (N_12584,N_11313,N_11555);
nor U12585 (N_12585,N_11338,N_10612);
nand U12586 (N_12586,N_11794,N_11598);
or U12587 (N_12587,N_11301,N_10626);
xnor U12588 (N_12588,N_11092,N_11755);
or U12589 (N_12589,N_10658,N_11732);
nor U12590 (N_12590,N_10832,N_10724);
and U12591 (N_12591,N_10744,N_10915);
or U12592 (N_12592,N_11818,N_11671);
or U12593 (N_12593,N_11030,N_10633);
nand U12594 (N_12594,N_11213,N_11370);
or U12595 (N_12595,N_11461,N_11813);
nand U12596 (N_12596,N_11390,N_11263);
nand U12597 (N_12597,N_11752,N_10897);
nor U12598 (N_12598,N_10510,N_10891);
nor U12599 (N_12599,N_11840,N_11963);
xor U12600 (N_12600,N_11409,N_11232);
nand U12601 (N_12601,N_11385,N_11454);
xor U12602 (N_12602,N_10757,N_10884);
nor U12603 (N_12603,N_10751,N_11309);
nor U12604 (N_12604,N_11290,N_10755);
or U12605 (N_12605,N_11204,N_11278);
nand U12606 (N_12606,N_10805,N_11417);
or U12607 (N_12607,N_11756,N_11017);
xnor U12608 (N_12608,N_11269,N_11842);
xnor U12609 (N_12609,N_11289,N_10758);
nor U12610 (N_12610,N_11393,N_10606);
and U12611 (N_12611,N_11927,N_11268);
or U12612 (N_12612,N_11034,N_10917);
nand U12613 (N_12613,N_11847,N_11776);
nor U12614 (N_12614,N_11932,N_11913);
xor U12615 (N_12615,N_11019,N_11427);
xor U12616 (N_12616,N_11516,N_10782);
nand U12617 (N_12617,N_11148,N_10646);
xnor U12618 (N_12618,N_11426,N_10957);
or U12619 (N_12619,N_10877,N_11658);
nand U12620 (N_12620,N_11661,N_11249);
xnor U12621 (N_12621,N_11119,N_11355);
or U12622 (N_12622,N_11614,N_11608);
nor U12623 (N_12623,N_10651,N_10677);
and U12624 (N_12624,N_11483,N_10748);
nand U12625 (N_12625,N_11145,N_10735);
and U12626 (N_12626,N_11112,N_11477);
and U12627 (N_12627,N_11481,N_11951);
xor U12628 (N_12628,N_10992,N_11291);
nor U12629 (N_12629,N_10712,N_11111);
xor U12630 (N_12630,N_11542,N_11146);
nor U12631 (N_12631,N_11738,N_11630);
nor U12632 (N_12632,N_11040,N_11468);
or U12633 (N_12633,N_10577,N_11885);
nor U12634 (N_12634,N_10521,N_10733);
nand U12635 (N_12635,N_10971,N_11359);
nand U12636 (N_12636,N_11331,N_10797);
and U12637 (N_12637,N_11042,N_11398);
or U12638 (N_12638,N_10828,N_11022);
or U12639 (N_12639,N_11382,N_11619);
xnor U12640 (N_12640,N_11587,N_11860);
nand U12641 (N_12641,N_10719,N_10503);
and U12642 (N_12642,N_11744,N_11800);
and U12643 (N_12643,N_10508,N_10929);
or U12644 (N_12644,N_11990,N_11900);
nand U12645 (N_12645,N_11038,N_11371);
xor U12646 (N_12646,N_11412,N_11132);
and U12647 (N_12647,N_11960,N_11325);
nand U12648 (N_12648,N_11469,N_10979);
nand U12649 (N_12649,N_10763,N_10919);
or U12650 (N_12650,N_11805,N_11773);
xnor U12651 (N_12651,N_10625,N_11449);
nor U12652 (N_12652,N_11339,N_11694);
nor U12653 (N_12653,N_11583,N_10728);
nor U12654 (N_12654,N_11557,N_10993);
or U12655 (N_12655,N_10941,N_11258);
nand U12656 (N_12656,N_11916,N_10670);
and U12657 (N_12657,N_11921,N_10725);
and U12658 (N_12658,N_10965,N_10799);
or U12659 (N_12659,N_10840,N_10721);
nor U12660 (N_12660,N_11016,N_11050);
nor U12661 (N_12661,N_11102,N_10908);
and U12662 (N_12662,N_11201,N_10869);
and U12663 (N_12663,N_11561,N_11107);
and U12664 (N_12664,N_11231,N_11364);
xnor U12665 (N_12665,N_11981,N_10821);
and U12666 (N_12666,N_11245,N_11552);
xor U12667 (N_12667,N_11013,N_11219);
nor U12668 (N_12668,N_11789,N_11233);
and U12669 (N_12669,N_10602,N_11926);
xor U12670 (N_12670,N_11460,N_11802);
xor U12671 (N_12671,N_10868,N_10823);
nand U12672 (N_12672,N_11989,N_11845);
nand U12673 (N_12673,N_10885,N_11954);
nor U12674 (N_12674,N_11513,N_11236);
xor U12675 (N_12675,N_11859,N_11924);
and U12676 (N_12676,N_11825,N_11048);
nand U12677 (N_12677,N_11904,N_11023);
nor U12678 (N_12678,N_10663,N_11995);
xor U12679 (N_12679,N_10783,N_10901);
nand U12680 (N_12680,N_10707,N_10686);
xor U12681 (N_12681,N_10672,N_11160);
nand U12682 (N_12682,N_11329,N_11556);
nor U12683 (N_12683,N_11529,N_11123);
xnor U12684 (N_12684,N_11533,N_11003);
nor U12685 (N_12685,N_11998,N_10982);
nand U12686 (N_12686,N_10627,N_11997);
or U12687 (N_12687,N_11388,N_11757);
or U12688 (N_12688,N_11764,N_11293);
nand U12689 (N_12689,N_11855,N_10730);
or U12690 (N_12690,N_11898,N_10835);
nand U12691 (N_12691,N_10940,N_11937);
nand U12692 (N_12692,N_10997,N_11352);
or U12693 (N_12693,N_11131,N_11994);
or U12694 (N_12694,N_10972,N_10682);
and U12695 (N_12695,N_10854,N_10575);
nand U12696 (N_12696,N_11686,N_11172);
xnor U12697 (N_12697,N_11283,N_11973);
or U12698 (N_12698,N_11260,N_11874);
or U12699 (N_12699,N_11730,N_11976);
and U12700 (N_12700,N_11302,N_11473);
xor U12701 (N_12701,N_11171,N_10528);
and U12702 (N_12702,N_11480,N_11273);
nand U12703 (N_12703,N_10973,N_11225);
nand U12704 (N_12704,N_11357,N_10714);
and U12705 (N_12705,N_10787,N_11062);
or U12706 (N_12706,N_10581,N_11474);
nand U12707 (N_12707,N_11693,N_10761);
xor U12708 (N_12708,N_11581,N_11745);
nand U12709 (N_12709,N_10741,N_11872);
or U12710 (N_12710,N_10894,N_11640);
and U12711 (N_12711,N_11833,N_11883);
nor U12712 (N_12712,N_11597,N_10968);
xor U12713 (N_12713,N_11563,N_10830);
and U12714 (N_12714,N_10765,N_11056);
xor U12715 (N_12715,N_10826,N_11224);
or U12716 (N_12716,N_10632,N_11501);
nand U12717 (N_12717,N_10931,N_11311);
xor U12718 (N_12718,N_11384,N_11775);
xnor U12719 (N_12719,N_10527,N_10731);
or U12720 (N_12720,N_11713,N_11416);
nand U12721 (N_12721,N_11189,N_11137);
or U12722 (N_12722,N_11154,N_10862);
nor U12723 (N_12723,N_10519,N_11280);
nand U12724 (N_12724,N_10935,N_10848);
xor U12725 (N_12725,N_11620,N_10533);
nand U12726 (N_12726,N_11684,N_11252);
and U12727 (N_12727,N_11627,N_10985);
or U12728 (N_12728,N_11330,N_10865);
or U12729 (N_12729,N_10501,N_11282);
nand U12730 (N_12730,N_10597,N_11549);
or U12731 (N_12731,N_10813,N_11109);
and U12732 (N_12732,N_10822,N_11525);
nor U12733 (N_12733,N_11434,N_10756);
or U12734 (N_12734,N_10773,N_11176);
nand U12735 (N_12735,N_11945,N_11223);
xor U12736 (N_12736,N_10604,N_11372);
nand U12737 (N_12737,N_10699,N_11341);
nor U12738 (N_12738,N_11036,N_11484);
xor U12739 (N_12739,N_10856,N_11340);
and U12740 (N_12740,N_11634,N_11931);
nand U12741 (N_12741,N_11606,N_10879);
nor U12742 (N_12742,N_11115,N_10946);
xnor U12743 (N_12743,N_10615,N_10864);
xor U12744 (N_12744,N_10895,N_10902);
nand U12745 (N_12745,N_11853,N_11573);
xnor U12746 (N_12746,N_10975,N_10600);
nor U12747 (N_12747,N_10700,N_10657);
and U12748 (N_12748,N_10984,N_10836);
nand U12749 (N_12749,N_10762,N_11342);
nor U12750 (N_12750,N_11230,N_11468);
nor U12751 (N_12751,N_10608,N_11297);
xnor U12752 (N_12752,N_11404,N_11476);
nand U12753 (N_12753,N_11539,N_11999);
nand U12754 (N_12754,N_10553,N_10748);
and U12755 (N_12755,N_11038,N_10716);
nand U12756 (N_12756,N_10616,N_11871);
nor U12757 (N_12757,N_11194,N_10580);
nand U12758 (N_12758,N_11027,N_11955);
and U12759 (N_12759,N_11203,N_11901);
and U12760 (N_12760,N_11264,N_11944);
or U12761 (N_12761,N_11482,N_10533);
xor U12762 (N_12762,N_11625,N_10554);
nor U12763 (N_12763,N_11324,N_11297);
or U12764 (N_12764,N_11812,N_11098);
and U12765 (N_12765,N_11509,N_10646);
xor U12766 (N_12766,N_10658,N_11156);
and U12767 (N_12767,N_11907,N_11421);
nor U12768 (N_12768,N_11300,N_11642);
and U12769 (N_12769,N_11386,N_11704);
and U12770 (N_12770,N_11121,N_10902);
xor U12771 (N_12771,N_10927,N_11335);
xnor U12772 (N_12772,N_11818,N_10788);
or U12773 (N_12773,N_11764,N_10634);
nand U12774 (N_12774,N_11103,N_11399);
and U12775 (N_12775,N_10556,N_11901);
and U12776 (N_12776,N_11802,N_10890);
nor U12777 (N_12777,N_11949,N_11467);
nor U12778 (N_12778,N_11409,N_10694);
and U12779 (N_12779,N_10682,N_11449);
and U12780 (N_12780,N_10717,N_11612);
xor U12781 (N_12781,N_11338,N_11427);
nand U12782 (N_12782,N_11595,N_10697);
and U12783 (N_12783,N_10881,N_11009);
and U12784 (N_12784,N_11483,N_10754);
nand U12785 (N_12785,N_11811,N_10906);
and U12786 (N_12786,N_10538,N_11218);
or U12787 (N_12787,N_11345,N_11323);
or U12788 (N_12788,N_10997,N_11616);
nand U12789 (N_12789,N_11515,N_11268);
nor U12790 (N_12790,N_11121,N_11767);
xor U12791 (N_12791,N_10619,N_11516);
xnor U12792 (N_12792,N_10669,N_11085);
or U12793 (N_12793,N_11758,N_11076);
or U12794 (N_12794,N_10682,N_10554);
nor U12795 (N_12795,N_10897,N_11310);
or U12796 (N_12796,N_11338,N_11104);
or U12797 (N_12797,N_10994,N_10516);
nor U12798 (N_12798,N_11960,N_11083);
nor U12799 (N_12799,N_10541,N_11591);
xnor U12800 (N_12800,N_11500,N_11033);
or U12801 (N_12801,N_10945,N_10531);
and U12802 (N_12802,N_11077,N_11982);
or U12803 (N_12803,N_10934,N_10790);
nand U12804 (N_12804,N_10695,N_11056);
xor U12805 (N_12805,N_11492,N_10679);
or U12806 (N_12806,N_11586,N_11121);
nand U12807 (N_12807,N_11468,N_11253);
nand U12808 (N_12808,N_11354,N_11326);
xnor U12809 (N_12809,N_11088,N_10529);
xnor U12810 (N_12810,N_11757,N_11032);
xnor U12811 (N_12811,N_11407,N_10702);
xor U12812 (N_12812,N_11005,N_11279);
nor U12813 (N_12813,N_11384,N_11429);
nor U12814 (N_12814,N_11483,N_11348);
or U12815 (N_12815,N_11927,N_11344);
nand U12816 (N_12816,N_11821,N_10559);
xnor U12817 (N_12817,N_10999,N_11046);
or U12818 (N_12818,N_11506,N_11988);
and U12819 (N_12819,N_10804,N_11581);
xor U12820 (N_12820,N_11805,N_10773);
xnor U12821 (N_12821,N_11957,N_11078);
nor U12822 (N_12822,N_10569,N_10766);
nor U12823 (N_12823,N_11176,N_10891);
nand U12824 (N_12824,N_11941,N_11793);
nand U12825 (N_12825,N_11781,N_11603);
xor U12826 (N_12826,N_10912,N_11340);
or U12827 (N_12827,N_11717,N_11658);
xnor U12828 (N_12828,N_10503,N_11124);
or U12829 (N_12829,N_11775,N_10643);
or U12830 (N_12830,N_11979,N_10720);
nor U12831 (N_12831,N_10687,N_10726);
nor U12832 (N_12832,N_11434,N_11909);
xnor U12833 (N_12833,N_11597,N_11562);
or U12834 (N_12834,N_11901,N_11748);
xnor U12835 (N_12835,N_11000,N_11892);
nor U12836 (N_12836,N_10587,N_11058);
nand U12837 (N_12837,N_10794,N_11846);
nand U12838 (N_12838,N_11798,N_11291);
nand U12839 (N_12839,N_10683,N_11996);
xnor U12840 (N_12840,N_11698,N_10955);
nor U12841 (N_12841,N_11686,N_10731);
or U12842 (N_12842,N_11407,N_11012);
nand U12843 (N_12843,N_11642,N_10879);
xor U12844 (N_12844,N_11449,N_11429);
xnor U12845 (N_12845,N_10806,N_10669);
nor U12846 (N_12846,N_10558,N_11580);
or U12847 (N_12847,N_11874,N_11989);
nor U12848 (N_12848,N_10565,N_11949);
nand U12849 (N_12849,N_11630,N_11979);
or U12850 (N_12850,N_10950,N_10965);
nand U12851 (N_12851,N_10597,N_11884);
nor U12852 (N_12852,N_11218,N_11104);
xor U12853 (N_12853,N_11104,N_10950);
xor U12854 (N_12854,N_10728,N_11729);
nor U12855 (N_12855,N_11073,N_10621);
and U12856 (N_12856,N_11211,N_11243);
xnor U12857 (N_12857,N_10977,N_11574);
and U12858 (N_12858,N_10556,N_10769);
xor U12859 (N_12859,N_11010,N_11392);
or U12860 (N_12860,N_10553,N_10830);
nor U12861 (N_12861,N_11255,N_10813);
and U12862 (N_12862,N_10719,N_10680);
and U12863 (N_12863,N_11800,N_10906);
nor U12864 (N_12864,N_10987,N_11235);
nand U12865 (N_12865,N_11175,N_11234);
nand U12866 (N_12866,N_11814,N_11115);
nor U12867 (N_12867,N_11191,N_11664);
and U12868 (N_12868,N_11410,N_10770);
and U12869 (N_12869,N_11509,N_11782);
and U12870 (N_12870,N_11167,N_11246);
xor U12871 (N_12871,N_10788,N_11683);
or U12872 (N_12872,N_10998,N_11724);
xnor U12873 (N_12873,N_10772,N_10614);
nor U12874 (N_12874,N_11419,N_11532);
xor U12875 (N_12875,N_10809,N_11589);
or U12876 (N_12876,N_11893,N_10634);
and U12877 (N_12877,N_11729,N_11124);
nor U12878 (N_12878,N_11095,N_11628);
nor U12879 (N_12879,N_11016,N_11269);
or U12880 (N_12880,N_11845,N_10960);
nor U12881 (N_12881,N_11814,N_11370);
nand U12882 (N_12882,N_10837,N_11767);
nor U12883 (N_12883,N_11399,N_11190);
nor U12884 (N_12884,N_11451,N_10697);
nand U12885 (N_12885,N_11846,N_11779);
xor U12886 (N_12886,N_10529,N_11064);
and U12887 (N_12887,N_11967,N_10878);
or U12888 (N_12888,N_10854,N_11536);
xor U12889 (N_12889,N_10765,N_11236);
nand U12890 (N_12890,N_11895,N_10772);
nand U12891 (N_12891,N_10648,N_11749);
and U12892 (N_12892,N_10559,N_10773);
xnor U12893 (N_12893,N_11837,N_11554);
xnor U12894 (N_12894,N_10651,N_11614);
or U12895 (N_12895,N_10931,N_10608);
or U12896 (N_12896,N_11460,N_11562);
nand U12897 (N_12897,N_11463,N_11869);
nor U12898 (N_12898,N_10715,N_11363);
xor U12899 (N_12899,N_11859,N_10934);
and U12900 (N_12900,N_11375,N_10959);
nand U12901 (N_12901,N_10666,N_11399);
and U12902 (N_12902,N_11556,N_11014);
nand U12903 (N_12903,N_11027,N_11950);
or U12904 (N_12904,N_11991,N_11450);
nor U12905 (N_12905,N_11015,N_11294);
xor U12906 (N_12906,N_11887,N_10728);
nand U12907 (N_12907,N_11633,N_11981);
nor U12908 (N_12908,N_10561,N_11522);
and U12909 (N_12909,N_11836,N_11145);
nor U12910 (N_12910,N_10691,N_11040);
xnor U12911 (N_12911,N_11310,N_11801);
or U12912 (N_12912,N_11067,N_11749);
and U12913 (N_12913,N_11662,N_10971);
nand U12914 (N_12914,N_10707,N_11296);
or U12915 (N_12915,N_11634,N_11502);
xnor U12916 (N_12916,N_11175,N_11140);
nand U12917 (N_12917,N_11955,N_11672);
nor U12918 (N_12918,N_11438,N_11114);
or U12919 (N_12919,N_10686,N_11498);
nand U12920 (N_12920,N_11209,N_11703);
or U12921 (N_12921,N_11405,N_10723);
nand U12922 (N_12922,N_10940,N_10946);
nor U12923 (N_12923,N_11873,N_10888);
nor U12924 (N_12924,N_11059,N_10500);
or U12925 (N_12925,N_11040,N_10704);
xnor U12926 (N_12926,N_10868,N_11832);
or U12927 (N_12927,N_10926,N_11241);
nand U12928 (N_12928,N_10731,N_11796);
nand U12929 (N_12929,N_11789,N_11935);
nor U12930 (N_12930,N_10733,N_11537);
nand U12931 (N_12931,N_11321,N_11285);
nand U12932 (N_12932,N_11804,N_10597);
nor U12933 (N_12933,N_11427,N_11801);
or U12934 (N_12934,N_11903,N_10665);
or U12935 (N_12935,N_11596,N_10899);
nand U12936 (N_12936,N_11220,N_11467);
xnor U12937 (N_12937,N_11111,N_11551);
nand U12938 (N_12938,N_10796,N_10896);
xor U12939 (N_12939,N_11829,N_11456);
and U12940 (N_12940,N_11094,N_11611);
and U12941 (N_12941,N_11106,N_11988);
xnor U12942 (N_12942,N_11473,N_11044);
and U12943 (N_12943,N_11089,N_11093);
and U12944 (N_12944,N_11323,N_10717);
or U12945 (N_12945,N_11379,N_11413);
xnor U12946 (N_12946,N_11059,N_10549);
nand U12947 (N_12947,N_10604,N_11393);
xor U12948 (N_12948,N_11779,N_11606);
xnor U12949 (N_12949,N_10761,N_10630);
nand U12950 (N_12950,N_10731,N_11908);
nand U12951 (N_12951,N_11664,N_11632);
nor U12952 (N_12952,N_11402,N_11199);
xnor U12953 (N_12953,N_11726,N_11105);
or U12954 (N_12954,N_11318,N_10596);
nor U12955 (N_12955,N_11919,N_11023);
xor U12956 (N_12956,N_10924,N_11367);
nor U12957 (N_12957,N_11106,N_11622);
nor U12958 (N_12958,N_11882,N_11264);
and U12959 (N_12959,N_11297,N_11174);
xnor U12960 (N_12960,N_11260,N_11460);
and U12961 (N_12961,N_11674,N_11745);
nand U12962 (N_12962,N_11077,N_10622);
nand U12963 (N_12963,N_10733,N_10679);
nand U12964 (N_12964,N_11507,N_11241);
nor U12965 (N_12965,N_10703,N_11243);
nand U12966 (N_12966,N_11568,N_11120);
and U12967 (N_12967,N_10793,N_10594);
or U12968 (N_12968,N_11284,N_11341);
and U12969 (N_12969,N_11378,N_11532);
nor U12970 (N_12970,N_11648,N_10789);
xor U12971 (N_12971,N_11869,N_11520);
xnor U12972 (N_12972,N_11099,N_10816);
nor U12973 (N_12973,N_10791,N_11341);
xor U12974 (N_12974,N_10557,N_11537);
nand U12975 (N_12975,N_11994,N_11540);
and U12976 (N_12976,N_11038,N_11679);
nand U12977 (N_12977,N_11659,N_11712);
and U12978 (N_12978,N_11003,N_11777);
nor U12979 (N_12979,N_11593,N_11355);
nor U12980 (N_12980,N_11828,N_10949);
or U12981 (N_12981,N_11878,N_11914);
and U12982 (N_12982,N_10882,N_10901);
xnor U12983 (N_12983,N_11419,N_11739);
nand U12984 (N_12984,N_10974,N_11602);
nand U12985 (N_12985,N_11353,N_11539);
nand U12986 (N_12986,N_11929,N_11047);
xnor U12987 (N_12987,N_10522,N_11858);
or U12988 (N_12988,N_11953,N_11531);
and U12989 (N_12989,N_10826,N_11544);
nor U12990 (N_12990,N_10898,N_11499);
or U12991 (N_12991,N_10616,N_11635);
xor U12992 (N_12992,N_11663,N_11687);
or U12993 (N_12993,N_11886,N_11032);
nand U12994 (N_12994,N_11994,N_11232);
nor U12995 (N_12995,N_10748,N_11177);
or U12996 (N_12996,N_11173,N_11328);
nor U12997 (N_12997,N_11838,N_11417);
or U12998 (N_12998,N_10589,N_11221);
nor U12999 (N_12999,N_10704,N_11982);
or U13000 (N_13000,N_10909,N_10544);
xor U13001 (N_13001,N_10956,N_10711);
nand U13002 (N_13002,N_11437,N_10897);
or U13003 (N_13003,N_11316,N_10601);
or U13004 (N_13004,N_11349,N_11621);
nand U13005 (N_13005,N_11645,N_11844);
or U13006 (N_13006,N_11038,N_11275);
nand U13007 (N_13007,N_11338,N_11671);
or U13008 (N_13008,N_11991,N_10582);
and U13009 (N_13009,N_10559,N_11595);
or U13010 (N_13010,N_10639,N_11427);
and U13011 (N_13011,N_11676,N_10606);
xnor U13012 (N_13012,N_10909,N_11707);
nand U13013 (N_13013,N_11040,N_11246);
or U13014 (N_13014,N_11119,N_11214);
nand U13015 (N_13015,N_11656,N_11598);
or U13016 (N_13016,N_11582,N_10568);
and U13017 (N_13017,N_11522,N_11100);
nand U13018 (N_13018,N_10578,N_10873);
nand U13019 (N_13019,N_11218,N_11949);
and U13020 (N_13020,N_11464,N_10559);
nand U13021 (N_13021,N_11765,N_10843);
and U13022 (N_13022,N_11463,N_11074);
nor U13023 (N_13023,N_11663,N_11169);
xor U13024 (N_13024,N_11042,N_11370);
and U13025 (N_13025,N_11363,N_10852);
nor U13026 (N_13026,N_11019,N_11157);
or U13027 (N_13027,N_11079,N_10609);
and U13028 (N_13028,N_11611,N_11801);
and U13029 (N_13029,N_10909,N_11844);
nand U13030 (N_13030,N_10571,N_11459);
xor U13031 (N_13031,N_11828,N_11043);
nor U13032 (N_13032,N_11307,N_11694);
nand U13033 (N_13033,N_11342,N_11501);
and U13034 (N_13034,N_11365,N_10637);
nor U13035 (N_13035,N_10608,N_11383);
and U13036 (N_13036,N_11228,N_10776);
or U13037 (N_13037,N_10606,N_11864);
xnor U13038 (N_13038,N_10817,N_10643);
or U13039 (N_13039,N_10631,N_11945);
or U13040 (N_13040,N_11259,N_11019);
nor U13041 (N_13041,N_11587,N_11419);
xnor U13042 (N_13042,N_11122,N_11288);
nor U13043 (N_13043,N_10557,N_11123);
or U13044 (N_13044,N_10943,N_11415);
nor U13045 (N_13045,N_11941,N_11400);
nor U13046 (N_13046,N_10911,N_10542);
nor U13047 (N_13047,N_11022,N_11691);
nor U13048 (N_13048,N_11880,N_11996);
xnor U13049 (N_13049,N_11031,N_10518);
and U13050 (N_13050,N_10709,N_10628);
nor U13051 (N_13051,N_11478,N_11324);
xor U13052 (N_13052,N_11794,N_11494);
xnor U13053 (N_13053,N_11449,N_11226);
and U13054 (N_13054,N_11784,N_10507);
nor U13055 (N_13055,N_11265,N_11560);
nand U13056 (N_13056,N_10996,N_10690);
nand U13057 (N_13057,N_10750,N_11149);
nor U13058 (N_13058,N_11175,N_10917);
or U13059 (N_13059,N_10765,N_11981);
or U13060 (N_13060,N_11876,N_10671);
xnor U13061 (N_13061,N_10680,N_11257);
nand U13062 (N_13062,N_10822,N_11857);
nor U13063 (N_13063,N_11856,N_11064);
xnor U13064 (N_13064,N_11564,N_11451);
or U13065 (N_13065,N_10912,N_11316);
nor U13066 (N_13066,N_10708,N_10982);
nand U13067 (N_13067,N_11720,N_11134);
or U13068 (N_13068,N_10957,N_11448);
nor U13069 (N_13069,N_10975,N_11034);
nor U13070 (N_13070,N_11508,N_11800);
xor U13071 (N_13071,N_11072,N_11099);
nor U13072 (N_13072,N_11105,N_11180);
xnor U13073 (N_13073,N_11307,N_11860);
xnor U13074 (N_13074,N_10820,N_11166);
nor U13075 (N_13075,N_11633,N_11862);
xor U13076 (N_13076,N_11003,N_11956);
nor U13077 (N_13077,N_10778,N_11308);
nor U13078 (N_13078,N_11681,N_10802);
or U13079 (N_13079,N_11075,N_10800);
or U13080 (N_13080,N_11779,N_11890);
nand U13081 (N_13081,N_11450,N_11750);
or U13082 (N_13082,N_11087,N_11048);
xor U13083 (N_13083,N_10662,N_10511);
xnor U13084 (N_13084,N_11910,N_10574);
or U13085 (N_13085,N_10620,N_10927);
nor U13086 (N_13086,N_11232,N_11121);
xnor U13087 (N_13087,N_11023,N_11581);
nand U13088 (N_13088,N_10878,N_11998);
or U13089 (N_13089,N_10607,N_11282);
and U13090 (N_13090,N_10525,N_10861);
and U13091 (N_13091,N_10536,N_10743);
nand U13092 (N_13092,N_11936,N_10987);
nand U13093 (N_13093,N_10849,N_10981);
nor U13094 (N_13094,N_11708,N_11261);
or U13095 (N_13095,N_11009,N_11112);
nor U13096 (N_13096,N_11120,N_10537);
xnor U13097 (N_13097,N_10560,N_11819);
or U13098 (N_13098,N_11912,N_10562);
xor U13099 (N_13099,N_10799,N_11440);
xnor U13100 (N_13100,N_10799,N_11386);
nor U13101 (N_13101,N_10868,N_11355);
or U13102 (N_13102,N_11804,N_10659);
and U13103 (N_13103,N_11118,N_10926);
nand U13104 (N_13104,N_11706,N_10941);
and U13105 (N_13105,N_10674,N_11076);
and U13106 (N_13106,N_11718,N_11059);
nand U13107 (N_13107,N_11069,N_11667);
xnor U13108 (N_13108,N_10685,N_10645);
nand U13109 (N_13109,N_10836,N_11611);
xor U13110 (N_13110,N_10750,N_10648);
nand U13111 (N_13111,N_11117,N_10724);
nand U13112 (N_13112,N_11040,N_11578);
nand U13113 (N_13113,N_11011,N_11397);
nand U13114 (N_13114,N_11463,N_10794);
and U13115 (N_13115,N_11864,N_11322);
nor U13116 (N_13116,N_11265,N_11341);
nor U13117 (N_13117,N_10875,N_11888);
or U13118 (N_13118,N_11869,N_11275);
xor U13119 (N_13119,N_11910,N_10506);
or U13120 (N_13120,N_11687,N_10716);
or U13121 (N_13121,N_11262,N_11424);
nand U13122 (N_13122,N_11262,N_11920);
or U13123 (N_13123,N_11186,N_10676);
nor U13124 (N_13124,N_11522,N_11176);
nand U13125 (N_13125,N_11614,N_11378);
nor U13126 (N_13126,N_10828,N_11337);
xnor U13127 (N_13127,N_11402,N_11753);
nand U13128 (N_13128,N_11196,N_10960);
and U13129 (N_13129,N_10558,N_10749);
xor U13130 (N_13130,N_11760,N_10900);
or U13131 (N_13131,N_11797,N_10592);
nand U13132 (N_13132,N_10553,N_10871);
nand U13133 (N_13133,N_10904,N_11533);
nand U13134 (N_13134,N_10739,N_11076);
xor U13135 (N_13135,N_11142,N_11472);
nor U13136 (N_13136,N_11142,N_11621);
or U13137 (N_13137,N_10500,N_11211);
or U13138 (N_13138,N_11393,N_10889);
nand U13139 (N_13139,N_11351,N_10522);
xnor U13140 (N_13140,N_11973,N_11959);
nand U13141 (N_13141,N_11309,N_11599);
nand U13142 (N_13142,N_11293,N_11564);
or U13143 (N_13143,N_11758,N_10918);
xnor U13144 (N_13144,N_10581,N_11878);
nand U13145 (N_13145,N_10576,N_10694);
nor U13146 (N_13146,N_11296,N_11872);
xor U13147 (N_13147,N_11683,N_11494);
nor U13148 (N_13148,N_11777,N_11813);
nand U13149 (N_13149,N_10800,N_11781);
xnor U13150 (N_13150,N_11310,N_11937);
nand U13151 (N_13151,N_11783,N_11851);
xor U13152 (N_13152,N_10570,N_10924);
nor U13153 (N_13153,N_11009,N_10810);
and U13154 (N_13154,N_11978,N_10636);
or U13155 (N_13155,N_10968,N_11396);
nor U13156 (N_13156,N_10762,N_11196);
nor U13157 (N_13157,N_11404,N_11570);
and U13158 (N_13158,N_11760,N_10687);
nand U13159 (N_13159,N_11711,N_10740);
nor U13160 (N_13160,N_10779,N_11243);
nor U13161 (N_13161,N_11270,N_10782);
nor U13162 (N_13162,N_10726,N_11145);
nand U13163 (N_13163,N_11477,N_11464);
and U13164 (N_13164,N_11629,N_11865);
or U13165 (N_13165,N_11328,N_10951);
xnor U13166 (N_13166,N_11434,N_10680);
nand U13167 (N_13167,N_11840,N_10649);
xnor U13168 (N_13168,N_11412,N_11550);
or U13169 (N_13169,N_11781,N_10825);
xnor U13170 (N_13170,N_11739,N_11789);
nor U13171 (N_13171,N_11652,N_11842);
nand U13172 (N_13172,N_10618,N_10522);
xnor U13173 (N_13173,N_10898,N_11476);
and U13174 (N_13174,N_11707,N_11982);
xnor U13175 (N_13175,N_11195,N_11712);
nor U13176 (N_13176,N_10884,N_10941);
xor U13177 (N_13177,N_11809,N_11693);
and U13178 (N_13178,N_11175,N_11534);
and U13179 (N_13179,N_11450,N_10827);
and U13180 (N_13180,N_11094,N_11123);
nor U13181 (N_13181,N_10530,N_11988);
xor U13182 (N_13182,N_11426,N_11959);
nor U13183 (N_13183,N_11293,N_11443);
xnor U13184 (N_13184,N_11081,N_11283);
nor U13185 (N_13185,N_10765,N_10843);
nor U13186 (N_13186,N_11821,N_11434);
xnor U13187 (N_13187,N_11623,N_10852);
nand U13188 (N_13188,N_10722,N_10849);
xor U13189 (N_13189,N_11784,N_11571);
nor U13190 (N_13190,N_11777,N_11231);
nand U13191 (N_13191,N_10687,N_11915);
xor U13192 (N_13192,N_10848,N_11135);
nor U13193 (N_13193,N_10685,N_11244);
nor U13194 (N_13194,N_11880,N_11369);
nor U13195 (N_13195,N_10848,N_11977);
nor U13196 (N_13196,N_11621,N_11223);
nor U13197 (N_13197,N_10731,N_10532);
xnor U13198 (N_13198,N_10849,N_11175);
or U13199 (N_13199,N_11867,N_11572);
xor U13200 (N_13200,N_11740,N_11583);
or U13201 (N_13201,N_11274,N_10599);
and U13202 (N_13202,N_11694,N_11186);
or U13203 (N_13203,N_11242,N_11982);
xnor U13204 (N_13204,N_10879,N_11739);
xnor U13205 (N_13205,N_10624,N_11068);
nor U13206 (N_13206,N_10891,N_11590);
or U13207 (N_13207,N_11108,N_10901);
xor U13208 (N_13208,N_11019,N_11954);
or U13209 (N_13209,N_10944,N_10952);
nor U13210 (N_13210,N_10829,N_11244);
xor U13211 (N_13211,N_11983,N_10887);
nand U13212 (N_13212,N_11529,N_11023);
xnor U13213 (N_13213,N_11461,N_11258);
nor U13214 (N_13214,N_11782,N_11956);
xnor U13215 (N_13215,N_11551,N_11163);
nor U13216 (N_13216,N_11344,N_10685);
and U13217 (N_13217,N_11180,N_11443);
or U13218 (N_13218,N_11528,N_11722);
xnor U13219 (N_13219,N_11679,N_10999);
nor U13220 (N_13220,N_11825,N_10714);
nor U13221 (N_13221,N_11164,N_11657);
and U13222 (N_13222,N_11630,N_11474);
nor U13223 (N_13223,N_11581,N_10759);
nor U13224 (N_13224,N_10925,N_10626);
nand U13225 (N_13225,N_11282,N_10816);
or U13226 (N_13226,N_11219,N_11875);
nor U13227 (N_13227,N_11162,N_11133);
xor U13228 (N_13228,N_11386,N_11080);
nand U13229 (N_13229,N_11934,N_11778);
xnor U13230 (N_13230,N_11094,N_10820);
xnor U13231 (N_13231,N_11697,N_11131);
and U13232 (N_13232,N_10508,N_11090);
nand U13233 (N_13233,N_11983,N_11780);
xnor U13234 (N_13234,N_11327,N_11151);
xnor U13235 (N_13235,N_11085,N_11067);
or U13236 (N_13236,N_11525,N_10757);
xnor U13237 (N_13237,N_11794,N_11121);
and U13238 (N_13238,N_10600,N_10560);
nor U13239 (N_13239,N_10673,N_11543);
or U13240 (N_13240,N_11816,N_10947);
and U13241 (N_13241,N_11244,N_10548);
nor U13242 (N_13242,N_10698,N_11168);
xnor U13243 (N_13243,N_11609,N_11923);
nand U13244 (N_13244,N_11057,N_11432);
xor U13245 (N_13245,N_11858,N_11230);
xor U13246 (N_13246,N_11128,N_11791);
nand U13247 (N_13247,N_10995,N_11329);
xnor U13248 (N_13248,N_11537,N_11981);
or U13249 (N_13249,N_11037,N_10924);
and U13250 (N_13250,N_11763,N_11988);
nand U13251 (N_13251,N_10639,N_11140);
xnor U13252 (N_13252,N_11731,N_11464);
nand U13253 (N_13253,N_10930,N_11658);
xnor U13254 (N_13254,N_11077,N_10603);
xor U13255 (N_13255,N_11150,N_11637);
or U13256 (N_13256,N_11176,N_11120);
nand U13257 (N_13257,N_11221,N_11846);
nor U13258 (N_13258,N_11016,N_10859);
nand U13259 (N_13259,N_11598,N_11051);
nor U13260 (N_13260,N_11766,N_11006);
nand U13261 (N_13261,N_10606,N_11536);
nor U13262 (N_13262,N_11592,N_11997);
xnor U13263 (N_13263,N_11753,N_11496);
or U13264 (N_13264,N_10821,N_10838);
and U13265 (N_13265,N_11982,N_10801);
xnor U13266 (N_13266,N_11013,N_11447);
xor U13267 (N_13267,N_11831,N_11959);
nand U13268 (N_13268,N_11057,N_11820);
or U13269 (N_13269,N_11330,N_11920);
and U13270 (N_13270,N_11893,N_11078);
and U13271 (N_13271,N_11824,N_11647);
nand U13272 (N_13272,N_11575,N_10863);
nand U13273 (N_13273,N_11665,N_11634);
and U13274 (N_13274,N_10662,N_11114);
and U13275 (N_13275,N_11467,N_10807);
xnor U13276 (N_13276,N_10790,N_10530);
nor U13277 (N_13277,N_10821,N_11326);
nor U13278 (N_13278,N_11162,N_11000);
and U13279 (N_13279,N_11969,N_10701);
nor U13280 (N_13280,N_11490,N_11500);
nand U13281 (N_13281,N_11606,N_10762);
or U13282 (N_13282,N_11942,N_10788);
nor U13283 (N_13283,N_11392,N_11522);
nand U13284 (N_13284,N_11008,N_11992);
xor U13285 (N_13285,N_11659,N_10847);
nor U13286 (N_13286,N_11140,N_11220);
and U13287 (N_13287,N_11737,N_11068);
or U13288 (N_13288,N_11575,N_10793);
and U13289 (N_13289,N_11390,N_11963);
xnor U13290 (N_13290,N_11322,N_11048);
nand U13291 (N_13291,N_10848,N_10918);
xor U13292 (N_13292,N_11164,N_11990);
nor U13293 (N_13293,N_10592,N_11107);
and U13294 (N_13294,N_11505,N_11474);
and U13295 (N_13295,N_11758,N_10879);
xor U13296 (N_13296,N_11444,N_11410);
and U13297 (N_13297,N_11309,N_10907);
nand U13298 (N_13298,N_11796,N_11011);
nor U13299 (N_13299,N_10895,N_11118);
xnor U13300 (N_13300,N_11308,N_11357);
xor U13301 (N_13301,N_11972,N_10897);
nor U13302 (N_13302,N_11860,N_10747);
and U13303 (N_13303,N_11089,N_11079);
xor U13304 (N_13304,N_11515,N_11661);
xor U13305 (N_13305,N_11062,N_11158);
nand U13306 (N_13306,N_10937,N_11729);
nor U13307 (N_13307,N_11182,N_10933);
xor U13308 (N_13308,N_10777,N_10616);
nor U13309 (N_13309,N_11505,N_11111);
nor U13310 (N_13310,N_11439,N_10939);
and U13311 (N_13311,N_10978,N_11876);
xor U13312 (N_13312,N_11456,N_10590);
nand U13313 (N_13313,N_11061,N_11983);
nand U13314 (N_13314,N_10675,N_11868);
xor U13315 (N_13315,N_11291,N_10811);
xnor U13316 (N_13316,N_11200,N_10879);
xnor U13317 (N_13317,N_11887,N_11722);
nor U13318 (N_13318,N_10792,N_11660);
and U13319 (N_13319,N_10886,N_10556);
or U13320 (N_13320,N_11805,N_11720);
and U13321 (N_13321,N_11464,N_11455);
xor U13322 (N_13322,N_11870,N_11142);
xor U13323 (N_13323,N_10514,N_11582);
and U13324 (N_13324,N_10912,N_11906);
and U13325 (N_13325,N_11194,N_11631);
and U13326 (N_13326,N_11993,N_11694);
and U13327 (N_13327,N_10850,N_11268);
nor U13328 (N_13328,N_11216,N_11519);
and U13329 (N_13329,N_11785,N_11535);
nor U13330 (N_13330,N_11916,N_11571);
nand U13331 (N_13331,N_11818,N_10802);
xnor U13332 (N_13332,N_11841,N_11204);
nand U13333 (N_13333,N_10660,N_10813);
nor U13334 (N_13334,N_11850,N_10519);
and U13335 (N_13335,N_11748,N_11634);
nand U13336 (N_13336,N_11386,N_10594);
xor U13337 (N_13337,N_10798,N_11074);
nor U13338 (N_13338,N_10968,N_11317);
nand U13339 (N_13339,N_11367,N_11659);
xor U13340 (N_13340,N_11620,N_11580);
nor U13341 (N_13341,N_11465,N_10646);
nor U13342 (N_13342,N_11794,N_10838);
nand U13343 (N_13343,N_11285,N_10954);
xor U13344 (N_13344,N_10983,N_10954);
or U13345 (N_13345,N_11266,N_11040);
or U13346 (N_13346,N_11225,N_11113);
xor U13347 (N_13347,N_11425,N_11824);
or U13348 (N_13348,N_11003,N_11541);
nor U13349 (N_13349,N_11940,N_11734);
or U13350 (N_13350,N_10708,N_11858);
nor U13351 (N_13351,N_11826,N_11294);
nand U13352 (N_13352,N_11409,N_11688);
nand U13353 (N_13353,N_11040,N_10835);
and U13354 (N_13354,N_11101,N_10571);
xnor U13355 (N_13355,N_11592,N_11664);
nor U13356 (N_13356,N_11333,N_10865);
nor U13357 (N_13357,N_11191,N_10833);
and U13358 (N_13358,N_11708,N_11879);
xnor U13359 (N_13359,N_10661,N_10848);
or U13360 (N_13360,N_10659,N_11085);
nor U13361 (N_13361,N_10523,N_11687);
or U13362 (N_13362,N_11269,N_10970);
or U13363 (N_13363,N_11062,N_11334);
nor U13364 (N_13364,N_11553,N_11316);
and U13365 (N_13365,N_11394,N_11265);
xnor U13366 (N_13366,N_10565,N_11367);
nand U13367 (N_13367,N_10670,N_10988);
xor U13368 (N_13368,N_11648,N_11660);
and U13369 (N_13369,N_11919,N_10952);
or U13370 (N_13370,N_11470,N_11634);
nand U13371 (N_13371,N_11469,N_11136);
nand U13372 (N_13372,N_10684,N_11382);
and U13373 (N_13373,N_11497,N_11802);
or U13374 (N_13374,N_11808,N_10734);
and U13375 (N_13375,N_11810,N_11990);
xnor U13376 (N_13376,N_11906,N_11059);
or U13377 (N_13377,N_11205,N_10968);
nand U13378 (N_13378,N_11127,N_10534);
nand U13379 (N_13379,N_10911,N_11556);
and U13380 (N_13380,N_10765,N_11732);
xor U13381 (N_13381,N_11010,N_11750);
nor U13382 (N_13382,N_11826,N_10522);
or U13383 (N_13383,N_11587,N_11925);
or U13384 (N_13384,N_11925,N_11146);
xnor U13385 (N_13385,N_11551,N_11216);
nor U13386 (N_13386,N_11506,N_11837);
xor U13387 (N_13387,N_11863,N_11920);
nand U13388 (N_13388,N_11289,N_11963);
nand U13389 (N_13389,N_11852,N_11692);
and U13390 (N_13390,N_10997,N_11611);
and U13391 (N_13391,N_10984,N_11047);
nor U13392 (N_13392,N_11734,N_10856);
nand U13393 (N_13393,N_11949,N_11906);
nand U13394 (N_13394,N_11931,N_11434);
or U13395 (N_13395,N_10516,N_11412);
xor U13396 (N_13396,N_11242,N_10847);
nand U13397 (N_13397,N_11367,N_11214);
or U13398 (N_13398,N_10595,N_11913);
or U13399 (N_13399,N_10546,N_11340);
xor U13400 (N_13400,N_11110,N_11492);
and U13401 (N_13401,N_10766,N_10555);
or U13402 (N_13402,N_10998,N_11236);
nor U13403 (N_13403,N_11674,N_11162);
nor U13404 (N_13404,N_11173,N_11547);
xnor U13405 (N_13405,N_11342,N_11465);
xor U13406 (N_13406,N_11344,N_11211);
nor U13407 (N_13407,N_11034,N_10982);
xor U13408 (N_13408,N_10682,N_11550);
nor U13409 (N_13409,N_11784,N_10531);
and U13410 (N_13410,N_10627,N_11410);
nor U13411 (N_13411,N_10698,N_11396);
nor U13412 (N_13412,N_11215,N_11893);
xnor U13413 (N_13413,N_11448,N_11265);
xnor U13414 (N_13414,N_11092,N_11205);
or U13415 (N_13415,N_11543,N_10939);
nor U13416 (N_13416,N_10913,N_11706);
or U13417 (N_13417,N_11921,N_11334);
xor U13418 (N_13418,N_10604,N_11401);
xor U13419 (N_13419,N_11944,N_10829);
xor U13420 (N_13420,N_11004,N_11704);
xnor U13421 (N_13421,N_11049,N_11388);
nor U13422 (N_13422,N_11690,N_11713);
and U13423 (N_13423,N_10601,N_11975);
nor U13424 (N_13424,N_10534,N_10832);
xor U13425 (N_13425,N_11611,N_11512);
xor U13426 (N_13426,N_11788,N_10877);
xor U13427 (N_13427,N_11255,N_11593);
xor U13428 (N_13428,N_11848,N_11371);
or U13429 (N_13429,N_11775,N_11123);
nand U13430 (N_13430,N_11880,N_10956);
xnor U13431 (N_13431,N_10604,N_11185);
and U13432 (N_13432,N_11539,N_10737);
or U13433 (N_13433,N_10536,N_11262);
and U13434 (N_13434,N_10715,N_10662);
or U13435 (N_13435,N_10914,N_11881);
nand U13436 (N_13436,N_11982,N_11878);
or U13437 (N_13437,N_11321,N_10901);
nand U13438 (N_13438,N_11330,N_11298);
or U13439 (N_13439,N_11014,N_10739);
or U13440 (N_13440,N_11880,N_11935);
or U13441 (N_13441,N_11081,N_11487);
or U13442 (N_13442,N_11840,N_11814);
and U13443 (N_13443,N_10508,N_11334);
xnor U13444 (N_13444,N_11074,N_11194);
nand U13445 (N_13445,N_11606,N_10587);
xnor U13446 (N_13446,N_11386,N_11788);
nand U13447 (N_13447,N_10853,N_10923);
nand U13448 (N_13448,N_10947,N_11062);
xor U13449 (N_13449,N_11487,N_10532);
or U13450 (N_13450,N_11918,N_11668);
xor U13451 (N_13451,N_11235,N_11689);
nor U13452 (N_13452,N_11823,N_11033);
and U13453 (N_13453,N_11031,N_10972);
and U13454 (N_13454,N_10712,N_10540);
or U13455 (N_13455,N_11206,N_11963);
and U13456 (N_13456,N_10691,N_10900);
nand U13457 (N_13457,N_10765,N_11824);
nor U13458 (N_13458,N_10638,N_11634);
nor U13459 (N_13459,N_11765,N_10848);
xnor U13460 (N_13460,N_11725,N_11952);
and U13461 (N_13461,N_11712,N_11696);
nand U13462 (N_13462,N_10590,N_10655);
and U13463 (N_13463,N_11760,N_10733);
and U13464 (N_13464,N_11463,N_11400);
and U13465 (N_13465,N_11971,N_10710);
nor U13466 (N_13466,N_11936,N_10627);
nor U13467 (N_13467,N_10645,N_11301);
nor U13468 (N_13468,N_11449,N_11078);
nor U13469 (N_13469,N_11976,N_11133);
xor U13470 (N_13470,N_10740,N_11867);
and U13471 (N_13471,N_11515,N_11240);
nor U13472 (N_13472,N_11205,N_10590);
and U13473 (N_13473,N_10626,N_11690);
xnor U13474 (N_13474,N_10842,N_11530);
xor U13475 (N_13475,N_11772,N_10733);
or U13476 (N_13476,N_10574,N_10937);
or U13477 (N_13477,N_11363,N_11654);
or U13478 (N_13478,N_11560,N_10716);
nor U13479 (N_13479,N_11957,N_10757);
nand U13480 (N_13480,N_10531,N_11184);
nor U13481 (N_13481,N_11330,N_11562);
nand U13482 (N_13482,N_11037,N_11305);
and U13483 (N_13483,N_10644,N_11750);
xnor U13484 (N_13484,N_10790,N_11000);
or U13485 (N_13485,N_10838,N_10578);
xor U13486 (N_13486,N_11327,N_11696);
or U13487 (N_13487,N_11129,N_11398);
and U13488 (N_13488,N_11396,N_11553);
xor U13489 (N_13489,N_11294,N_11531);
nor U13490 (N_13490,N_11137,N_11303);
nor U13491 (N_13491,N_11402,N_11482);
and U13492 (N_13492,N_10943,N_11134);
nand U13493 (N_13493,N_11567,N_11267);
and U13494 (N_13494,N_10543,N_10984);
nand U13495 (N_13495,N_11895,N_11208);
or U13496 (N_13496,N_10841,N_10815);
xnor U13497 (N_13497,N_10997,N_10703);
nand U13498 (N_13498,N_11270,N_11794);
nor U13499 (N_13499,N_10960,N_11757);
nand U13500 (N_13500,N_12776,N_12679);
nor U13501 (N_13501,N_13445,N_12630);
and U13502 (N_13502,N_12726,N_12376);
nand U13503 (N_13503,N_13465,N_12451);
nand U13504 (N_13504,N_12710,N_12764);
and U13505 (N_13505,N_12212,N_13377);
nor U13506 (N_13506,N_13493,N_12491);
xor U13507 (N_13507,N_12247,N_13091);
and U13508 (N_13508,N_12879,N_12463);
or U13509 (N_13509,N_13315,N_13177);
and U13510 (N_13510,N_13470,N_13454);
nand U13511 (N_13511,N_13074,N_12238);
nand U13512 (N_13512,N_12880,N_12772);
nand U13513 (N_13513,N_12915,N_12937);
and U13514 (N_13514,N_12081,N_12158);
nor U13515 (N_13515,N_12246,N_12171);
xor U13516 (N_13516,N_13239,N_12185);
xnor U13517 (N_13517,N_12154,N_13040);
nand U13518 (N_13518,N_12524,N_12893);
nand U13519 (N_13519,N_12333,N_12117);
and U13520 (N_13520,N_12616,N_12049);
nor U13521 (N_13521,N_12177,N_12912);
nor U13522 (N_13522,N_12973,N_12399);
nor U13523 (N_13523,N_12403,N_13310);
nand U13524 (N_13524,N_13477,N_12511);
or U13525 (N_13525,N_12291,N_12188);
xor U13526 (N_13526,N_13029,N_13007);
or U13527 (N_13527,N_13405,N_12671);
and U13528 (N_13528,N_13443,N_12900);
and U13529 (N_13529,N_12813,N_13487);
nand U13530 (N_13530,N_12766,N_12902);
nor U13531 (N_13531,N_13394,N_12221);
and U13532 (N_13532,N_13168,N_13042);
nor U13533 (N_13533,N_13233,N_12642);
xor U13534 (N_13534,N_13428,N_13408);
xor U13535 (N_13535,N_12295,N_12182);
and U13536 (N_13536,N_13367,N_13257);
nand U13537 (N_13537,N_12856,N_12311);
nand U13538 (N_13538,N_12480,N_12521);
nor U13539 (N_13539,N_13277,N_12738);
xnor U13540 (N_13540,N_12601,N_12901);
nor U13541 (N_13541,N_13237,N_13240);
or U13542 (N_13542,N_13137,N_12692);
or U13543 (N_13543,N_12280,N_13324);
or U13544 (N_13544,N_12819,N_12352);
or U13545 (N_13545,N_12120,N_13354);
nor U13546 (N_13546,N_13104,N_12839);
xnor U13547 (N_13547,N_13109,N_12509);
xor U13548 (N_13548,N_12674,N_12097);
or U13549 (N_13549,N_12771,N_12709);
nor U13550 (N_13550,N_12327,N_12217);
and U13551 (N_13551,N_12862,N_13182);
and U13552 (N_13552,N_13131,N_12818);
and U13553 (N_13553,N_12334,N_12335);
and U13554 (N_13554,N_12495,N_12932);
xor U13555 (N_13555,N_12331,N_13458);
and U13556 (N_13556,N_12066,N_13144);
xor U13557 (N_13557,N_12379,N_13245);
and U13558 (N_13558,N_12603,N_12696);
nor U13559 (N_13559,N_12223,N_12047);
xnor U13560 (N_13560,N_12040,N_13406);
nand U13561 (N_13561,N_13432,N_12474);
or U13562 (N_13562,N_12865,N_13398);
or U13563 (N_13563,N_12492,N_12014);
nand U13564 (N_13564,N_12790,N_13489);
or U13565 (N_13565,N_12211,N_12914);
nand U13566 (N_13566,N_12847,N_12557);
and U13567 (N_13567,N_12980,N_13474);
or U13568 (N_13568,N_13384,N_12949);
or U13569 (N_13569,N_12852,N_12091);
xnor U13570 (N_13570,N_12874,N_13490);
nor U13571 (N_13571,N_12001,N_12442);
or U13572 (N_13572,N_13356,N_12367);
or U13573 (N_13573,N_12168,N_13190);
or U13574 (N_13574,N_12791,N_12634);
nand U13575 (N_13575,N_12614,N_12271);
or U13576 (N_13576,N_13434,N_13393);
and U13577 (N_13577,N_12167,N_13056);
and U13578 (N_13578,N_12477,N_13385);
or U13579 (N_13579,N_13412,N_12476);
nor U13580 (N_13580,N_12964,N_12660);
nand U13581 (N_13581,N_12008,N_12998);
xnor U13582 (N_13582,N_12780,N_12868);
nand U13583 (N_13583,N_13279,N_13025);
nand U13584 (N_13584,N_12712,N_12782);
xnor U13585 (N_13585,N_13299,N_12861);
and U13586 (N_13586,N_13469,N_12121);
xnor U13587 (N_13587,N_13140,N_13455);
or U13588 (N_13588,N_12253,N_12454);
nand U13589 (N_13589,N_12808,N_12134);
or U13590 (N_13590,N_12722,N_12105);
nand U13591 (N_13591,N_13271,N_13323);
xnor U13592 (N_13592,N_12923,N_13147);
xnor U13593 (N_13593,N_13222,N_12456);
nand U13594 (N_13594,N_12213,N_13345);
nor U13595 (N_13595,N_12582,N_12200);
xor U13596 (N_13596,N_12360,N_12229);
nor U13597 (N_13597,N_12162,N_12377);
nor U13598 (N_13598,N_13159,N_12669);
or U13599 (N_13599,N_12199,N_12531);
nor U13600 (N_13600,N_13055,N_12163);
nor U13601 (N_13601,N_12827,N_12611);
and U13602 (N_13602,N_12542,N_13347);
nor U13603 (N_13603,N_12924,N_12760);
and U13604 (N_13604,N_12899,N_12686);
and U13605 (N_13605,N_13242,N_12954);
and U13606 (N_13606,N_12731,N_13484);
xor U13607 (N_13607,N_13423,N_12513);
nor U13608 (N_13608,N_13223,N_12962);
and U13609 (N_13609,N_12636,N_12984);
and U13610 (N_13610,N_12683,N_12386);
nand U13611 (N_13611,N_13246,N_12920);
and U13612 (N_13612,N_12708,N_12112);
nand U13613 (N_13613,N_12483,N_13352);
nor U13614 (N_13614,N_12801,N_12183);
nand U13615 (N_13615,N_13146,N_13273);
nor U13616 (N_13616,N_12210,N_12309);
xnor U13617 (N_13617,N_12036,N_13017);
nor U13618 (N_13618,N_12995,N_13250);
xnor U13619 (N_13619,N_12422,N_13107);
nand U13620 (N_13620,N_13337,N_13100);
nor U13621 (N_13621,N_12499,N_12882);
xnor U13622 (N_13622,N_13106,N_12059);
nor U13623 (N_13623,N_12665,N_12762);
or U13624 (N_13624,N_12979,N_13123);
or U13625 (N_13625,N_12944,N_12982);
nor U13626 (N_13626,N_13047,N_13411);
nor U13627 (N_13627,N_13036,N_12272);
xnor U13628 (N_13628,N_13339,N_13387);
nand U13629 (N_13629,N_12983,N_12314);
nand U13630 (N_13630,N_12942,N_12232);
or U13631 (N_13631,N_13480,N_12549);
and U13632 (N_13632,N_12872,N_12805);
and U13633 (N_13633,N_12651,N_13022);
nor U13634 (N_13634,N_12249,N_12481);
nand U13635 (N_13635,N_12437,N_12448);
nand U13636 (N_13636,N_12159,N_12149);
nor U13637 (N_13637,N_12080,N_12695);
nor U13638 (N_13638,N_12986,N_12054);
nor U13639 (N_13639,N_12967,N_12510);
or U13640 (N_13640,N_12089,N_12786);
nand U13641 (N_13641,N_13390,N_13117);
xor U13642 (N_13642,N_13000,N_13261);
or U13643 (N_13643,N_12888,N_13082);
or U13644 (N_13644,N_12673,N_13101);
or U13645 (N_13645,N_13202,N_12290);
nand U13646 (N_13646,N_12936,N_12627);
and U13647 (N_13647,N_12816,N_13181);
nand U13648 (N_13648,N_12435,N_12370);
xor U13649 (N_13649,N_13446,N_13050);
or U13650 (N_13650,N_12754,N_13062);
nor U13651 (N_13651,N_12490,N_12508);
nor U13652 (N_13652,N_12729,N_12341);
xnor U13653 (N_13653,N_12706,N_13197);
and U13654 (N_13654,N_12270,N_12560);
xnor U13655 (N_13655,N_12220,N_12802);
and U13656 (N_13656,N_12160,N_13355);
and U13657 (N_13657,N_12237,N_12599);
nor U13658 (N_13658,N_13450,N_13461);
nor U13659 (N_13659,N_13155,N_13012);
and U13660 (N_13660,N_13497,N_13176);
nand U13661 (N_13661,N_13189,N_12575);
xnor U13662 (N_13662,N_12714,N_13021);
nor U13663 (N_13663,N_12432,N_12610);
nand U13664 (N_13664,N_12767,N_12250);
xnor U13665 (N_13665,N_12606,N_12053);
or U13666 (N_13666,N_13068,N_12007);
xor U13667 (N_13667,N_12684,N_12356);
xor U13668 (N_13668,N_13110,N_13462);
and U13669 (N_13669,N_13327,N_13171);
and U13670 (N_13670,N_12812,N_12427);
xnor U13671 (N_13671,N_13172,N_13466);
nand U13672 (N_13672,N_12433,N_13481);
nand U13673 (N_13673,N_12548,N_12803);
xnor U13674 (N_13674,N_12324,N_12023);
nand U13675 (N_13675,N_12364,N_13067);
and U13676 (N_13676,N_12006,N_12544);
nand U13677 (N_13677,N_12903,N_13280);
nand U13678 (N_13678,N_12203,N_12359);
nand U13679 (N_13679,N_12688,N_13495);
nor U13680 (N_13680,N_12301,N_12534);
xor U13681 (N_13681,N_12296,N_13096);
or U13682 (N_13682,N_12394,N_12361);
nor U13683 (N_13683,N_13061,N_13275);
xnor U13684 (N_13684,N_13128,N_13429);
xnor U13685 (N_13685,N_12447,N_12953);
nand U13686 (N_13686,N_13369,N_13205);
nor U13687 (N_13687,N_12537,N_12886);
or U13688 (N_13688,N_13483,N_12648);
and U13689 (N_13689,N_12908,N_12116);
xor U13690 (N_13690,N_12822,N_12486);
nor U13691 (N_13691,N_13361,N_12743);
xor U13692 (N_13692,N_12419,N_13206);
or U13693 (N_13693,N_12877,N_12917);
xnor U13694 (N_13694,N_13213,N_13145);
or U13695 (N_13695,N_13449,N_12957);
nor U13696 (N_13696,N_13373,N_12532);
xnor U13697 (N_13697,N_13286,N_13396);
nor U13698 (N_13698,N_12000,N_12153);
or U13699 (N_13699,N_13203,N_12189);
nor U13700 (N_13700,N_12172,N_13169);
nor U13701 (N_13701,N_13456,N_12587);
nor U13702 (N_13702,N_12533,N_13416);
nor U13703 (N_13703,N_12104,N_12793);
and U13704 (N_13704,N_12191,N_12501);
or U13705 (N_13705,N_12411,N_12099);
or U13706 (N_13706,N_12292,N_12682);
nor U13707 (N_13707,N_12758,N_12863);
and U13708 (N_13708,N_12781,N_13249);
nand U13709 (N_13709,N_12798,N_12389);
nor U13710 (N_13710,N_13311,N_13251);
nand U13711 (N_13711,N_12538,N_12174);
xor U13712 (N_13712,N_12817,N_13312);
and U13713 (N_13713,N_13217,N_12430);
xor U13714 (N_13714,N_13350,N_12079);
and U13715 (N_13715,N_12670,N_13143);
xnor U13716 (N_13716,N_12343,N_12550);
nand U13717 (N_13717,N_13325,N_12909);
or U13718 (N_13718,N_12694,N_13424);
nor U13719 (N_13719,N_12315,N_12947);
nand U13720 (N_13720,N_13027,N_12933);
nor U13721 (N_13721,N_13116,N_12069);
or U13722 (N_13722,N_12680,N_12527);
nand U13723 (N_13723,N_12431,N_13016);
and U13724 (N_13724,N_12573,N_13316);
nor U13725 (N_13725,N_12558,N_12392);
or U13726 (N_13726,N_13289,N_12385);
or U13727 (N_13727,N_12308,N_12348);
nand U13728 (N_13728,N_13404,N_12146);
nor U13729 (N_13729,N_12244,N_12063);
nand U13730 (N_13730,N_12241,N_12702);
nor U13731 (N_13731,N_13329,N_13086);
xor U13732 (N_13732,N_12077,N_13248);
nand U13733 (N_13733,N_12485,N_12928);
nand U13734 (N_13734,N_12181,N_13302);
xnor U13735 (N_13735,N_12413,N_12208);
xor U13736 (N_13736,N_12952,N_12038);
xnor U13737 (N_13737,N_13340,N_12552);
and U13738 (N_13738,N_12316,N_12843);
nor U13739 (N_13739,N_12225,N_12259);
nand U13740 (N_13740,N_13122,N_13064);
nand U13741 (N_13741,N_12342,N_12029);
nand U13742 (N_13742,N_12581,N_12365);
nand U13743 (N_13743,N_13437,N_12417);
or U13744 (N_13744,N_13447,N_13431);
nor U13745 (N_13745,N_12161,N_12281);
or U13746 (N_13746,N_13183,N_12825);
nand U13747 (N_13747,N_12258,N_13113);
and U13748 (N_13748,N_12164,N_12974);
xor U13749 (N_13749,N_12997,N_12655);
or U13750 (N_13750,N_12494,N_12078);
xor U13751 (N_13751,N_12742,N_12590);
xnor U13752 (N_13752,N_12028,N_12337);
and U13753 (N_13753,N_13204,N_12592);
nor U13754 (N_13754,N_12283,N_13232);
or U13755 (N_13755,N_13051,N_12329);
nand U13756 (N_13756,N_12057,N_12500);
or U13757 (N_13757,N_12242,N_13180);
nor U13758 (N_13758,N_12133,N_13215);
nand U13759 (N_13759,N_12022,N_13414);
nor U13760 (N_13760,N_12834,N_12138);
or U13761 (N_13761,N_12551,N_12588);
nor U13762 (N_13762,N_12891,N_12777);
and U13763 (N_13763,N_12916,N_12815);
xnor U13764 (N_13764,N_12778,N_13003);
xor U13765 (N_13765,N_12958,N_13392);
and U13766 (N_13766,N_13342,N_12410);
xnor U13767 (N_13767,N_12058,N_13254);
nor U13768 (N_13768,N_13258,N_12773);
xnor U13769 (N_13769,N_13179,N_12678);
nand U13770 (N_13770,N_12248,N_12522);
or U13771 (N_13771,N_12140,N_13492);
and U13772 (N_13772,N_12721,N_12641);
xor U13773 (N_13773,N_12257,N_12535);
xnor U13774 (N_13774,N_12027,N_12689);
xnor U13775 (N_13775,N_12226,N_13139);
nand U13776 (N_13776,N_12113,N_13093);
nor U13777 (N_13777,N_12875,N_12111);
or U13778 (N_13778,N_13336,N_13089);
and U13779 (N_13779,N_13276,N_13148);
nand U13780 (N_13780,N_12514,N_12449);
nor U13781 (N_13781,N_12092,N_13372);
nand U13782 (N_13782,N_13207,N_13058);
nand U13783 (N_13783,N_12945,N_12012);
and U13784 (N_13784,N_13314,N_12589);
nor U13785 (N_13785,N_12128,N_12612);
and U13786 (N_13786,N_13192,N_13282);
nor U13787 (N_13787,N_13228,N_13072);
and U13788 (N_13788,N_12278,N_12647);
or U13789 (N_13789,N_12855,N_12889);
and U13790 (N_13790,N_12675,N_12026);
xor U13791 (N_13791,N_12993,N_12845);
and U13792 (N_13792,N_13442,N_12322);
xor U13793 (N_13793,N_13220,N_13191);
or U13794 (N_13794,N_12288,N_13209);
nand U13795 (N_13795,N_13344,N_13438);
nor U13796 (N_13796,N_13305,N_12123);
and U13797 (N_13797,N_12137,N_12262);
nand U13798 (N_13798,N_12130,N_12593);
nor U13799 (N_13799,N_12905,N_12347);
and U13800 (N_13800,N_12735,N_12646);
nor U13801 (N_13801,N_12934,N_12939);
xor U13802 (N_13802,N_12718,N_12975);
nand U13803 (N_13803,N_12373,N_13320);
xor U13804 (N_13804,N_13225,N_13391);
and U13805 (N_13805,N_12887,N_12010);
xnor U13806 (N_13806,N_12724,N_13125);
or U13807 (N_13807,N_12227,N_13317);
or U13808 (N_13808,N_13313,N_12520);
and U13809 (N_13809,N_13001,N_12369);
nand U13810 (N_13810,N_12717,N_12779);
and U13811 (N_13811,N_13409,N_13135);
nand U13812 (N_13812,N_12205,N_12629);
nand U13813 (N_13813,N_13138,N_12677);
and U13814 (N_13814,N_12615,N_12363);
xnor U13815 (N_13815,N_13368,N_12382);
and U13816 (N_13816,N_12401,N_12190);
xnor U13817 (N_13817,N_12372,N_12032);
nor U13818 (N_13818,N_12266,N_12693);
or U13819 (N_13819,N_12970,N_12326);
nor U13820 (N_13820,N_13141,N_12497);
nor U13821 (N_13821,N_12961,N_13063);
and U13822 (N_13822,N_12255,N_13039);
and U13823 (N_13823,N_12951,N_12635);
nor U13824 (N_13824,N_13076,N_13224);
nor U13825 (N_13825,N_13219,N_13362);
and U13826 (N_13826,N_13380,N_12775);
xnor U13827 (N_13827,N_12090,N_13366);
and U13828 (N_13828,N_12201,N_12384);
or U13829 (N_13829,N_12658,N_12263);
nand U13830 (N_13830,N_12977,N_13436);
or U13831 (N_13831,N_13208,N_12019);
nand U13832 (N_13832,N_12921,N_12016);
nor U13833 (N_13833,N_13023,N_13360);
xor U13834 (N_13834,N_12155,N_13243);
nand U13835 (N_13835,N_13266,N_13486);
or U13836 (N_13836,N_12734,N_13292);
or U13837 (N_13837,N_12306,N_13482);
or U13838 (N_13838,N_13126,N_12193);
nand U13839 (N_13839,N_13475,N_13186);
xor U13840 (N_13840,N_12186,N_12375);
nor U13841 (N_13841,N_12748,N_13170);
nor U13842 (N_13842,N_13468,N_12371);
and U13843 (N_13843,N_12725,N_13389);
or U13844 (N_13844,N_13085,N_12554);
xnor U13845 (N_13845,N_12453,N_12108);
or U13846 (N_13846,N_12571,N_13066);
nand U13847 (N_13847,N_12021,N_12799);
or U13848 (N_13848,N_12085,N_12374);
xor U13849 (N_13849,N_12992,N_12842);
xor U13850 (N_13850,N_13160,N_12062);
and U13851 (N_13851,N_12383,N_12340);
or U13852 (N_13852,N_12585,N_12956);
nand U13853 (N_13853,N_12289,N_13165);
and U13854 (N_13854,N_12700,N_13478);
nand U13855 (N_13855,N_13298,N_12763);
nor U13856 (N_13856,N_12114,N_13133);
nor U13857 (N_13857,N_12739,N_12755);
and U13858 (N_13858,N_12691,N_13151);
or U13859 (N_13859,N_12011,N_12857);
xor U13860 (N_13860,N_13473,N_12279);
or U13861 (N_13861,N_12765,N_13363);
nand U13862 (N_13862,N_12609,N_12598);
or U13863 (N_13863,N_12515,N_12713);
xor U13864 (N_13864,N_12506,N_12355);
or U13865 (N_13865,N_12661,N_13166);
nand U13866 (N_13866,N_13163,N_12656);
or U13867 (N_13867,N_12122,N_12434);
and U13868 (N_13868,N_12547,N_12037);
and U13869 (N_13869,N_12564,N_12142);
xnor U13870 (N_13870,N_13008,N_12539);
xnor U13871 (N_13871,N_12676,N_12621);
or U13872 (N_13872,N_13158,N_12837);
or U13873 (N_13873,N_12439,N_12395);
nand U13874 (N_13874,N_13400,N_12144);
nor U13875 (N_13875,N_13346,N_12003);
nand U13876 (N_13876,N_12666,N_13014);
or U13877 (N_13877,N_12475,N_12943);
xor U13878 (N_13878,N_12468,N_13041);
xnor U13879 (N_13879,N_12894,N_12990);
and U13880 (N_13880,N_12195,N_13262);
nand U13881 (N_13881,N_12633,N_12488);
and U13882 (N_13882,N_13498,N_13046);
nand U13883 (N_13883,N_13378,N_12745);
nand U13884 (N_13884,N_13453,N_12358);
nor U13885 (N_13885,N_12095,N_12366);
nor U13886 (N_13886,N_13118,N_12747);
nand U13887 (N_13887,N_13297,N_12789);
nor U13888 (N_13888,N_13244,N_12784);
nor U13889 (N_13889,N_12141,N_12645);
nand U13890 (N_13890,N_12800,N_12653);
xor U13891 (N_13891,N_12015,N_12096);
nor U13892 (N_13892,N_12406,N_12436);
nor U13893 (N_13893,N_12218,N_13081);
nor U13894 (N_13894,N_12867,N_13371);
and U13895 (N_13895,N_12804,N_12126);
nand U13896 (N_13896,N_12457,N_13494);
and U13897 (N_13897,N_13381,N_12197);
or U13898 (N_13898,N_12568,N_12440);
nor U13899 (N_13899,N_13334,N_13120);
xnor U13900 (N_13900,N_12004,N_12536);
nor U13901 (N_13901,N_12580,N_13349);
nor U13902 (N_13902,N_12344,N_13195);
xor U13903 (N_13903,N_12543,N_13149);
nand U13904 (N_13904,N_13175,N_13038);
nor U13905 (N_13905,N_12854,N_13005);
and U13906 (N_13906,N_12088,N_13032);
nor U13907 (N_13907,N_12354,N_12046);
nand U13908 (N_13908,N_12424,N_12649);
nand U13909 (N_13909,N_13059,N_12727);
xor U13910 (N_13910,N_12319,N_12728);
or U13911 (N_13911,N_12836,N_12397);
or U13912 (N_13912,N_12323,N_13167);
xor U13913 (N_13913,N_12198,N_12409);
xor U13914 (N_13914,N_12761,N_12050);
and U13915 (N_13915,N_13471,N_12751);
nand U13916 (N_13916,N_12178,N_12043);
and U13917 (N_13917,N_12873,N_13427);
or U13918 (N_13918,N_13294,N_13034);
nand U13919 (N_13919,N_12883,N_13296);
nand U13920 (N_13920,N_12576,N_13402);
nor U13921 (N_13921,N_12756,N_13370);
nor U13922 (N_13922,N_12657,N_12041);
nand U13923 (N_13923,N_12788,N_12446);
nor U13924 (N_13924,N_13395,N_13087);
and U13925 (N_13925,N_12192,N_12024);
nor U13926 (N_13926,N_13200,N_12482);
xnor U13927 (N_13927,N_12876,N_12444);
nand U13928 (N_13928,N_12018,N_12595);
nor U13929 (N_13929,N_13365,N_13364);
nand U13930 (N_13930,N_12740,N_13024);
or U13931 (N_13931,N_13084,N_12139);
nor U13932 (N_13932,N_12254,N_12732);
and U13933 (N_13933,N_13071,N_13425);
nor U13934 (N_13934,N_12643,N_12525);
nor U13935 (N_13935,N_13010,N_12084);
xnor U13936 (N_13936,N_12971,N_13013);
nor U13937 (N_13937,N_12807,N_12216);
nand U13938 (N_13938,N_13150,N_12968);
nand U13939 (N_13939,N_12898,N_12559);
xnor U13940 (N_13940,N_13173,N_12567);
nor U13941 (N_13941,N_12297,N_13353);
or U13942 (N_13942,N_12060,N_12512);
nand U13943 (N_13943,N_13057,N_12586);
and U13944 (N_13944,N_12849,N_12231);
and U13945 (N_13945,N_13335,N_12579);
nand U13946 (N_13946,N_12707,N_12002);
and U13947 (N_13947,N_12904,N_12505);
xnor U13948 (N_13948,N_12033,N_12907);
nand U13949 (N_13949,N_12787,N_12838);
xnor U13950 (N_13950,N_12166,N_13304);
or U13951 (N_13951,N_13226,N_12150);
nand U13952 (N_13952,N_13092,N_12770);
nand U13953 (N_13953,N_13083,N_13422);
and U13954 (N_13954,N_12067,N_12821);
or U13955 (N_13955,N_13070,N_12135);
nand U13956 (N_13956,N_13241,N_13121);
xor U13957 (N_13957,N_12276,N_13154);
or U13958 (N_13958,N_13460,N_12698);
nand U13959 (N_13959,N_13111,N_12380);
nor U13960 (N_13960,N_12562,N_12991);
nor U13961 (N_13961,N_12604,N_12737);
nand U13962 (N_13962,N_12034,N_12136);
nor U13963 (N_13963,N_12622,N_13090);
xnor U13964 (N_13964,N_12287,N_13374);
and U13965 (N_13965,N_13463,N_12602);
and U13966 (N_13966,N_12966,N_13193);
nor U13967 (N_13967,N_13102,N_12179);
nor U13968 (N_13968,N_12517,N_13383);
or U13969 (N_13969,N_12206,N_12273);
and U13970 (N_13970,N_12871,N_12769);
nand U13971 (N_13971,N_12031,N_12996);
xnor U13972 (N_13972,N_12072,N_12711);
xor U13973 (N_13973,N_12911,N_12093);
or U13974 (N_13974,N_12074,N_12608);
or U13975 (N_13975,N_12858,N_12701);
and U13976 (N_13976,N_12125,N_12890);
and U13977 (N_13977,N_13479,N_12526);
or U13978 (N_13978,N_13080,N_12425);
nand U13979 (N_13979,N_12407,N_12321);
xnor U13980 (N_13980,N_12357,N_13015);
nor U13981 (N_13981,N_13075,N_12180);
nor U13982 (N_13982,N_13263,N_13134);
xnor U13983 (N_13983,N_12420,N_12672);
nand U13984 (N_13984,N_13306,N_12809);
and U13985 (N_13985,N_13234,N_12631);
and U13986 (N_13986,N_12460,N_12083);
xnor U13987 (N_13987,N_12426,N_13221);
nor U13988 (N_13988,N_12269,N_13399);
or U13989 (N_13989,N_13351,N_12507);
and U13990 (N_13990,N_13114,N_12100);
nand U13991 (N_13991,N_13332,N_13035);
nand U13992 (N_13992,N_12349,N_12175);
or U13993 (N_13993,N_12594,N_12299);
and U13994 (N_13994,N_12294,N_12864);
nand U13995 (N_13995,N_13069,N_12502);
xnor U13996 (N_13996,N_12832,N_13295);
nand U13997 (N_13997,N_12565,N_12184);
or U13998 (N_13998,N_13132,N_13303);
or U13999 (N_13999,N_12009,N_12685);
nand U14000 (N_14000,N_12070,N_12039);
and U14001 (N_14001,N_12204,N_13287);
xnor U14002 (N_14002,N_13044,N_13285);
xnor U14003 (N_14003,N_12640,N_12277);
or U14004 (N_14004,N_13439,N_12236);
nor U14005 (N_14005,N_12256,N_12129);
and U14006 (N_14006,N_12267,N_13293);
nor U14007 (N_14007,N_12840,N_12624);
nor U14008 (N_14008,N_13229,N_13318);
xor U14009 (N_14009,N_13331,N_12963);
nor U14010 (N_14010,N_12013,N_12935);
and U14011 (N_14011,N_12398,N_13330);
and U14012 (N_14012,N_12844,N_13321);
or U14013 (N_14013,N_13417,N_12668);
and U14014 (N_14014,N_13230,N_12325);
or U14015 (N_14015,N_12332,N_12638);
and U14016 (N_14016,N_12496,N_13283);
xor U14017 (N_14017,N_12265,N_12307);
nand U14018 (N_14018,N_13020,N_12165);
nand U14019 (N_14019,N_13343,N_12071);
or U14020 (N_14020,N_12438,N_12268);
nor U14021 (N_14021,N_12351,N_12716);
nand U14022 (N_14022,N_12919,N_12393);
or U14023 (N_14023,N_12597,N_12429);
and U14024 (N_14024,N_13328,N_12469);
and U14025 (N_14025,N_12017,N_12170);
and U14026 (N_14026,N_12042,N_13157);
nand U14027 (N_14027,N_13185,N_12224);
nor U14028 (N_14028,N_12264,N_12148);
nor U14029 (N_14029,N_12487,N_12423);
and U14030 (N_14030,N_12626,N_12941);
and U14031 (N_14031,N_12312,N_13270);
nor U14032 (N_14032,N_13073,N_12402);
nor U14033 (N_14033,N_13476,N_12619);
nand U14034 (N_14034,N_12405,N_12994);
nand U14035 (N_14035,N_13018,N_13156);
nor U14036 (N_14036,N_12467,N_12985);
and U14037 (N_14037,N_12318,N_13333);
xor U14038 (N_14038,N_12304,N_12897);
nand U14039 (N_14039,N_12157,N_12662);
xnor U14040 (N_14040,N_12569,N_13199);
nand U14041 (N_14041,N_12082,N_12650);
nor U14042 (N_14042,N_13448,N_12330);
and U14043 (N_14043,N_12068,N_12052);
or U14044 (N_14044,N_12723,N_13174);
xnor U14045 (N_14045,N_13433,N_13359);
nor U14046 (N_14046,N_12044,N_12811);
nor U14047 (N_14047,N_12965,N_12131);
or U14048 (N_14048,N_12545,N_12878);
nor U14049 (N_14049,N_12418,N_13098);
and U14050 (N_14050,N_13326,N_13435);
and U14051 (N_14051,N_13290,N_13403);
or U14052 (N_14052,N_12613,N_12464);
or U14053 (N_14053,N_12783,N_12228);
xor U14054 (N_14054,N_12831,N_13264);
and U14055 (N_14055,N_12285,N_12404);
xnor U14056 (N_14056,N_13060,N_13397);
nand U14057 (N_14057,N_12681,N_12946);
and U14058 (N_14058,N_12313,N_12132);
and U14059 (N_14059,N_12086,N_12841);
nand U14060 (N_14060,N_13260,N_13218);
and U14061 (N_14061,N_12300,N_12194);
nor U14062 (N_14062,N_12151,N_12346);
and U14063 (N_14063,N_13124,N_12774);
or U14064 (N_14064,N_12336,N_12950);
and U14065 (N_14065,N_12350,N_13212);
xor U14066 (N_14066,N_12302,N_12215);
nand U14067 (N_14067,N_12570,N_13338);
xor U14068 (N_14068,N_12896,N_13028);
or U14069 (N_14069,N_12744,N_13009);
or U14070 (N_14070,N_13130,N_12455);
nor U14071 (N_14071,N_13194,N_12759);
or U14072 (N_14072,N_12637,N_12048);
or U14073 (N_14073,N_13187,N_13099);
and U14074 (N_14074,N_12103,N_13401);
and U14075 (N_14075,N_13247,N_12378);
nand U14076 (N_14076,N_13033,N_12233);
and U14077 (N_14077,N_13357,N_13054);
or U14078 (N_14078,N_12866,N_13037);
nand U14079 (N_14079,N_13485,N_13162);
xor U14080 (N_14080,N_12918,N_12320);
and U14081 (N_14081,N_12196,N_12927);
nand U14082 (N_14082,N_12541,N_12516);
nor U14083 (N_14083,N_12458,N_13004);
and U14084 (N_14084,N_12362,N_12390);
or U14085 (N_14085,N_12757,N_12959);
nand U14086 (N_14086,N_12929,N_12275);
xor U14087 (N_14087,N_12555,N_13201);
nand U14088 (N_14088,N_13152,N_12035);
xor U14089 (N_14089,N_13236,N_13211);
nand U14090 (N_14090,N_12623,N_12396);
and U14091 (N_14091,N_13136,N_12940);
and U14092 (N_14092,N_12885,N_12503);
and U14093 (N_14093,N_12219,N_12461);
or U14094 (N_14094,N_13030,N_13108);
and U14095 (N_14095,N_13472,N_13269);
xnor U14096 (N_14096,N_12110,N_12736);
nor U14097 (N_14097,N_12753,N_13272);
xnor U14098 (N_14098,N_13142,N_12504);
xor U14099 (N_14099,N_13415,N_13235);
nor U14100 (N_14100,N_13079,N_12387);
nor U14101 (N_14101,N_12605,N_12820);
xnor U14102 (N_14102,N_13413,N_13419);
nor U14103 (N_14103,N_12851,N_13119);
or U14104 (N_14104,N_12574,N_12388);
or U14105 (N_14105,N_12222,N_12797);
or U14106 (N_14106,N_12591,N_12690);
xor U14107 (N_14107,N_13255,N_12561);
nor U14108 (N_14108,N_12870,N_12830);
or U14109 (N_14109,N_13268,N_12261);
and U14110 (N_14110,N_13048,N_13031);
or U14111 (N_14111,N_12999,N_12910);
and U14112 (N_14112,N_13309,N_12972);
or U14113 (N_14113,N_13043,N_12230);
nor U14114 (N_14114,N_12214,N_12795);
or U14115 (N_14115,N_12750,N_12310);
or U14116 (N_14116,N_12715,N_12628);
nor U14117 (N_14117,N_13375,N_12796);
or U14118 (N_14118,N_13105,N_12260);
xnor U14119 (N_14119,N_12169,N_12282);
nand U14120 (N_14120,N_12906,N_12152);
nand U14121 (N_14121,N_12828,N_13386);
nand U14122 (N_14122,N_12752,N_12293);
nor U14123 (N_14123,N_12607,N_12540);
nand U14124 (N_14124,N_12835,N_12484);
nor U14125 (N_14125,N_12073,N_12465);
xor U14126 (N_14126,N_12566,N_12584);
and U14127 (N_14127,N_12005,N_13011);
nand U14128 (N_14128,N_12076,N_12639);
or U14129 (N_14129,N_13026,N_12826);
xor U14130 (N_14130,N_12452,N_12948);
and U14131 (N_14131,N_12466,N_12473);
nor U14132 (N_14132,N_12518,N_12098);
nor U14133 (N_14133,N_12338,N_12733);
xnor U14134 (N_14134,N_13358,N_13095);
nand U14135 (N_14135,N_12833,N_12529);
xnor U14136 (N_14136,N_13440,N_13452);
and U14137 (N_14137,N_13379,N_13002);
xnor U14138 (N_14138,N_12176,N_12412);
or U14139 (N_14139,N_12353,N_12644);
xor U14140 (N_14140,N_12768,N_12235);
xor U14141 (N_14141,N_12926,N_12583);
nand U14142 (N_14142,N_13284,N_12978);
xor U14143 (N_14143,N_12853,N_13227);
or U14144 (N_14144,N_13161,N_12345);
or U14145 (N_14145,N_12530,N_12704);
nor U14146 (N_14146,N_12450,N_13103);
nor U14147 (N_14147,N_12976,N_12470);
and U14148 (N_14148,N_13300,N_12284);
and U14149 (N_14149,N_12519,N_12075);
nor U14150 (N_14150,N_12719,N_12578);
and U14151 (N_14151,N_12055,N_12652);
nor U14152 (N_14152,N_13153,N_13265);
or U14153 (N_14153,N_13256,N_13307);
or U14154 (N_14154,N_12065,N_13006);
xnor U14155 (N_14155,N_13115,N_13278);
or U14156 (N_14156,N_13421,N_13499);
nor U14157 (N_14157,N_12955,N_12115);
or U14158 (N_14158,N_12303,N_12051);
and U14159 (N_14159,N_12869,N_12617);
nor U14160 (N_14160,N_12339,N_13094);
nor U14161 (N_14161,N_13322,N_12305);
and U14162 (N_14162,N_12119,N_13184);
and U14163 (N_14163,N_13291,N_12703);
xnor U14164 (N_14164,N_12523,N_12618);
nor U14165 (N_14165,N_13319,N_13019);
xnor U14166 (N_14166,N_12498,N_13097);
and U14167 (N_14167,N_13088,N_13459);
xor U14168 (N_14168,N_12025,N_12749);
nor U14169 (N_14169,N_13376,N_12145);
and U14170 (N_14170,N_12478,N_12416);
or U14171 (N_14171,N_12471,N_12730);
nor U14172 (N_14172,N_12118,N_13441);
nor U14173 (N_14173,N_12667,N_12892);
and U14174 (N_14174,N_12462,N_12859);
xnor U14175 (N_14175,N_12408,N_12699);
or U14176 (N_14176,N_13198,N_12988);
nand U14177 (N_14177,N_12445,N_13418);
xnor U14178 (N_14178,N_13488,N_12848);
nand U14179 (N_14179,N_12064,N_13281);
nor U14180 (N_14180,N_13467,N_12824);
nand U14181 (N_14181,N_12572,N_12600);
xnor U14182 (N_14182,N_12556,N_12931);
xnor U14183 (N_14183,N_12286,N_13252);
nor U14184 (N_14184,N_13231,N_12045);
nand U14185 (N_14185,N_12061,N_12687);
nor U14186 (N_14186,N_12596,N_12987);
nand U14187 (N_14187,N_12400,N_13259);
nand U14188 (N_14188,N_12298,N_12553);
xnor U14189 (N_14189,N_12846,N_13112);
nor U14190 (N_14190,N_12441,N_12391);
or U14191 (N_14191,N_13267,N_12654);
and U14192 (N_14192,N_13348,N_12632);
and U14193 (N_14193,N_12823,N_12546);
nand U14194 (N_14194,N_12020,N_13052);
or U14195 (N_14195,N_12925,N_12109);
or U14196 (N_14196,N_12317,N_13410);
or U14197 (N_14197,N_13420,N_12829);
xnor U14198 (N_14198,N_12107,N_12922);
or U14199 (N_14199,N_13457,N_13078);
and U14200 (N_14200,N_13444,N_12415);
nor U14201 (N_14201,N_12245,N_12697);
and U14202 (N_14202,N_12124,N_13274);
or U14203 (N_14203,N_13496,N_13388);
nor U14204 (N_14204,N_13045,N_12156);
nor U14205 (N_14205,N_13430,N_12792);
or U14206 (N_14206,N_12056,N_13053);
or U14207 (N_14207,N_13127,N_13216);
xnor U14208 (N_14208,N_12659,N_12806);
and U14209 (N_14209,N_12930,N_13308);
nor U14210 (N_14210,N_12094,N_13214);
or U14211 (N_14211,N_12106,N_12881);
nand U14212 (N_14212,N_13491,N_12030);
xnor U14213 (N_14213,N_12489,N_12664);
nor U14214 (N_14214,N_12421,N_12101);
xnor U14215 (N_14215,N_12850,N_12368);
or U14216 (N_14216,N_12810,N_13451);
and U14217 (N_14217,N_12969,N_12785);
xnor U14218 (N_14218,N_12663,N_12746);
nand U14219 (N_14219,N_13188,N_13301);
nand U14220 (N_14220,N_13238,N_12243);
nand U14221 (N_14221,N_12127,N_12251);
nand U14222 (N_14222,N_12240,N_12274);
nand U14223 (N_14223,N_13129,N_13407);
xor U14224 (N_14224,N_12479,N_12472);
and U14225 (N_14225,N_13341,N_12895);
nand U14226 (N_14226,N_12207,N_12860);
xor U14227 (N_14227,N_12381,N_12234);
and U14228 (N_14228,N_12720,N_12209);
and U14229 (N_14229,N_12884,N_13164);
nor U14230 (N_14230,N_12493,N_12741);
or U14231 (N_14231,N_12143,N_12102);
and U14232 (N_14232,N_13426,N_12443);
or U14233 (N_14233,N_13464,N_13196);
xnor U14234 (N_14234,N_13382,N_12428);
and U14235 (N_14235,N_12239,N_12981);
or U14236 (N_14236,N_13049,N_12625);
xnor U14237 (N_14237,N_12202,N_12620);
nor U14238 (N_14238,N_12459,N_12913);
nor U14239 (N_14239,N_13288,N_12328);
nor U14240 (N_14240,N_13210,N_12705);
xnor U14241 (N_14241,N_12147,N_13253);
or U14242 (N_14242,N_13077,N_12938);
nor U14243 (N_14243,N_12960,N_12794);
nor U14244 (N_14244,N_12414,N_12252);
and U14245 (N_14245,N_12563,N_12187);
xnor U14246 (N_14246,N_13178,N_12528);
and U14247 (N_14247,N_12989,N_12087);
nor U14248 (N_14248,N_13065,N_12814);
xnor U14249 (N_14249,N_12577,N_12173);
nand U14250 (N_14250,N_13150,N_12813);
or U14251 (N_14251,N_12358,N_12496);
and U14252 (N_14252,N_12884,N_12252);
and U14253 (N_14253,N_12446,N_13312);
or U14254 (N_14254,N_12480,N_12491);
nand U14255 (N_14255,N_12011,N_12975);
nor U14256 (N_14256,N_13464,N_12068);
xor U14257 (N_14257,N_13289,N_12672);
or U14258 (N_14258,N_12959,N_13361);
and U14259 (N_14259,N_12628,N_12946);
xor U14260 (N_14260,N_12373,N_12328);
or U14261 (N_14261,N_12016,N_13384);
xor U14262 (N_14262,N_12193,N_12910);
xnor U14263 (N_14263,N_12304,N_13119);
nor U14264 (N_14264,N_12346,N_12406);
nand U14265 (N_14265,N_13095,N_12956);
nand U14266 (N_14266,N_12975,N_12841);
nor U14267 (N_14267,N_12217,N_12845);
and U14268 (N_14268,N_12680,N_12266);
or U14269 (N_14269,N_12903,N_13072);
or U14270 (N_14270,N_13439,N_13068);
and U14271 (N_14271,N_12903,N_12160);
nor U14272 (N_14272,N_13474,N_13058);
xor U14273 (N_14273,N_13316,N_13448);
and U14274 (N_14274,N_13185,N_12150);
or U14275 (N_14275,N_12094,N_12634);
nand U14276 (N_14276,N_12875,N_13347);
xnor U14277 (N_14277,N_12258,N_13472);
or U14278 (N_14278,N_13025,N_12792);
and U14279 (N_14279,N_12053,N_13160);
and U14280 (N_14280,N_12039,N_12330);
and U14281 (N_14281,N_12867,N_12683);
and U14282 (N_14282,N_12518,N_12526);
xor U14283 (N_14283,N_12621,N_13059);
xor U14284 (N_14284,N_12579,N_13226);
nand U14285 (N_14285,N_12102,N_12041);
and U14286 (N_14286,N_12241,N_12983);
nand U14287 (N_14287,N_12262,N_12425);
or U14288 (N_14288,N_12411,N_13067);
or U14289 (N_14289,N_13388,N_13293);
xor U14290 (N_14290,N_12323,N_12763);
xnor U14291 (N_14291,N_12859,N_12360);
nor U14292 (N_14292,N_12750,N_13449);
and U14293 (N_14293,N_12668,N_12024);
nand U14294 (N_14294,N_12498,N_12397);
and U14295 (N_14295,N_12845,N_12498);
nor U14296 (N_14296,N_12581,N_12435);
nor U14297 (N_14297,N_12733,N_12828);
and U14298 (N_14298,N_12960,N_13265);
or U14299 (N_14299,N_12451,N_12036);
or U14300 (N_14300,N_13091,N_12538);
xor U14301 (N_14301,N_12161,N_12572);
or U14302 (N_14302,N_12071,N_13108);
nor U14303 (N_14303,N_12096,N_13244);
nand U14304 (N_14304,N_12917,N_12950);
nor U14305 (N_14305,N_12534,N_13409);
or U14306 (N_14306,N_12753,N_12876);
nand U14307 (N_14307,N_12831,N_13018);
and U14308 (N_14308,N_12356,N_12935);
xor U14309 (N_14309,N_12253,N_12501);
xnor U14310 (N_14310,N_12731,N_12763);
or U14311 (N_14311,N_12866,N_12206);
nand U14312 (N_14312,N_12632,N_12506);
nand U14313 (N_14313,N_12149,N_13406);
nand U14314 (N_14314,N_12308,N_12821);
xnor U14315 (N_14315,N_12498,N_13402);
xor U14316 (N_14316,N_12083,N_12867);
or U14317 (N_14317,N_12618,N_13207);
nand U14318 (N_14318,N_12074,N_12022);
and U14319 (N_14319,N_13077,N_13422);
nand U14320 (N_14320,N_12086,N_12598);
nand U14321 (N_14321,N_13019,N_12737);
xor U14322 (N_14322,N_12976,N_12926);
or U14323 (N_14323,N_12353,N_13475);
nor U14324 (N_14324,N_13413,N_12858);
and U14325 (N_14325,N_13495,N_12017);
xor U14326 (N_14326,N_13215,N_12087);
and U14327 (N_14327,N_13125,N_13071);
nor U14328 (N_14328,N_12102,N_12634);
and U14329 (N_14329,N_12975,N_12976);
and U14330 (N_14330,N_12812,N_13103);
nor U14331 (N_14331,N_12640,N_12602);
or U14332 (N_14332,N_12669,N_12171);
nor U14333 (N_14333,N_13417,N_12612);
xor U14334 (N_14334,N_13033,N_13417);
nand U14335 (N_14335,N_13460,N_12910);
nor U14336 (N_14336,N_12270,N_12531);
nand U14337 (N_14337,N_13062,N_13006);
nand U14338 (N_14338,N_12172,N_12765);
nor U14339 (N_14339,N_12810,N_13390);
nand U14340 (N_14340,N_12577,N_12396);
nand U14341 (N_14341,N_13420,N_12797);
or U14342 (N_14342,N_12477,N_12022);
and U14343 (N_14343,N_12685,N_13122);
nand U14344 (N_14344,N_12516,N_12408);
and U14345 (N_14345,N_13232,N_12329);
or U14346 (N_14346,N_13152,N_12314);
or U14347 (N_14347,N_12370,N_12938);
and U14348 (N_14348,N_12276,N_12667);
and U14349 (N_14349,N_12010,N_13062);
nand U14350 (N_14350,N_12576,N_12094);
or U14351 (N_14351,N_13081,N_12020);
and U14352 (N_14352,N_12672,N_12867);
and U14353 (N_14353,N_12830,N_12141);
nor U14354 (N_14354,N_12998,N_12457);
and U14355 (N_14355,N_12594,N_12483);
or U14356 (N_14356,N_13229,N_12077);
xor U14357 (N_14357,N_13111,N_12185);
xor U14358 (N_14358,N_12948,N_12295);
xor U14359 (N_14359,N_13389,N_13495);
or U14360 (N_14360,N_13304,N_13012);
nand U14361 (N_14361,N_12789,N_12819);
or U14362 (N_14362,N_13287,N_12543);
and U14363 (N_14363,N_12486,N_13372);
or U14364 (N_14364,N_13208,N_12425);
or U14365 (N_14365,N_13019,N_12695);
and U14366 (N_14366,N_12287,N_13117);
and U14367 (N_14367,N_12500,N_12503);
and U14368 (N_14368,N_12148,N_13471);
xnor U14369 (N_14369,N_13371,N_12615);
and U14370 (N_14370,N_13030,N_12130);
or U14371 (N_14371,N_12488,N_13202);
xor U14372 (N_14372,N_13171,N_12837);
xnor U14373 (N_14373,N_12485,N_12902);
xnor U14374 (N_14374,N_13086,N_13035);
or U14375 (N_14375,N_12523,N_12081);
xnor U14376 (N_14376,N_12333,N_13353);
nor U14377 (N_14377,N_12203,N_13181);
and U14378 (N_14378,N_12716,N_12720);
nand U14379 (N_14379,N_12909,N_13360);
or U14380 (N_14380,N_12025,N_12644);
xnor U14381 (N_14381,N_12373,N_12637);
or U14382 (N_14382,N_12903,N_12732);
nor U14383 (N_14383,N_12371,N_13374);
nand U14384 (N_14384,N_12630,N_12834);
or U14385 (N_14385,N_12275,N_13354);
nor U14386 (N_14386,N_13209,N_12147);
or U14387 (N_14387,N_13450,N_12104);
nand U14388 (N_14388,N_12303,N_13374);
or U14389 (N_14389,N_13131,N_12918);
and U14390 (N_14390,N_13477,N_13282);
nor U14391 (N_14391,N_13404,N_13302);
xnor U14392 (N_14392,N_12454,N_13030);
or U14393 (N_14393,N_13327,N_12444);
xnor U14394 (N_14394,N_12692,N_12684);
and U14395 (N_14395,N_13288,N_13089);
nand U14396 (N_14396,N_12425,N_12947);
xnor U14397 (N_14397,N_12865,N_12835);
and U14398 (N_14398,N_13499,N_12407);
xnor U14399 (N_14399,N_12498,N_12827);
nand U14400 (N_14400,N_12001,N_12680);
or U14401 (N_14401,N_12291,N_12501);
and U14402 (N_14402,N_12880,N_12055);
nor U14403 (N_14403,N_12992,N_12588);
nor U14404 (N_14404,N_13185,N_13019);
xnor U14405 (N_14405,N_12022,N_12282);
and U14406 (N_14406,N_12812,N_12556);
and U14407 (N_14407,N_13006,N_13459);
xnor U14408 (N_14408,N_12436,N_12214);
or U14409 (N_14409,N_13459,N_12118);
or U14410 (N_14410,N_12909,N_12838);
nor U14411 (N_14411,N_13084,N_13268);
xor U14412 (N_14412,N_12436,N_12983);
nor U14413 (N_14413,N_13180,N_12608);
nor U14414 (N_14414,N_12595,N_12126);
xor U14415 (N_14415,N_13319,N_12482);
or U14416 (N_14416,N_12778,N_13178);
nor U14417 (N_14417,N_12386,N_12119);
xnor U14418 (N_14418,N_12883,N_12712);
xor U14419 (N_14419,N_12475,N_12340);
nand U14420 (N_14420,N_12192,N_12521);
nand U14421 (N_14421,N_12870,N_12601);
nor U14422 (N_14422,N_12928,N_12950);
or U14423 (N_14423,N_12347,N_13304);
nor U14424 (N_14424,N_12324,N_13148);
and U14425 (N_14425,N_12230,N_12952);
nor U14426 (N_14426,N_12978,N_12530);
and U14427 (N_14427,N_12541,N_13157);
xnor U14428 (N_14428,N_12093,N_13171);
nand U14429 (N_14429,N_13113,N_13397);
nor U14430 (N_14430,N_12548,N_13413);
or U14431 (N_14431,N_13260,N_12450);
xor U14432 (N_14432,N_12867,N_12557);
or U14433 (N_14433,N_12237,N_12286);
xnor U14434 (N_14434,N_12267,N_12820);
xor U14435 (N_14435,N_13471,N_13247);
and U14436 (N_14436,N_13080,N_13014);
and U14437 (N_14437,N_12963,N_12458);
nor U14438 (N_14438,N_13199,N_12792);
nand U14439 (N_14439,N_13402,N_12005);
nor U14440 (N_14440,N_13491,N_13222);
and U14441 (N_14441,N_13415,N_12505);
xor U14442 (N_14442,N_12694,N_12065);
xnor U14443 (N_14443,N_13132,N_12986);
xnor U14444 (N_14444,N_13066,N_13123);
nor U14445 (N_14445,N_12945,N_12781);
xor U14446 (N_14446,N_12232,N_13120);
or U14447 (N_14447,N_12100,N_13047);
or U14448 (N_14448,N_12750,N_12719);
nor U14449 (N_14449,N_13206,N_12498);
or U14450 (N_14450,N_12347,N_12808);
and U14451 (N_14451,N_12678,N_12609);
and U14452 (N_14452,N_13031,N_13156);
and U14453 (N_14453,N_12298,N_12397);
nand U14454 (N_14454,N_12599,N_12710);
or U14455 (N_14455,N_12141,N_12399);
nand U14456 (N_14456,N_13138,N_12009);
nand U14457 (N_14457,N_13101,N_13278);
nor U14458 (N_14458,N_12083,N_12598);
or U14459 (N_14459,N_13316,N_12369);
nor U14460 (N_14460,N_12163,N_13377);
nor U14461 (N_14461,N_12778,N_12560);
or U14462 (N_14462,N_12775,N_12907);
xnor U14463 (N_14463,N_12244,N_12316);
or U14464 (N_14464,N_13408,N_12035);
nor U14465 (N_14465,N_12809,N_13484);
xnor U14466 (N_14466,N_12758,N_12899);
and U14467 (N_14467,N_12899,N_13291);
and U14468 (N_14468,N_13328,N_12614);
or U14469 (N_14469,N_12893,N_12648);
nor U14470 (N_14470,N_12245,N_12900);
xnor U14471 (N_14471,N_12346,N_12771);
nand U14472 (N_14472,N_13410,N_12476);
and U14473 (N_14473,N_13003,N_12067);
or U14474 (N_14474,N_12760,N_13345);
nand U14475 (N_14475,N_12711,N_12354);
and U14476 (N_14476,N_13235,N_13035);
nand U14477 (N_14477,N_13269,N_12600);
nor U14478 (N_14478,N_12040,N_12059);
and U14479 (N_14479,N_13283,N_12581);
or U14480 (N_14480,N_13238,N_12972);
nor U14481 (N_14481,N_12550,N_12968);
nor U14482 (N_14482,N_12794,N_12134);
or U14483 (N_14483,N_12861,N_12988);
and U14484 (N_14484,N_12061,N_12449);
nor U14485 (N_14485,N_12001,N_13145);
nor U14486 (N_14486,N_12229,N_13022);
or U14487 (N_14487,N_12789,N_13266);
xnor U14488 (N_14488,N_12228,N_13032);
nor U14489 (N_14489,N_12710,N_12718);
or U14490 (N_14490,N_13179,N_13106);
or U14491 (N_14491,N_12783,N_12131);
xnor U14492 (N_14492,N_12759,N_12163);
nor U14493 (N_14493,N_13206,N_12380);
and U14494 (N_14494,N_12216,N_13081);
or U14495 (N_14495,N_12488,N_12013);
nor U14496 (N_14496,N_12521,N_12625);
xor U14497 (N_14497,N_13212,N_12958);
nand U14498 (N_14498,N_13357,N_12962);
or U14499 (N_14499,N_13194,N_13101);
nor U14500 (N_14500,N_12077,N_12522);
xnor U14501 (N_14501,N_13346,N_12945);
nand U14502 (N_14502,N_12238,N_13309);
nor U14503 (N_14503,N_13130,N_12247);
nand U14504 (N_14504,N_12486,N_13439);
xor U14505 (N_14505,N_12271,N_12234);
and U14506 (N_14506,N_13199,N_12520);
nand U14507 (N_14507,N_12163,N_12421);
xnor U14508 (N_14508,N_12353,N_12227);
nand U14509 (N_14509,N_12430,N_12052);
xnor U14510 (N_14510,N_12957,N_13009);
nor U14511 (N_14511,N_13384,N_12629);
and U14512 (N_14512,N_12123,N_12912);
xnor U14513 (N_14513,N_12520,N_13214);
nor U14514 (N_14514,N_12900,N_12933);
nand U14515 (N_14515,N_13221,N_12090);
xnor U14516 (N_14516,N_12508,N_13282);
nor U14517 (N_14517,N_13135,N_13107);
or U14518 (N_14518,N_13292,N_12457);
and U14519 (N_14519,N_13309,N_12861);
xnor U14520 (N_14520,N_13396,N_12678);
nand U14521 (N_14521,N_13017,N_12836);
and U14522 (N_14522,N_12130,N_12150);
xnor U14523 (N_14523,N_12282,N_13124);
xor U14524 (N_14524,N_12441,N_12607);
xor U14525 (N_14525,N_13215,N_13316);
nor U14526 (N_14526,N_12573,N_12150);
xnor U14527 (N_14527,N_13340,N_13219);
nor U14528 (N_14528,N_13302,N_13260);
xnor U14529 (N_14529,N_13133,N_12865);
nand U14530 (N_14530,N_12335,N_13454);
or U14531 (N_14531,N_12345,N_13017);
xor U14532 (N_14532,N_12708,N_12255);
nor U14533 (N_14533,N_12854,N_12756);
and U14534 (N_14534,N_12911,N_12454);
or U14535 (N_14535,N_13156,N_13308);
xor U14536 (N_14536,N_12668,N_12680);
xor U14537 (N_14537,N_12540,N_13301);
xor U14538 (N_14538,N_12307,N_12561);
or U14539 (N_14539,N_12061,N_12316);
and U14540 (N_14540,N_12383,N_12364);
or U14541 (N_14541,N_12627,N_12027);
xor U14542 (N_14542,N_13205,N_13126);
nor U14543 (N_14543,N_13375,N_12568);
and U14544 (N_14544,N_12688,N_13429);
nor U14545 (N_14545,N_12516,N_13264);
and U14546 (N_14546,N_12485,N_12919);
and U14547 (N_14547,N_12232,N_12200);
xnor U14548 (N_14548,N_12599,N_12043);
xnor U14549 (N_14549,N_13090,N_12037);
and U14550 (N_14550,N_12194,N_13292);
xor U14551 (N_14551,N_12901,N_12027);
xor U14552 (N_14552,N_12018,N_12876);
nand U14553 (N_14553,N_13119,N_12789);
nor U14554 (N_14554,N_13204,N_13085);
and U14555 (N_14555,N_12551,N_13083);
nor U14556 (N_14556,N_12045,N_13077);
nand U14557 (N_14557,N_12506,N_13459);
and U14558 (N_14558,N_12502,N_12388);
and U14559 (N_14559,N_13043,N_12623);
xnor U14560 (N_14560,N_13326,N_12253);
nor U14561 (N_14561,N_12440,N_12891);
and U14562 (N_14562,N_12565,N_12876);
nand U14563 (N_14563,N_13146,N_12080);
xnor U14564 (N_14564,N_12912,N_12417);
nand U14565 (N_14565,N_12620,N_12398);
nor U14566 (N_14566,N_12742,N_12552);
nor U14567 (N_14567,N_12972,N_13434);
or U14568 (N_14568,N_13360,N_12636);
or U14569 (N_14569,N_12379,N_12182);
nor U14570 (N_14570,N_12066,N_12918);
and U14571 (N_14571,N_13443,N_12752);
or U14572 (N_14572,N_13478,N_12952);
nor U14573 (N_14573,N_12941,N_12449);
nor U14574 (N_14574,N_12598,N_13396);
nor U14575 (N_14575,N_13199,N_13139);
or U14576 (N_14576,N_13325,N_12407);
and U14577 (N_14577,N_13215,N_12676);
nor U14578 (N_14578,N_12964,N_12031);
xnor U14579 (N_14579,N_13185,N_12383);
xnor U14580 (N_14580,N_12466,N_12733);
and U14581 (N_14581,N_13228,N_13347);
nand U14582 (N_14582,N_12053,N_13168);
and U14583 (N_14583,N_12355,N_12491);
and U14584 (N_14584,N_13118,N_13007);
xor U14585 (N_14585,N_12703,N_13246);
or U14586 (N_14586,N_12370,N_12239);
xnor U14587 (N_14587,N_12232,N_12735);
and U14588 (N_14588,N_13283,N_12063);
nand U14589 (N_14589,N_12037,N_13172);
nand U14590 (N_14590,N_12423,N_12404);
or U14591 (N_14591,N_13448,N_12451);
or U14592 (N_14592,N_12764,N_12781);
nand U14593 (N_14593,N_12373,N_13096);
and U14594 (N_14594,N_13140,N_13439);
xnor U14595 (N_14595,N_12256,N_12907);
and U14596 (N_14596,N_12883,N_12099);
and U14597 (N_14597,N_13226,N_12580);
nand U14598 (N_14598,N_12543,N_12429);
and U14599 (N_14599,N_12304,N_12404);
nor U14600 (N_14600,N_12063,N_13284);
xor U14601 (N_14601,N_13320,N_12370);
and U14602 (N_14602,N_13161,N_13292);
and U14603 (N_14603,N_13307,N_13425);
or U14604 (N_14604,N_12298,N_13039);
or U14605 (N_14605,N_12729,N_12824);
xor U14606 (N_14606,N_12291,N_12387);
nor U14607 (N_14607,N_13254,N_13006);
or U14608 (N_14608,N_13229,N_12787);
nand U14609 (N_14609,N_13028,N_13026);
nor U14610 (N_14610,N_13319,N_12429);
and U14611 (N_14611,N_13198,N_13017);
or U14612 (N_14612,N_13215,N_12594);
and U14613 (N_14613,N_12128,N_13374);
xnor U14614 (N_14614,N_12682,N_13179);
nand U14615 (N_14615,N_13131,N_12178);
or U14616 (N_14616,N_12341,N_12318);
and U14617 (N_14617,N_12402,N_13245);
nand U14618 (N_14618,N_12028,N_12433);
xnor U14619 (N_14619,N_12014,N_12309);
and U14620 (N_14620,N_12881,N_13483);
or U14621 (N_14621,N_12011,N_13490);
nor U14622 (N_14622,N_12311,N_12711);
xnor U14623 (N_14623,N_12899,N_13028);
nand U14624 (N_14624,N_13346,N_13330);
or U14625 (N_14625,N_13367,N_13047);
and U14626 (N_14626,N_12628,N_12550);
nand U14627 (N_14627,N_12431,N_12564);
nor U14628 (N_14628,N_12385,N_12581);
nand U14629 (N_14629,N_12068,N_12139);
nor U14630 (N_14630,N_12650,N_12640);
nor U14631 (N_14631,N_12973,N_12059);
and U14632 (N_14632,N_13163,N_13441);
nand U14633 (N_14633,N_13312,N_12187);
nand U14634 (N_14634,N_12877,N_12832);
xnor U14635 (N_14635,N_12460,N_12020);
xnor U14636 (N_14636,N_12179,N_12738);
xnor U14637 (N_14637,N_12867,N_13408);
nand U14638 (N_14638,N_12273,N_13112);
nor U14639 (N_14639,N_12310,N_13166);
xor U14640 (N_14640,N_13470,N_12326);
and U14641 (N_14641,N_12202,N_12037);
nand U14642 (N_14642,N_12926,N_13293);
nand U14643 (N_14643,N_12790,N_12482);
nor U14644 (N_14644,N_12603,N_13013);
nand U14645 (N_14645,N_13212,N_12696);
nand U14646 (N_14646,N_12564,N_13354);
or U14647 (N_14647,N_13413,N_12427);
or U14648 (N_14648,N_12203,N_12014);
nor U14649 (N_14649,N_12621,N_13255);
nor U14650 (N_14650,N_12238,N_12099);
or U14651 (N_14651,N_12382,N_13070);
nor U14652 (N_14652,N_13260,N_12423);
xnor U14653 (N_14653,N_12540,N_12291);
or U14654 (N_14654,N_12549,N_13315);
xnor U14655 (N_14655,N_13024,N_12172);
or U14656 (N_14656,N_13424,N_13211);
and U14657 (N_14657,N_12880,N_13279);
nor U14658 (N_14658,N_13115,N_12029);
nor U14659 (N_14659,N_12101,N_13245);
nor U14660 (N_14660,N_12734,N_12748);
and U14661 (N_14661,N_13427,N_13291);
xor U14662 (N_14662,N_13417,N_13037);
nor U14663 (N_14663,N_12438,N_12533);
or U14664 (N_14664,N_13469,N_12372);
or U14665 (N_14665,N_13378,N_12223);
nor U14666 (N_14666,N_12974,N_12544);
xor U14667 (N_14667,N_12198,N_12001);
nor U14668 (N_14668,N_12420,N_13405);
xor U14669 (N_14669,N_12544,N_12160);
and U14670 (N_14670,N_12713,N_12970);
and U14671 (N_14671,N_12971,N_12177);
xor U14672 (N_14672,N_13082,N_12517);
nor U14673 (N_14673,N_12589,N_13433);
xor U14674 (N_14674,N_12436,N_12284);
and U14675 (N_14675,N_12339,N_13079);
nor U14676 (N_14676,N_12313,N_12304);
nand U14677 (N_14677,N_12560,N_12185);
xnor U14678 (N_14678,N_13486,N_12490);
nor U14679 (N_14679,N_12439,N_12309);
and U14680 (N_14680,N_13351,N_12784);
or U14681 (N_14681,N_13038,N_12068);
xor U14682 (N_14682,N_12399,N_12451);
or U14683 (N_14683,N_13421,N_12042);
nand U14684 (N_14684,N_13000,N_13240);
or U14685 (N_14685,N_13013,N_13494);
or U14686 (N_14686,N_12006,N_12171);
nor U14687 (N_14687,N_13381,N_12483);
nor U14688 (N_14688,N_12064,N_12431);
xor U14689 (N_14689,N_12770,N_13205);
and U14690 (N_14690,N_13324,N_13364);
nand U14691 (N_14691,N_12793,N_12399);
xnor U14692 (N_14692,N_12387,N_12184);
or U14693 (N_14693,N_12898,N_12619);
nand U14694 (N_14694,N_12508,N_12546);
xor U14695 (N_14695,N_12109,N_12445);
xor U14696 (N_14696,N_12906,N_13299);
or U14697 (N_14697,N_13283,N_12942);
nor U14698 (N_14698,N_12986,N_13222);
and U14699 (N_14699,N_12258,N_12334);
xor U14700 (N_14700,N_12633,N_12436);
and U14701 (N_14701,N_13431,N_12269);
or U14702 (N_14702,N_12117,N_12249);
or U14703 (N_14703,N_12061,N_13159);
nor U14704 (N_14704,N_12228,N_12537);
xnor U14705 (N_14705,N_12398,N_12107);
or U14706 (N_14706,N_12969,N_12001);
nor U14707 (N_14707,N_12241,N_12045);
nor U14708 (N_14708,N_12347,N_12556);
nand U14709 (N_14709,N_13326,N_12217);
or U14710 (N_14710,N_12323,N_12262);
and U14711 (N_14711,N_12251,N_12742);
xnor U14712 (N_14712,N_12556,N_13452);
xor U14713 (N_14713,N_12499,N_12014);
nand U14714 (N_14714,N_12290,N_13320);
nor U14715 (N_14715,N_12155,N_12985);
xor U14716 (N_14716,N_12490,N_12281);
nor U14717 (N_14717,N_12996,N_12899);
or U14718 (N_14718,N_13291,N_12606);
and U14719 (N_14719,N_12542,N_12483);
nand U14720 (N_14720,N_12437,N_12863);
and U14721 (N_14721,N_13227,N_12226);
xor U14722 (N_14722,N_13392,N_13260);
nor U14723 (N_14723,N_12712,N_12445);
xor U14724 (N_14724,N_12736,N_13259);
nand U14725 (N_14725,N_12097,N_12608);
and U14726 (N_14726,N_12030,N_13248);
xnor U14727 (N_14727,N_12255,N_12702);
and U14728 (N_14728,N_13059,N_12635);
nor U14729 (N_14729,N_13153,N_12397);
or U14730 (N_14730,N_12857,N_12719);
nor U14731 (N_14731,N_13050,N_13007);
nor U14732 (N_14732,N_12919,N_12477);
xor U14733 (N_14733,N_12105,N_13439);
xnor U14734 (N_14734,N_12104,N_13491);
nor U14735 (N_14735,N_12633,N_12611);
or U14736 (N_14736,N_13247,N_13287);
nand U14737 (N_14737,N_12006,N_12245);
or U14738 (N_14738,N_13489,N_12450);
and U14739 (N_14739,N_12326,N_13446);
and U14740 (N_14740,N_12246,N_13048);
nor U14741 (N_14741,N_13185,N_12675);
nor U14742 (N_14742,N_12965,N_12688);
and U14743 (N_14743,N_12322,N_13163);
or U14744 (N_14744,N_12230,N_12561);
xnor U14745 (N_14745,N_12996,N_12101);
and U14746 (N_14746,N_12993,N_13444);
or U14747 (N_14747,N_13340,N_13187);
and U14748 (N_14748,N_12566,N_13474);
and U14749 (N_14749,N_12446,N_13255);
and U14750 (N_14750,N_12261,N_12592);
nor U14751 (N_14751,N_13437,N_12849);
and U14752 (N_14752,N_12996,N_12449);
and U14753 (N_14753,N_13164,N_12176);
nor U14754 (N_14754,N_12655,N_13149);
nand U14755 (N_14755,N_12490,N_12014);
or U14756 (N_14756,N_12606,N_12035);
and U14757 (N_14757,N_12869,N_13280);
xor U14758 (N_14758,N_12141,N_13404);
nor U14759 (N_14759,N_12462,N_12932);
and U14760 (N_14760,N_12625,N_13312);
nand U14761 (N_14761,N_12119,N_12018);
nand U14762 (N_14762,N_13397,N_12821);
and U14763 (N_14763,N_12899,N_13206);
nor U14764 (N_14764,N_13167,N_12613);
or U14765 (N_14765,N_12116,N_12641);
nor U14766 (N_14766,N_12096,N_13195);
and U14767 (N_14767,N_13414,N_12962);
nand U14768 (N_14768,N_12451,N_12126);
and U14769 (N_14769,N_13181,N_13251);
or U14770 (N_14770,N_12816,N_12769);
and U14771 (N_14771,N_12072,N_13031);
xor U14772 (N_14772,N_13336,N_13278);
nand U14773 (N_14773,N_13479,N_12778);
or U14774 (N_14774,N_13449,N_12813);
and U14775 (N_14775,N_13301,N_13123);
or U14776 (N_14776,N_12529,N_13259);
nor U14777 (N_14777,N_12136,N_12798);
xnor U14778 (N_14778,N_13003,N_13208);
nor U14779 (N_14779,N_12330,N_12920);
and U14780 (N_14780,N_13146,N_12037);
or U14781 (N_14781,N_13016,N_13447);
nand U14782 (N_14782,N_12404,N_12803);
and U14783 (N_14783,N_13011,N_13272);
or U14784 (N_14784,N_12216,N_12452);
nor U14785 (N_14785,N_12863,N_13044);
and U14786 (N_14786,N_13093,N_12638);
or U14787 (N_14787,N_12604,N_12257);
xnor U14788 (N_14788,N_13366,N_13456);
nor U14789 (N_14789,N_13392,N_12637);
nor U14790 (N_14790,N_12210,N_12475);
and U14791 (N_14791,N_12772,N_12644);
nor U14792 (N_14792,N_12939,N_12455);
xor U14793 (N_14793,N_13000,N_12851);
and U14794 (N_14794,N_12596,N_12603);
nor U14795 (N_14795,N_12326,N_12474);
nor U14796 (N_14796,N_12917,N_12613);
and U14797 (N_14797,N_12565,N_12358);
xnor U14798 (N_14798,N_13039,N_13135);
xor U14799 (N_14799,N_13260,N_12111);
and U14800 (N_14800,N_13166,N_13104);
xor U14801 (N_14801,N_12850,N_12562);
nor U14802 (N_14802,N_13298,N_13276);
and U14803 (N_14803,N_13173,N_12488);
xnor U14804 (N_14804,N_12700,N_12431);
or U14805 (N_14805,N_12639,N_12331);
nor U14806 (N_14806,N_13380,N_13036);
nor U14807 (N_14807,N_13018,N_13056);
or U14808 (N_14808,N_12093,N_12097);
nand U14809 (N_14809,N_12355,N_13205);
nor U14810 (N_14810,N_12818,N_12714);
and U14811 (N_14811,N_13082,N_12199);
nor U14812 (N_14812,N_13401,N_12619);
and U14813 (N_14813,N_13301,N_13053);
nand U14814 (N_14814,N_12190,N_12980);
nand U14815 (N_14815,N_12216,N_12211);
nor U14816 (N_14816,N_12159,N_12656);
nand U14817 (N_14817,N_12085,N_12985);
nand U14818 (N_14818,N_13158,N_12027);
xor U14819 (N_14819,N_12515,N_12337);
or U14820 (N_14820,N_13110,N_13330);
xor U14821 (N_14821,N_12074,N_12994);
nand U14822 (N_14822,N_12381,N_12718);
or U14823 (N_14823,N_13329,N_13355);
or U14824 (N_14824,N_13309,N_12298);
or U14825 (N_14825,N_13443,N_12810);
or U14826 (N_14826,N_12925,N_12290);
and U14827 (N_14827,N_12907,N_12183);
and U14828 (N_14828,N_12484,N_12451);
and U14829 (N_14829,N_12977,N_12441);
xor U14830 (N_14830,N_13194,N_12743);
xnor U14831 (N_14831,N_12045,N_12688);
nand U14832 (N_14832,N_12179,N_12430);
or U14833 (N_14833,N_12890,N_12525);
or U14834 (N_14834,N_12205,N_12601);
or U14835 (N_14835,N_13329,N_13331);
and U14836 (N_14836,N_12776,N_12491);
nor U14837 (N_14837,N_12727,N_13243);
nor U14838 (N_14838,N_13212,N_12748);
or U14839 (N_14839,N_13344,N_12783);
nor U14840 (N_14840,N_12239,N_12582);
or U14841 (N_14841,N_13070,N_12377);
or U14842 (N_14842,N_13239,N_12375);
and U14843 (N_14843,N_12497,N_12918);
xnor U14844 (N_14844,N_12262,N_13150);
nand U14845 (N_14845,N_12641,N_12702);
xnor U14846 (N_14846,N_13461,N_13436);
and U14847 (N_14847,N_13044,N_13171);
nor U14848 (N_14848,N_13109,N_13178);
nor U14849 (N_14849,N_13038,N_12400);
or U14850 (N_14850,N_12439,N_12432);
and U14851 (N_14851,N_12071,N_13249);
or U14852 (N_14852,N_13009,N_12746);
xor U14853 (N_14853,N_12452,N_12178);
and U14854 (N_14854,N_12172,N_13336);
and U14855 (N_14855,N_12775,N_12204);
xor U14856 (N_14856,N_13202,N_13238);
xor U14857 (N_14857,N_13246,N_12338);
nand U14858 (N_14858,N_13107,N_12373);
xnor U14859 (N_14859,N_13317,N_12611);
xor U14860 (N_14860,N_12277,N_12409);
xnor U14861 (N_14861,N_12775,N_12685);
nand U14862 (N_14862,N_12598,N_13205);
and U14863 (N_14863,N_12610,N_12416);
and U14864 (N_14864,N_12518,N_12657);
or U14865 (N_14865,N_12621,N_12836);
xnor U14866 (N_14866,N_12325,N_12871);
nor U14867 (N_14867,N_12523,N_12806);
xnor U14868 (N_14868,N_13204,N_12121);
nand U14869 (N_14869,N_13134,N_13203);
nor U14870 (N_14870,N_13359,N_12881);
or U14871 (N_14871,N_12776,N_13116);
nor U14872 (N_14872,N_13199,N_12611);
xnor U14873 (N_14873,N_12973,N_13011);
xor U14874 (N_14874,N_13297,N_12984);
nor U14875 (N_14875,N_12659,N_12407);
nor U14876 (N_14876,N_12620,N_13468);
or U14877 (N_14877,N_12458,N_13159);
xor U14878 (N_14878,N_12335,N_13176);
xor U14879 (N_14879,N_13471,N_12201);
and U14880 (N_14880,N_13057,N_12541);
nor U14881 (N_14881,N_13153,N_13097);
or U14882 (N_14882,N_12040,N_13214);
and U14883 (N_14883,N_12351,N_13164);
and U14884 (N_14884,N_13421,N_12469);
xor U14885 (N_14885,N_12093,N_12545);
xor U14886 (N_14886,N_12951,N_12129);
nand U14887 (N_14887,N_12690,N_12073);
or U14888 (N_14888,N_12326,N_12776);
and U14889 (N_14889,N_12885,N_13313);
nor U14890 (N_14890,N_13293,N_13134);
xnor U14891 (N_14891,N_12140,N_12588);
nand U14892 (N_14892,N_12300,N_12036);
or U14893 (N_14893,N_12607,N_13004);
and U14894 (N_14894,N_12459,N_13332);
nor U14895 (N_14895,N_13233,N_12957);
or U14896 (N_14896,N_12845,N_12259);
nand U14897 (N_14897,N_13144,N_13172);
nor U14898 (N_14898,N_12911,N_12863);
or U14899 (N_14899,N_12313,N_13252);
and U14900 (N_14900,N_12214,N_12934);
xnor U14901 (N_14901,N_13088,N_12751);
or U14902 (N_14902,N_12078,N_12575);
xor U14903 (N_14903,N_12865,N_12861);
or U14904 (N_14904,N_12955,N_13006);
nor U14905 (N_14905,N_12314,N_13297);
nor U14906 (N_14906,N_12358,N_12684);
and U14907 (N_14907,N_12823,N_12037);
and U14908 (N_14908,N_12635,N_13126);
nor U14909 (N_14909,N_12432,N_12375);
and U14910 (N_14910,N_12757,N_12436);
nor U14911 (N_14911,N_12756,N_13255);
or U14912 (N_14912,N_12968,N_12777);
nand U14913 (N_14913,N_12769,N_13498);
nor U14914 (N_14914,N_12509,N_12475);
and U14915 (N_14915,N_12252,N_13489);
nor U14916 (N_14916,N_12821,N_12827);
xor U14917 (N_14917,N_13168,N_12970);
nor U14918 (N_14918,N_13220,N_13081);
nand U14919 (N_14919,N_12915,N_12172);
nor U14920 (N_14920,N_12406,N_12916);
or U14921 (N_14921,N_13228,N_13262);
and U14922 (N_14922,N_12814,N_12213);
xor U14923 (N_14923,N_12178,N_13268);
xor U14924 (N_14924,N_13230,N_12051);
or U14925 (N_14925,N_12194,N_12945);
nand U14926 (N_14926,N_12350,N_12638);
or U14927 (N_14927,N_12931,N_12673);
or U14928 (N_14928,N_12922,N_13302);
nand U14929 (N_14929,N_12634,N_12629);
nor U14930 (N_14930,N_13403,N_13223);
nand U14931 (N_14931,N_12774,N_13487);
or U14932 (N_14932,N_12618,N_12259);
nand U14933 (N_14933,N_13204,N_12267);
or U14934 (N_14934,N_12445,N_12847);
and U14935 (N_14935,N_12333,N_12091);
xnor U14936 (N_14936,N_12633,N_13484);
xor U14937 (N_14937,N_13201,N_13417);
or U14938 (N_14938,N_12632,N_13183);
and U14939 (N_14939,N_13286,N_13322);
or U14940 (N_14940,N_12444,N_12622);
nand U14941 (N_14941,N_13481,N_13144);
or U14942 (N_14942,N_12228,N_12963);
xnor U14943 (N_14943,N_12222,N_12123);
nand U14944 (N_14944,N_12874,N_13155);
nand U14945 (N_14945,N_12198,N_13381);
nor U14946 (N_14946,N_12669,N_12252);
or U14947 (N_14947,N_12770,N_13136);
nor U14948 (N_14948,N_13338,N_12361);
nand U14949 (N_14949,N_12299,N_13322);
xor U14950 (N_14950,N_13373,N_12391);
or U14951 (N_14951,N_13079,N_12319);
and U14952 (N_14952,N_13206,N_12122);
nand U14953 (N_14953,N_12527,N_12470);
xnor U14954 (N_14954,N_13279,N_13486);
nor U14955 (N_14955,N_13227,N_12873);
nor U14956 (N_14956,N_12956,N_12214);
or U14957 (N_14957,N_13351,N_12947);
xor U14958 (N_14958,N_12666,N_12366);
xor U14959 (N_14959,N_12905,N_12273);
nand U14960 (N_14960,N_12475,N_13365);
or U14961 (N_14961,N_13065,N_12237);
nand U14962 (N_14962,N_13370,N_12750);
and U14963 (N_14963,N_12537,N_12780);
and U14964 (N_14964,N_12681,N_12965);
xor U14965 (N_14965,N_12212,N_12057);
nor U14966 (N_14966,N_12132,N_13429);
and U14967 (N_14967,N_12695,N_13338);
and U14968 (N_14968,N_12059,N_12320);
and U14969 (N_14969,N_13219,N_12533);
nor U14970 (N_14970,N_13394,N_13357);
or U14971 (N_14971,N_13455,N_12733);
or U14972 (N_14972,N_12241,N_12611);
and U14973 (N_14973,N_12012,N_12168);
xnor U14974 (N_14974,N_13065,N_12993);
or U14975 (N_14975,N_12761,N_12918);
or U14976 (N_14976,N_12024,N_12112);
nor U14977 (N_14977,N_12254,N_13187);
nor U14978 (N_14978,N_12096,N_13309);
xor U14979 (N_14979,N_13144,N_12746);
and U14980 (N_14980,N_12675,N_12587);
and U14981 (N_14981,N_12912,N_13094);
xor U14982 (N_14982,N_13251,N_13133);
xor U14983 (N_14983,N_12681,N_13148);
and U14984 (N_14984,N_12316,N_12060);
nor U14985 (N_14985,N_12109,N_12213);
and U14986 (N_14986,N_13404,N_12926);
nor U14987 (N_14987,N_12421,N_13047);
xor U14988 (N_14988,N_12808,N_12581);
nand U14989 (N_14989,N_12283,N_13057);
nor U14990 (N_14990,N_12675,N_13118);
or U14991 (N_14991,N_12730,N_13437);
and U14992 (N_14992,N_12006,N_12068);
nor U14993 (N_14993,N_13166,N_12885);
and U14994 (N_14994,N_12497,N_13134);
and U14995 (N_14995,N_12271,N_12002);
or U14996 (N_14996,N_12212,N_12860);
nor U14997 (N_14997,N_12192,N_12299);
nand U14998 (N_14998,N_13147,N_12877);
nand U14999 (N_14999,N_12866,N_12779);
xnor UO_0 (O_0,N_13550,N_14147);
nor UO_1 (O_1,N_13741,N_14342);
or UO_2 (O_2,N_14350,N_13785);
and UO_3 (O_3,N_14826,N_14849);
nand UO_4 (O_4,N_14365,N_13592);
nand UO_5 (O_5,N_14320,N_13889);
xor UO_6 (O_6,N_14260,N_14156);
xor UO_7 (O_7,N_14123,N_13861);
nor UO_8 (O_8,N_14482,N_14374);
nor UO_9 (O_9,N_13723,N_14282);
nor UO_10 (O_10,N_14354,N_14872);
xnor UO_11 (O_11,N_13835,N_14939);
and UO_12 (O_12,N_14825,N_13912);
or UO_13 (O_13,N_14300,N_13990);
or UO_14 (O_14,N_14064,N_13583);
and UO_15 (O_15,N_13570,N_14929);
and UO_16 (O_16,N_14405,N_13679);
xnor UO_17 (O_17,N_13950,N_14540);
nand UO_18 (O_18,N_14041,N_13956);
nand UO_19 (O_19,N_13981,N_14583);
xor UO_20 (O_20,N_14544,N_13724);
or UO_21 (O_21,N_14148,N_14711);
or UO_22 (O_22,N_13585,N_13658);
and UO_23 (O_23,N_14690,N_14254);
nor UO_24 (O_24,N_14643,N_14670);
nand UO_25 (O_25,N_14718,N_14336);
and UO_26 (O_26,N_13574,N_14003);
nor UO_27 (O_27,N_13731,N_14833);
nand UO_28 (O_28,N_14289,N_13774);
or UO_29 (O_29,N_13817,N_13862);
nand UO_30 (O_30,N_14757,N_14664);
xor UO_31 (O_31,N_13729,N_14605);
and UO_32 (O_32,N_14580,N_13893);
nor UO_33 (O_33,N_13852,N_14774);
nor UO_34 (O_34,N_14706,N_14899);
and UO_35 (O_35,N_13984,N_14158);
nand UO_36 (O_36,N_13538,N_13790);
nor UO_37 (O_37,N_14674,N_14275);
nand UO_38 (O_38,N_14911,N_14961);
and UO_39 (O_39,N_14036,N_14351);
and UO_40 (O_40,N_14914,N_14904);
or UO_41 (O_41,N_14302,N_13680);
nand UO_42 (O_42,N_14235,N_14842);
nand UO_43 (O_43,N_14181,N_13962);
nor UO_44 (O_44,N_14986,N_14788);
and UO_45 (O_45,N_13930,N_14952);
or UO_46 (O_46,N_14109,N_14527);
xnor UO_47 (O_47,N_13725,N_14995);
xnor UO_48 (O_48,N_14547,N_14566);
xnor UO_49 (O_49,N_14010,N_14530);
nand UO_50 (O_50,N_14067,N_14874);
xnor UO_51 (O_51,N_13843,N_14283);
xnor UO_52 (O_52,N_14719,N_14061);
nor UO_53 (O_53,N_14864,N_14529);
or UO_54 (O_54,N_14733,N_14875);
xnor UO_55 (O_55,N_14345,N_14328);
xnor UO_56 (O_56,N_14212,N_14416);
nand UO_57 (O_57,N_14494,N_14548);
nand UO_58 (O_58,N_14198,N_14533);
nor UO_59 (O_59,N_14555,N_14829);
nor UO_60 (O_60,N_14075,N_14252);
nor UO_61 (O_61,N_13824,N_14159);
and UO_62 (O_62,N_13749,N_14411);
nor UO_63 (O_63,N_14209,N_14463);
and UO_64 (O_64,N_13779,N_14660);
xor UO_65 (O_65,N_13701,N_13672);
nor UO_66 (O_66,N_14388,N_14855);
nand UO_67 (O_67,N_14931,N_14110);
and UO_68 (O_68,N_13619,N_13839);
xnor UO_69 (O_69,N_14955,N_13595);
and UO_70 (O_70,N_13963,N_14713);
nand UO_71 (O_71,N_13863,N_14843);
and UO_72 (O_72,N_13961,N_14224);
nand UO_73 (O_73,N_13987,N_14907);
nand UO_74 (O_74,N_14989,N_14944);
nand UO_75 (O_75,N_13694,N_13593);
nor UO_76 (O_76,N_14069,N_14267);
and UO_77 (O_77,N_13949,N_14403);
nor UO_78 (O_78,N_13763,N_13503);
xnor UO_79 (O_79,N_14174,N_14753);
nand UO_80 (O_80,N_13581,N_14508);
xnor UO_81 (O_81,N_14293,N_14380);
or UO_82 (O_82,N_14065,N_14987);
xnor UO_83 (O_83,N_13911,N_13696);
xor UO_84 (O_84,N_14795,N_14606);
or UO_85 (O_85,N_13983,N_14701);
xor UO_86 (O_86,N_13744,N_13756);
xor UO_87 (O_87,N_13653,N_14358);
nand UO_88 (O_88,N_13666,N_13752);
nor UO_89 (O_89,N_13792,N_14838);
nand UO_90 (O_90,N_13746,N_14820);
nand UO_91 (O_91,N_13925,N_14404);
nand UO_92 (O_92,N_14216,N_13836);
and UO_93 (O_93,N_14432,N_14251);
nor UO_94 (O_94,N_13557,N_14349);
xor UO_95 (O_95,N_14692,N_14896);
xnor UO_96 (O_96,N_14563,N_14098);
and UO_97 (O_97,N_13762,N_13934);
nand UO_98 (O_98,N_14142,N_14621);
xor UO_99 (O_99,N_13565,N_14383);
xnor UO_100 (O_100,N_13998,N_13602);
and UO_101 (O_101,N_14290,N_14364);
or UO_102 (O_102,N_14005,N_13966);
xnor UO_103 (O_103,N_14766,N_14327);
xor UO_104 (O_104,N_14611,N_13936);
or UO_105 (O_105,N_14246,N_14515);
or UO_106 (O_106,N_13703,N_14756);
or UO_107 (O_107,N_14305,N_13829);
and UO_108 (O_108,N_13909,N_14724);
or UO_109 (O_109,N_13507,N_14568);
or UO_110 (O_110,N_14678,N_14011);
nand UO_111 (O_111,N_13767,N_14625);
and UO_112 (O_112,N_13657,N_14122);
xnor UO_113 (O_113,N_14071,N_14819);
or UO_114 (O_114,N_14748,N_13651);
or UO_115 (O_115,N_14448,N_14778);
nor UO_116 (O_116,N_13964,N_14296);
nand UO_117 (O_117,N_14916,N_14980);
xnor UO_118 (O_118,N_13778,N_14483);
nand UO_119 (O_119,N_13569,N_13900);
nor UO_120 (O_120,N_13627,N_14324);
and UO_121 (O_121,N_13868,N_14395);
or UO_122 (O_122,N_14006,N_14938);
nor UO_123 (O_123,N_13545,N_13504);
nor UO_124 (O_124,N_13944,N_13822);
nor UO_125 (O_125,N_13566,N_13562);
nand UO_126 (O_126,N_14867,N_14934);
nor UO_127 (O_127,N_14201,N_14593);
xor UO_128 (O_128,N_14859,N_14130);
nand UO_129 (O_129,N_14417,N_14306);
nor UO_130 (O_130,N_14789,N_13528);
xor UO_131 (O_131,N_14623,N_14474);
xor UO_132 (O_132,N_13548,N_14079);
nor UO_133 (O_133,N_13513,N_14090);
and UO_134 (O_134,N_14546,N_13572);
nand UO_135 (O_135,N_14612,N_14340);
or UO_136 (O_136,N_14759,N_14783);
nand UO_137 (O_137,N_14191,N_14108);
or UO_138 (O_138,N_14595,N_14465);
or UO_139 (O_139,N_14894,N_14173);
or UO_140 (O_140,N_14727,N_13973);
xnor UO_141 (O_141,N_14027,N_14832);
nand UO_142 (O_142,N_14433,N_13999);
or UO_143 (O_143,N_14900,N_13764);
nor UO_144 (O_144,N_14629,N_14967);
and UO_145 (O_145,N_14813,N_14261);
nand UO_146 (O_146,N_13618,N_14870);
nand UO_147 (O_147,N_13676,N_13643);
and UO_148 (O_148,N_13514,N_14263);
nor UO_149 (O_149,N_13877,N_13707);
nand UO_150 (O_150,N_14862,N_14725);
or UO_151 (O_151,N_14854,N_14019);
nor UO_152 (O_152,N_13979,N_14732);
nor UO_153 (O_153,N_13991,N_14384);
or UO_154 (O_154,N_14745,N_14406);
nand UO_155 (O_155,N_13727,N_14860);
or UO_156 (O_156,N_14182,N_14997);
or UO_157 (O_157,N_13649,N_13612);
xnor UO_158 (O_158,N_14419,N_13571);
or UO_159 (O_159,N_14648,N_14973);
nand UO_160 (O_160,N_14798,N_14343);
nor UO_161 (O_161,N_13568,N_14645);
or UO_162 (O_162,N_14062,N_14978);
and UO_163 (O_163,N_13804,N_14697);
nor UO_164 (O_164,N_14578,N_14150);
nand UO_165 (O_165,N_14205,N_14134);
and UO_166 (O_166,N_14428,N_14315);
xnor UO_167 (O_167,N_14236,N_14975);
nand UO_168 (O_168,N_14322,N_14219);
nor UO_169 (O_169,N_14603,N_14063);
nor UO_170 (O_170,N_14276,N_14074);
xnor UO_171 (O_171,N_13717,N_13512);
nor UO_172 (O_172,N_14534,N_14434);
and UO_173 (O_173,N_13831,N_14673);
nand UO_174 (O_174,N_14886,N_14392);
or UO_175 (O_175,N_14707,N_14966);
or UO_176 (O_176,N_14381,N_14225);
nand UO_177 (O_177,N_14023,N_14478);
nand UO_178 (O_178,N_13765,N_14423);
nor UO_179 (O_179,N_14704,N_13738);
nor UO_180 (O_180,N_13815,N_14270);
and UO_181 (O_181,N_14523,N_14379);
nand UO_182 (O_182,N_13630,N_14910);
nand UO_183 (O_183,N_14097,N_14279);
and UO_184 (O_184,N_13505,N_13806);
nor UO_185 (O_185,N_14880,N_14323);
or UO_186 (O_186,N_14335,N_13664);
and UO_187 (O_187,N_14585,N_13515);
or UO_188 (O_188,N_14743,N_14273);
or UO_189 (O_189,N_14895,N_14848);
xor UO_190 (O_190,N_14571,N_13748);
nand UO_191 (O_191,N_14565,N_14971);
and UO_192 (O_192,N_14991,N_13784);
nor UO_193 (O_193,N_13635,N_14758);
or UO_194 (O_194,N_13854,N_13549);
nor UO_195 (O_195,N_13770,N_13921);
and UO_196 (O_196,N_14081,N_14086);
and UO_197 (O_197,N_14947,N_13743);
and UO_198 (O_198,N_14425,N_14514);
and UO_199 (O_199,N_14893,N_13842);
nand UO_200 (O_200,N_14536,N_14981);
xor UO_201 (O_201,N_14356,N_13830);
nand UO_202 (O_202,N_14772,N_14815);
and UO_203 (O_203,N_14175,N_14538);
and UO_204 (O_204,N_14076,N_14339);
or UO_205 (O_205,N_14811,N_13637);
and UO_206 (O_206,N_13754,N_14835);
or UO_207 (O_207,N_13511,N_13985);
nand UO_208 (O_208,N_13786,N_14927);
nor UO_209 (O_209,N_13706,N_13888);
nand UO_210 (O_210,N_14171,N_13776);
xor UO_211 (O_211,N_14338,N_14087);
xnor UO_212 (O_212,N_14196,N_14146);
or UO_213 (O_213,N_14822,N_14072);
and UO_214 (O_214,N_14229,N_13808);
nand UO_215 (O_215,N_13878,N_14915);
and UO_216 (O_216,N_14637,N_13675);
or UO_217 (O_217,N_14232,N_14667);
and UO_218 (O_218,N_14988,N_14919);
nand UO_219 (O_219,N_13789,N_14321);
and UO_220 (O_220,N_14310,N_13918);
or UO_221 (O_221,N_13659,N_14227);
nand UO_222 (O_222,N_13782,N_14035);
xnor UO_223 (O_223,N_14769,N_14000);
xnor UO_224 (O_224,N_13768,N_13975);
or UO_225 (O_225,N_13642,N_14284);
xnor UO_226 (O_226,N_14999,N_14576);
and UO_227 (O_227,N_13965,N_14444);
and UO_228 (O_228,N_14785,N_13825);
or UO_229 (O_229,N_14857,N_14901);
or UO_230 (O_230,N_14741,N_14657);
nand UO_231 (O_231,N_13688,N_14599);
nand UO_232 (O_232,N_14627,N_14638);
xor UO_233 (O_233,N_14461,N_14303);
xnor UO_234 (O_234,N_13932,N_14326);
nor UO_235 (O_235,N_14683,N_14962);
xnor UO_236 (O_236,N_13536,N_13614);
nor UO_237 (O_237,N_14045,N_14972);
or UO_238 (O_238,N_14584,N_13544);
nor UO_239 (O_239,N_14165,N_13695);
and UO_240 (O_240,N_13584,N_13733);
nand UO_241 (O_241,N_14631,N_14168);
and UO_242 (O_242,N_14841,N_14178);
nand UO_243 (O_243,N_14172,N_14295);
and UO_244 (O_244,N_14518,N_13547);
nor UO_245 (O_245,N_14601,N_13908);
xor UO_246 (O_246,N_13628,N_14091);
nand UO_247 (O_247,N_14715,N_13941);
xor UO_248 (O_248,N_14736,N_14721);
xnor UO_249 (O_249,N_14133,N_13753);
nor UO_250 (O_250,N_14368,N_14332);
or UO_251 (O_251,N_14591,N_14389);
and UO_252 (O_252,N_14531,N_14945);
nand UO_253 (O_253,N_14837,N_14926);
or UO_254 (O_254,N_13606,N_13750);
or UO_255 (O_255,N_13891,N_14028);
nor UO_256 (O_256,N_13940,N_13976);
xnor UO_257 (O_257,N_14390,N_14528);
and UO_258 (O_258,N_14470,N_14702);
xor UO_259 (O_259,N_13787,N_13690);
xnor UO_260 (O_260,N_13794,N_14213);
nor UO_261 (O_261,N_14441,N_14865);
xor UO_262 (O_262,N_14139,N_14382);
or UO_263 (O_263,N_14477,N_14179);
xor UO_264 (O_264,N_14956,N_13638);
xnor UO_265 (O_265,N_14255,N_14426);
nor UO_266 (O_266,N_14614,N_13715);
xor UO_267 (O_267,N_14941,N_13874);
nor UO_268 (O_268,N_13736,N_13827);
or UO_269 (O_269,N_13541,N_13518);
nor UO_270 (O_270,N_13650,N_14370);
nand UO_271 (O_271,N_13948,N_14858);
xnor UO_272 (O_272,N_13864,N_14680);
nor UO_273 (O_273,N_14009,N_13834);
nand UO_274 (O_274,N_13919,N_14762);
xor UO_275 (O_275,N_14597,N_14298);
nor UO_276 (O_276,N_14633,N_13622);
nor UO_277 (O_277,N_14644,N_13957);
nand UO_278 (O_278,N_14656,N_14831);
xnor UO_279 (O_279,N_14497,N_13837);
nand UO_280 (O_280,N_14039,N_14024);
xor UO_281 (O_281,N_14669,N_14884);
nand UO_282 (O_282,N_14001,N_14163);
nor UO_283 (O_283,N_14472,N_13590);
and UO_284 (O_284,N_13751,N_14851);
or UO_285 (O_285,N_13886,N_14253);
xor UO_286 (O_286,N_14088,N_14113);
xnor UO_287 (O_287,N_14468,N_13561);
or UO_288 (O_288,N_14816,N_14008);
xnor UO_289 (O_289,N_14214,N_14963);
or UO_290 (O_290,N_14143,N_14983);
nand UO_291 (O_291,N_14511,N_14613);
or UO_292 (O_292,N_14476,N_13869);
or UO_293 (O_293,N_14455,N_13633);
xor UO_294 (O_294,N_13813,N_14698);
or UO_295 (O_295,N_13632,N_14622);
nor UO_296 (O_296,N_14266,N_13559);
nand UO_297 (O_297,N_14288,N_14723);
nand UO_298 (O_298,N_14693,N_13860);
or UO_299 (O_299,N_14722,N_14694);
nand UO_300 (O_300,N_14856,N_14830);
or UO_301 (O_301,N_13667,N_14249);
or UO_302 (O_302,N_14025,N_14866);
nor UO_303 (O_303,N_14887,N_14800);
and UO_304 (O_304,N_14687,N_13645);
nand UO_305 (O_305,N_13563,N_14539);
and UO_306 (O_306,N_14194,N_14125);
xor UO_307 (O_307,N_14046,N_14791);
xor UO_308 (O_308,N_14628,N_14121);
xor UO_309 (O_309,N_14850,N_13788);
and UO_310 (O_310,N_14532,N_13589);
nand UO_311 (O_311,N_14691,N_14094);
nor UO_312 (O_312,N_14211,N_13537);
nand UO_313 (O_313,N_14489,N_13755);
and UO_314 (O_314,N_13870,N_14127);
or UO_315 (O_315,N_13610,N_13519);
or UO_316 (O_316,N_13546,N_14132);
xnor UO_317 (O_317,N_13580,N_14863);
or UO_318 (O_318,N_13702,N_14869);
and UO_319 (O_319,N_14739,N_13989);
or UO_320 (O_320,N_13594,N_13578);
nand UO_321 (O_321,N_14786,N_13978);
nand UO_322 (O_322,N_13684,N_14281);
or UO_323 (O_323,N_13530,N_14274);
or UO_324 (O_324,N_13615,N_14602);
and UO_325 (O_325,N_14577,N_14215);
or UO_326 (O_326,N_13791,N_13579);
or UO_327 (O_327,N_14845,N_14562);
nand UO_328 (O_328,N_14188,N_14487);
xnor UO_329 (O_329,N_13895,N_13600);
and UO_330 (O_330,N_13904,N_14451);
nand UO_331 (O_331,N_13543,N_14760);
nor UO_332 (O_332,N_14953,N_14400);
nand UO_333 (O_333,N_14299,N_13661);
nor UO_334 (O_334,N_13654,N_14846);
xor UO_335 (O_335,N_14905,N_13847);
and UO_336 (O_336,N_14740,N_14466);
nor UO_337 (O_337,N_14427,N_14387);
or UO_338 (O_338,N_13714,N_14787);
or UO_339 (O_339,N_14550,N_14923);
xor UO_340 (O_340,N_13721,N_14458);
nor UO_341 (O_341,N_14844,N_13757);
nor UO_342 (O_342,N_14369,N_14549);
and UO_343 (O_343,N_14763,N_13691);
nor UO_344 (O_344,N_13665,N_13977);
xor UO_345 (O_345,N_14521,N_13995);
nor UO_346 (O_346,N_14709,N_13928);
nor UO_347 (O_347,N_13992,N_13634);
nor UO_348 (O_348,N_13802,N_14834);
nor UO_349 (O_349,N_14951,N_14506);
xnor UO_350 (O_350,N_13687,N_14898);
nand UO_351 (O_351,N_14101,N_14499);
nand UO_352 (O_352,N_14847,N_14582);
or UO_353 (O_353,N_13613,N_14446);
and UO_354 (O_354,N_14319,N_14516);
nor UO_355 (O_355,N_14840,N_14918);
and UO_356 (O_356,N_13971,N_14357);
nor UO_357 (O_357,N_13951,N_13742);
or UO_358 (O_358,N_13828,N_13849);
nor UO_359 (O_359,N_13508,N_14545);
nand UO_360 (O_360,N_14537,N_14280);
xnor UO_361 (O_361,N_13814,N_13556);
or UO_362 (O_362,N_14782,N_13532);
or UO_363 (O_363,N_14436,N_14728);
nor UO_364 (O_364,N_14137,N_13929);
nand UO_365 (O_365,N_14240,N_14022);
nand UO_366 (O_366,N_14111,N_13551);
xor UO_367 (O_367,N_14618,N_14187);
and UO_368 (O_368,N_13883,N_13996);
or UO_369 (O_369,N_14031,N_14735);
or UO_370 (O_370,N_14313,N_14177);
or UO_371 (O_371,N_14976,N_14512);
and UO_372 (O_372,N_13641,N_14592);
nand UO_373 (O_373,N_14202,N_13838);
nand UO_374 (O_374,N_13737,N_14341);
xnor UO_375 (O_375,N_13884,N_14943);
nor UO_376 (O_376,N_14647,N_14291);
nand UO_377 (O_377,N_14654,N_14239);
nand UO_378 (O_378,N_14491,N_13720);
xor UO_379 (O_379,N_13529,N_13960);
xnor UO_380 (O_380,N_14964,N_14457);
nor UO_381 (O_381,N_14102,N_14985);
nand UO_382 (O_382,N_14588,N_14309);
nand UO_383 (O_383,N_14292,N_14386);
nand UO_384 (O_384,N_13777,N_13783);
nand UO_385 (O_385,N_13599,N_14827);
nor UO_386 (O_386,N_13576,N_14112);
xnor UO_387 (O_387,N_13826,N_13531);
or UO_388 (O_388,N_14573,N_13509);
nand UO_389 (O_389,N_14556,N_14818);
nand UO_390 (O_390,N_14151,N_14821);
nand UO_391 (O_391,N_13734,N_14522);
nor UO_392 (O_392,N_14836,N_14207);
nand UO_393 (O_393,N_14128,N_13967);
nor UO_394 (O_394,N_14083,N_14804);
xor UO_395 (O_395,N_14594,N_13608);
or UO_396 (O_396,N_14708,N_14714);
xnor UO_397 (O_397,N_14402,N_13887);
nand UO_398 (O_398,N_14828,N_13501);
nand UO_399 (O_399,N_14761,N_14301);
xor UO_400 (O_400,N_14107,N_13697);
xnor UO_401 (O_401,N_14770,N_13876);
and UO_402 (O_402,N_13597,N_14703);
nor UO_403 (O_403,N_14913,N_14141);
xnor UO_404 (O_404,N_14093,N_13970);
or UO_405 (O_405,N_14218,N_14498);
or UO_406 (O_406,N_14180,N_14587);
or UO_407 (O_407,N_14567,N_14272);
or UO_408 (O_408,N_13502,N_14060);
xnor UO_409 (O_409,N_13739,N_13732);
nand UO_410 (O_410,N_13905,N_13994);
nor UO_411 (O_411,N_13718,N_14409);
and UO_412 (O_412,N_14259,N_14784);
or UO_413 (O_413,N_14812,N_14742);
nor UO_414 (O_414,N_14286,N_14334);
nor UO_415 (O_415,N_14641,N_13916);
or UO_416 (O_416,N_13626,N_13506);
nor UO_417 (O_417,N_14073,N_13517);
nand UO_418 (O_418,N_14959,N_13982);
nor UO_419 (O_419,N_14017,N_14230);
and UO_420 (O_420,N_13554,N_14208);
nor UO_421 (O_421,N_13914,N_14814);
and UO_422 (O_422,N_14192,N_14636);
and UO_423 (O_423,N_13685,N_13624);
or UO_424 (O_424,N_13605,N_14755);
nor UO_425 (O_425,N_14183,N_13577);
nand UO_426 (O_426,N_13972,N_14676);
or UO_427 (O_427,N_14940,N_14502);
nor UO_428 (O_428,N_14659,N_13534);
xnor UO_429 (O_429,N_14979,N_13609);
and UO_430 (O_430,N_14247,N_14467);
xnor UO_431 (O_431,N_14590,N_14412);
nor UO_432 (O_432,N_14294,N_14355);
xor UO_433 (O_433,N_14161,N_14688);
and UO_434 (O_434,N_14653,N_13866);
xnor UO_435 (O_435,N_13773,N_14505);
xnor UO_436 (O_436,N_14777,N_14485);
nor UO_437 (O_437,N_14089,N_14696);
or UO_438 (O_438,N_14554,N_14226);
xnor UO_439 (O_439,N_13616,N_14135);
or UO_440 (O_440,N_14600,N_14347);
nand UO_441 (O_441,N_13903,N_14100);
and UO_442 (O_442,N_13892,N_14195);
or UO_443 (O_443,N_13601,N_13698);
nand UO_444 (O_444,N_14776,N_14699);
xnor UO_445 (O_445,N_13699,N_13681);
xnor UO_446 (O_446,N_14439,N_14803);
nand UO_447 (O_447,N_13719,N_13907);
xor UO_448 (O_448,N_14047,N_13678);
or UO_449 (O_449,N_14105,N_14507);
nor UO_450 (O_450,N_13604,N_13625);
xor UO_451 (O_451,N_14095,N_14542);
xor UO_452 (O_452,N_14256,N_14807);
nand UO_453 (O_453,N_13939,N_14993);
nor UO_454 (O_454,N_14839,N_13758);
nand UO_455 (O_455,N_13598,N_14352);
nor UO_456 (O_456,N_14312,N_14903);
or UO_457 (O_457,N_13730,N_14375);
nand UO_458 (O_458,N_14797,N_14632);
or UO_459 (O_459,N_13882,N_13573);
or UO_460 (O_460,N_14262,N_14790);
and UO_461 (O_461,N_14026,N_13652);
nand UO_462 (O_462,N_13663,N_14131);
or UO_463 (O_463,N_14705,N_14331);
nand UO_464 (O_464,N_14948,N_14344);
xnor UO_465 (O_465,N_14459,N_14808);
nand UO_466 (O_466,N_14937,N_13823);
or UO_467 (O_467,N_14149,N_14169);
and UO_468 (O_468,N_13620,N_14435);
nand UO_469 (O_469,N_13709,N_14136);
or UO_470 (O_470,N_14124,N_14186);
and UO_471 (O_471,N_14360,N_14559);
and UO_472 (O_472,N_14220,N_14325);
xnor UO_473 (O_473,N_14579,N_14333);
nor UO_474 (O_474,N_13564,N_14033);
nor UO_475 (O_475,N_13558,N_14421);
nand UO_476 (O_476,N_14015,N_13587);
and UO_477 (O_477,N_14968,N_13582);
and UO_478 (O_478,N_13523,N_13901);
or UO_479 (O_479,N_13931,N_14243);
xor UO_480 (O_480,N_14116,N_14646);
nor UO_481 (O_481,N_14396,N_14391);
and UO_482 (O_482,N_14138,N_14484);
and UO_483 (O_483,N_14397,N_14932);
and UO_484 (O_484,N_14145,N_14367);
and UO_485 (O_485,N_14068,N_14604);
xor UO_486 (O_486,N_14608,N_13810);
or UO_487 (O_487,N_14413,N_14348);
nand UO_488 (O_488,N_13867,N_13716);
and UO_489 (O_489,N_14004,N_13910);
nor UO_490 (O_490,N_14596,N_13894);
and UO_491 (O_491,N_14233,N_13596);
nor UO_492 (O_492,N_14437,N_13588);
nor UO_493 (O_493,N_13811,N_13969);
xor UO_494 (O_494,N_13821,N_13692);
xnor UO_495 (O_495,N_14543,N_13591);
or UO_496 (O_496,N_14767,N_13670);
or UO_497 (O_497,N_13611,N_14630);
nand UO_498 (O_498,N_13683,N_14480);
nand UO_499 (O_499,N_13747,N_14385);
nand UO_500 (O_500,N_14949,N_14902);
nor UO_501 (O_501,N_14607,N_14077);
xnor UO_502 (O_502,N_14479,N_13816);
xor UO_503 (O_503,N_13803,N_14551);
or UO_504 (O_504,N_14021,N_13524);
or UO_505 (O_505,N_14889,N_13937);
xnor UO_506 (O_506,N_14311,N_13660);
and UO_507 (O_507,N_14754,N_14184);
nand UO_508 (O_508,N_14394,N_14969);
xor UO_509 (O_509,N_14040,N_14581);
nand UO_510 (O_510,N_14445,N_14809);
and UO_511 (O_511,N_14410,N_14558);
xnor UO_512 (O_512,N_13668,N_14525);
or UO_513 (O_513,N_14560,N_13872);
nor UO_514 (O_514,N_14720,N_13820);
nand UO_515 (O_515,N_14672,N_14731);
xor UO_516 (O_516,N_14935,N_14965);
and UO_517 (O_517,N_13525,N_14377);
xnor UO_518 (O_518,N_14883,N_14675);
and UO_519 (O_519,N_14199,N_14099);
and UO_520 (O_520,N_13974,N_13745);
nand UO_521 (O_521,N_14307,N_14450);
nand UO_522 (O_522,N_14399,N_13924);
or UO_523 (O_523,N_14710,N_14269);
xnor UO_524 (O_524,N_14737,N_13879);
nor UO_525 (O_525,N_14014,N_14624);
or UO_526 (O_526,N_14154,N_14030);
and UO_527 (O_527,N_14114,N_14126);
xnor UO_528 (O_528,N_14257,N_14185);
xnor UO_529 (O_529,N_14876,N_13769);
xor UO_530 (O_530,N_13796,N_14050);
xnor UO_531 (O_531,N_13942,N_13516);
nand UO_532 (O_532,N_14152,N_14176);
nand UO_533 (O_533,N_14059,N_14572);
or UO_534 (O_534,N_14885,N_13700);
nand UO_535 (O_535,N_13527,N_13959);
nor UO_536 (O_536,N_13922,N_14946);
xnor UO_537 (O_537,N_13902,N_13728);
nand UO_538 (O_538,N_14793,N_14689);
xor UO_539 (O_539,N_13677,N_14449);
nand UO_540 (O_540,N_13993,N_13759);
nor UO_541 (O_541,N_13906,N_13781);
xnor UO_542 (O_542,N_14553,N_14817);
and UO_543 (O_543,N_14258,N_14610);
nand UO_544 (O_544,N_14650,N_14574);
nor UO_545 (O_545,N_13710,N_13656);
or UO_546 (O_546,N_14401,N_13898);
or UO_547 (O_547,N_14129,N_14998);
nor UO_548 (O_548,N_13980,N_14626);
and UO_549 (O_549,N_13881,N_13801);
nor UO_550 (O_550,N_14881,N_13760);
or UO_551 (O_551,N_14044,N_14570);
and UO_552 (O_552,N_13819,N_14634);
or UO_553 (O_553,N_14695,N_14729);
nand UO_554 (O_554,N_14655,N_14048);
nand UO_555 (O_555,N_13832,N_13708);
xor UO_556 (O_556,N_14032,N_13521);
xor UO_557 (O_557,N_14373,N_14250);
or UO_558 (O_558,N_13935,N_14917);
or UO_559 (O_559,N_14658,N_13693);
or UO_560 (O_560,N_14277,N_14443);
and UO_561 (O_561,N_14304,N_14996);
nand UO_562 (O_562,N_14609,N_14203);
nand UO_563 (O_563,N_14712,N_13938);
nor UO_564 (O_564,N_14504,N_14771);
or UO_565 (O_565,N_14806,N_14888);
or UO_566 (O_566,N_14029,N_13812);
nor UO_567 (O_567,N_14287,N_13947);
xor UO_568 (O_568,N_14314,N_14430);
nand UO_569 (O_569,N_13841,N_14242);
xnor UO_570 (O_570,N_14552,N_13890);
and UO_571 (O_571,N_14237,N_13851);
and UO_572 (O_572,N_14084,N_14317);
xnor UO_573 (O_573,N_14564,N_13631);
nor UO_574 (O_574,N_14897,N_13621);
nor UO_575 (O_575,N_13552,N_14206);
nor UO_576 (O_576,N_14747,N_14921);
xnor UO_577 (O_577,N_13856,N_14773);
xor UO_578 (O_578,N_13875,N_14140);
nor UO_579 (O_579,N_13535,N_14746);
nand UO_580 (O_580,N_14974,N_14376);
nand UO_581 (O_581,N_14475,N_13923);
xnor UO_582 (O_582,N_14056,N_14920);
or UO_583 (O_583,N_14665,N_14120);
and UO_584 (O_584,N_13711,N_14942);
xor UO_585 (O_585,N_14429,N_13818);
nor UO_586 (O_586,N_13555,N_13674);
or UO_587 (O_587,N_14265,N_14160);
nor UO_588 (O_588,N_13647,N_14557);
or UO_589 (O_589,N_14078,N_14170);
and UO_590 (O_590,N_13848,N_14234);
xor UO_591 (O_591,N_14197,N_14471);
or UO_592 (O_592,N_13805,N_14096);
nand UO_593 (O_593,N_14794,N_14775);
nand UO_594 (O_594,N_13953,N_14268);
and UO_595 (O_595,N_13682,N_13915);
or UO_596 (O_596,N_13917,N_13617);
and UO_597 (O_597,N_13807,N_13644);
or UO_598 (O_598,N_14738,N_14469);
nand UO_599 (O_599,N_14635,N_14353);
or UO_600 (O_600,N_13560,N_14868);
xor UO_601 (O_601,N_13926,N_14764);
and UO_602 (O_602,N_14823,N_14057);
nor UO_603 (O_603,N_14503,N_14792);
and UO_604 (O_604,N_14909,N_14796);
and UO_605 (O_605,N_14153,N_14906);
and UO_606 (O_606,N_14361,N_14810);
and UO_607 (O_607,N_14744,N_14238);
nand UO_608 (O_608,N_13858,N_14990);
nand UO_609 (O_609,N_13809,N_14510);
and UO_610 (O_610,N_14049,N_13761);
or UO_611 (O_611,N_14002,N_14318);
or UO_612 (O_612,N_14569,N_13705);
or UO_613 (O_613,N_13798,N_14070);
and UO_614 (O_614,N_13575,N_13945);
nand UO_615 (O_615,N_14241,N_14541);
and UO_616 (O_616,N_14700,N_13539);
nand UO_617 (O_617,N_13857,N_13952);
nor UO_618 (O_618,N_14012,N_14912);
or UO_619 (O_619,N_13933,N_14752);
and UO_620 (O_620,N_14651,N_14085);
xnor UO_621 (O_621,N_14285,N_14977);
and UO_622 (O_622,N_14051,N_14730);
nor UO_623 (O_623,N_14765,N_14244);
xnor UO_624 (O_624,N_14994,N_13873);
and UO_625 (O_625,N_13855,N_14231);
and UO_626 (O_626,N_13713,N_14481);
xnor UO_627 (O_627,N_14431,N_14228);
nand UO_628 (O_628,N_14166,N_14092);
nand UO_629 (O_629,N_14442,N_14362);
nor UO_630 (O_630,N_14970,N_13880);
nor UO_631 (O_631,N_13607,N_14805);
and UO_632 (O_632,N_14055,N_14933);
nor UO_633 (O_633,N_14058,N_13844);
xor UO_634 (O_634,N_14640,N_14824);
or UO_635 (O_635,N_14780,N_14892);
xor UO_636 (O_636,N_14217,N_14853);
or UO_637 (O_637,N_14157,N_14891);
nand UO_638 (O_638,N_13899,N_13865);
or UO_639 (O_639,N_14462,N_14278);
nor UO_640 (O_640,N_14861,N_14750);
or UO_641 (O_641,N_14118,N_13689);
or UO_642 (O_642,N_14366,N_14117);
nand UO_643 (O_643,N_13639,N_14193);
xnor UO_644 (O_644,N_14992,N_13567);
xnor UO_645 (O_645,N_14668,N_14054);
and UO_646 (O_646,N_14922,N_13520);
nor UO_647 (O_647,N_14359,N_14424);
nand UO_648 (O_648,N_14042,N_14615);
or UO_649 (O_649,N_14513,N_14104);
nand UO_650 (O_650,N_14018,N_14308);
and UO_651 (O_651,N_14877,N_14456);
xor UO_652 (O_652,N_14407,N_14080);
nand UO_653 (O_653,N_14495,N_14043);
nand UO_654 (O_654,N_14666,N_14501);
xor UO_655 (O_655,N_13846,N_13673);
nor UO_656 (O_656,N_13648,N_13526);
nor UO_657 (O_657,N_13603,N_14016);
and UO_658 (O_658,N_14488,N_13655);
nor UO_659 (O_659,N_14871,N_14768);
xnor UO_660 (O_660,N_14930,N_13845);
or UO_661 (O_661,N_14264,N_14248);
and UO_662 (O_662,N_14535,N_14679);
and UO_663 (O_663,N_14363,N_14685);
nand UO_664 (O_664,N_13646,N_14879);
or UO_665 (O_665,N_14371,N_14493);
or UO_666 (O_666,N_13533,N_14189);
nand UO_667 (O_667,N_14779,N_14802);
nand UO_668 (O_668,N_14034,N_14398);
and UO_669 (O_669,N_13686,N_14928);
nand UO_670 (O_670,N_14144,N_14984);
nand UO_671 (O_671,N_14223,N_13800);
nand UO_672 (O_672,N_14337,N_14052);
xor UO_673 (O_673,N_13522,N_14677);
or UO_674 (O_674,N_13726,N_14155);
nor UO_675 (O_675,N_14222,N_13586);
or UO_676 (O_676,N_14473,N_14717);
and UO_677 (O_677,N_14013,N_13671);
or UO_678 (O_678,N_14453,N_14799);
or UO_679 (O_679,N_14642,N_14221);
and UO_680 (O_680,N_14749,N_13840);
nor UO_681 (O_681,N_13553,N_14346);
nor UO_682 (O_682,N_14020,N_14393);
xor UO_683 (O_683,N_14496,N_13735);
or UO_684 (O_684,N_14103,N_14204);
and UO_685 (O_685,N_14297,N_14639);
xnor UO_686 (O_686,N_14329,N_13920);
nand UO_687 (O_687,N_13986,N_13722);
xnor UO_688 (O_688,N_13958,N_13954);
nand UO_689 (O_689,N_13833,N_14616);
nand UO_690 (O_690,N_13669,N_14663);
or UO_691 (O_691,N_13740,N_13859);
nand UO_692 (O_692,N_14519,N_13897);
nor UO_693 (O_693,N_14520,N_13712);
or UO_694 (O_694,N_14982,N_14106);
nand UO_695 (O_695,N_14878,N_14751);
nand UO_696 (O_696,N_14561,N_14408);
nand UO_697 (O_697,N_13799,N_13780);
and UO_698 (O_698,N_14452,N_14649);
or UO_699 (O_699,N_14682,N_13500);
nor UO_700 (O_700,N_14440,N_14619);
or UO_701 (O_701,N_13885,N_14734);
xor UO_702 (O_702,N_13510,N_14007);
or UO_703 (O_703,N_13640,N_14526);
xor UO_704 (O_704,N_13988,N_14575);
and UO_705 (O_705,N_14438,N_14924);
xor UO_706 (O_706,N_14330,N_13623);
nor UO_707 (O_707,N_14852,N_13540);
and UO_708 (O_708,N_14524,N_14681);
nand UO_709 (O_709,N_14415,N_13636);
nand UO_710 (O_710,N_14950,N_14486);
or UO_711 (O_711,N_14958,N_13943);
or UO_712 (O_712,N_14908,N_14418);
and UO_713 (O_713,N_14957,N_14726);
nand UO_714 (O_714,N_14801,N_14037);
and UO_715 (O_715,N_13913,N_14671);
nand UO_716 (O_716,N_14684,N_13662);
and UO_717 (O_717,N_14500,N_14960);
nor UO_718 (O_718,N_14119,N_14617);
xor UO_719 (O_719,N_13793,N_14925);
xor UO_720 (O_720,N_13775,N_13997);
nand UO_721 (O_721,N_14454,N_14038);
nor UO_722 (O_722,N_14661,N_14464);
xnor UO_723 (O_723,N_13871,N_14082);
nor UO_724 (O_724,N_14164,N_13896);
nor UO_725 (O_725,N_14414,N_14652);
nand UO_726 (O_726,N_14954,N_14115);
nand UO_727 (O_727,N_14882,N_14372);
xor UO_728 (O_728,N_13955,N_13771);
xor UO_729 (O_729,N_14162,N_14167);
and UO_730 (O_730,N_13946,N_14716);
nand UO_731 (O_731,N_13766,N_14053);
or UO_732 (O_732,N_14662,N_13704);
nor UO_733 (O_733,N_14781,N_14378);
nor UO_734 (O_734,N_13853,N_14509);
nand UO_735 (O_735,N_14245,N_14420);
nand UO_736 (O_736,N_14598,N_14490);
or UO_737 (O_737,N_14271,N_14586);
and UO_738 (O_738,N_14936,N_14066);
xnor UO_739 (O_739,N_14517,N_13850);
or UO_740 (O_740,N_13927,N_14686);
xor UO_741 (O_741,N_14460,N_13772);
or UO_742 (O_742,N_14316,N_13542);
and UO_743 (O_743,N_14873,N_14447);
or UO_744 (O_744,N_13797,N_14190);
or UO_745 (O_745,N_13795,N_14890);
and UO_746 (O_746,N_13629,N_14492);
and UO_747 (O_747,N_14200,N_13968);
and UO_748 (O_748,N_14620,N_14589);
or UO_749 (O_749,N_14210,N_14422);
nor UO_750 (O_750,N_13578,N_14961);
nand UO_751 (O_751,N_14341,N_14585);
or UO_752 (O_752,N_13976,N_13621);
xor UO_753 (O_753,N_14162,N_14984);
nor UO_754 (O_754,N_14121,N_14471);
xor UO_755 (O_755,N_14737,N_14161);
nor UO_756 (O_756,N_13854,N_14814);
xnor UO_757 (O_757,N_13674,N_13965);
nand UO_758 (O_758,N_13718,N_14927);
or UO_759 (O_759,N_13510,N_14525);
or UO_760 (O_760,N_13524,N_14566);
xor UO_761 (O_761,N_14178,N_14706);
nand UO_762 (O_762,N_14636,N_14542);
or UO_763 (O_763,N_14751,N_13690);
and UO_764 (O_764,N_14938,N_14141);
nor UO_765 (O_765,N_14505,N_14730);
nor UO_766 (O_766,N_14684,N_14177);
and UO_767 (O_767,N_14372,N_13976);
nor UO_768 (O_768,N_13771,N_14037);
xor UO_769 (O_769,N_13648,N_14187);
nor UO_770 (O_770,N_14631,N_14157);
xor UO_771 (O_771,N_13653,N_14615);
and UO_772 (O_772,N_14519,N_13526);
nor UO_773 (O_773,N_14197,N_13940);
and UO_774 (O_774,N_14560,N_13991);
nor UO_775 (O_775,N_14967,N_13525);
xnor UO_776 (O_776,N_14425,N_14159);
xor UO_777 (O_777,N_14548,N_13611);
xor UO_778 (O_778,N_14184,N_14233);
nand UO_779 (O_779,N_14127,N_14204);
nand UO_780 (O_780,N_14032,N_14433);
nor UO_781 (O_781,N_13793,N_14020);
nor UO_782 (O_782,N_13759,N_14233);
xnor UO_783 (O_783,N_13923,N_14816);
nand UO_784 (O_784,N_14885,N_14247);
or UO_785 (O_785,N_14502,N_14305);
xor UO_786 (O_786,N_14908,N_14799);
and UO_787 (O_787,N_13854,N_14970);
xnor UO_788 (O_788,N_14420,N_14033);
xor UO_789 (O_789,N_13587,N_14750);
nor UO_790 (O_790,N_14985,N_13700);
nand UO_791 (O_791,N_14452,N_14965);
or UO_792 (O_792,N_14333,N_14549);
or UO_793 (O_793,N_14711,N_14942);
or UO_794 (O_794,N_13824,N_14870);
xnor UO_795 (O_795,N_13983,N_14085);
nand UO_796 (O_796,N_14436,N_13679);
or UO_797 (O_797,N_13869,N_14494);
xor UO_798 (O_798,N_13898,N_14005);
nor UO_799 (O_799,N_13895,N_14249);
nand UO_800 (O_800,N_13983,N_14995);
nor UO_801 (O_801,N_13541,N_14655);
nor UO_802 (O_802,N_14296,N_14212);
and UO_803 (O_803,N_14285,N_14622);
or UO_804 (O_804,N_14825,N_14118);
nor UO_805 (O_805,N_14795,N_13767);
or UO_806 (O_806,N_14625,N_13607);
and UO_807 (O_807,N_13693,N_13864);
nand UO_808 (O_808,N_14011,N_13695);
or UO_809 (O_809,N_14559,N_14064);
nand UO_810 (O_810,N_14453,N_13974);
xnor UO_811 (O_811,N_14403,N_13617);
or UO_812 (O_812,N_13943,N_14991);
and UO_813 (O_813,N_13681,N_14717);
xnor UO_814 (O_814,N_13847,N_14363);
nand UO_815 (O_815,N_14161,N_14574);
xnor UO_816 (O_816,N_13790,N_13709);
and UO_817 (O_817,N_14507,N_14135);
xor UO_818 (O_818,N_14478,N_13530);
or UO_819 (O_819,N_13893,N_13551);
nor UO_820 (O_820,N_13791,N_13989);
and UO_821 (O_821,N_13926,N_14067);
xnor UO_822 (O_822,N_13548,N_14977);
nand UO_823 (O_823,N_14737,N_14698);
and UO_824 (O_824,N_14129,N_14298);
or UO_825 (O_825,N_14345,N_13939);
and UO_826 (O_826,N_14670,N_13782);
and UO_827 (O_827,N_13898,N_14106);
or UO_828 (O_828,N_14578,N_13824);
nand UO_829 (O_829,N_14583,N_14231);
and UO_830 (O_830,N_14177,N_14191);
xor UO_831 (O_831,N_14541,N_14492);
nand UO_832 (O_832,N_13945,N_14867);
nand UO_833 (O_833,N_14967,N_14438);
xor UO_834 (O_834,N_14950,N_13529);
and UO_835 (O_835,N_14756,N_14018);
and UO_836 (O_836,N_13641,N_14448);
nand UO_837 (O_837,N_14246,N_13716);
or UO_838 (O_838,N_14915,N_13530);
nand UO_839 (O_839,N_14978,N_13508);
nand UO_840 (O_840,N_14076,N_14397);
and UO_841 (O_841,N_14469,N_14392);
or UO_842 (O_842,N_13811,N_13605);
xnor UO_843 (O_843,N_13965,N_14823);
and UO_844 (O_844,N_14242,N_13724);
and UO_845 (O_845,N_13513,N_14674);
nand UO_846 (O_846,N_13512,N_13841);
nand UO_847 (O_847,N_14165,N_14450);
xor UO_848 (O_848,N_13691,N_14152);
nand UO_849 (O_849,N_14342,N_14909);
and UO_850 (O_850,N_14720,N_14238);
and UO_851 (O_851,N_14249,N_13802);
or UO_852 (O_852,N_13935,N_14461);
xor UO_853 (O_853,N_14883,N_14175);
or UO_854 (O_854,N_14449,N_14583);
nand UO_855 (O_855,N_13715,N_14608);
xnor UO_856 (O_856,N_14699,N_13554);
and UO_857 (O_857,N_13943,N_14887);
xnor UO_858 (O_858,N_13618,N_14450);
and UO_859 (O_859,N_13847,N_14876);
nand UO_860 (O_860,N_14147,N_13703);
nand UO_861 (O_861,N_14404,N_14412);
nor UO_862 (O_862,N_14094,N_14331);
xnor UO_863 (O_863,N_13858,N_14364);
nor UO_864 (O_864,N_14473,N_14454);
and UO_865 (O_865,N_14704,N_13698);
nand UO_866 (O_866,N_14908,N_14132);
nor UO_867 (O_867,N_14435,N_14487);
xnor UO_868 (O_868,N_13595,N_13603);
or UO_869 (O_869,N_13714,N_14149);
nor UO_870 (O_870,N_14388,N_13838);
xnor UO_871 (O_871,N_14239,N_14535);
and UO_872 (O_872,N_13536,N_14289);
xor UO_873 (O_873,N_13894,N_14661);
nor UO_874 (O_874,N_14869,N_14842);
or UO_875 (O_875,N_14126,N_14826);
or UO_876 (O_876,N_14315,N_14575);
nand UO_877 (O_877,N_13996,N_14016);
nand UO_878 (O_878,N_13763,N_13877);
nand UO_879 (O_879,N_14016,N_14875);
nor UO_880 (O_880,N_13556,N_14871);
nor UO_881 (O_881,N_13949,N_14112);
or UO_882 (O_882,N_13911,N_14127);
and UO_883 (O_883,N_14335,N_13752);
xnor UO_884 (O_884,N_14594,N_14440);
xor UO_885 (O_885,N_14446,N_14933);
xor UO_886 (O_886,N_13686,N_13625);
xor UO_887 (O_887,N_13599,N_13588);
xor UO_888 (O_888,N_13829,N_13517);
nand UO_889 (O_889,N_14493,N_14248);
and UO_890 (O_890,N_14692,N_14406);
nand UO_891 (O_891,N_14815,N_14124);
nand UO_892 (O_892,N_14656,N_14878);
nor UO_893 (O_893,N_13969,N_13735);
xor UO_894 (O_894,N_13646,N_14551);
and UO_895 (O_895,N_14978,N_14812);
nand UO_896 (O_896,N_13716,N_14543);
nor UO_897 (O_897,N_13685,N_14329);
or UO_898 (O_898,N_14146,N_13954);
and UO_899 (O_899,N_14044,N_13813);
nor UO_900 (O_900,N_14308,N_13816);
nand UO_901 (O_901,N_14302,N_14752);
or UO_902 (O_902,N_14490,N_13936);
or UO_903 (O_903,N_13688,N_14542);
nor UO_904 (O_904,N_14225,N_14854);
or UO_905 (O_905,N_13689,N_13712);
and UO_906 (O_906,N_13863,N_14956);
and UO_907 (O_907,N_14601,N_14696);
xor UO_908 (O_908,N_14971,N_13930);
nand UO_909 (O_909,N_13699,N_14872);
xnor UO_910 (O_910,N_13858,N_13790);
nand UO_911 (O_911,N_13651,N_14198);
nor UO_912 (O_912,N_14314,N_14709);
and UO_913 (O_913,N_14085,N_13621);
xor UO_914 (O_914,N_14050,N_14920);
nand UO_915 (O_915,N_13593,N_13840);
xor UO_916 (O_916,N_13856,N_14476);
nor UO_917 (O_917,N_14332,N_14288);
xor UO_918 (O_918,N_13720,N_14002);
xnor UO_919 (O_919,N_13502,N_14485);
and UO_920 (O_920,N_14137,N_14565);
and UO_921 (O_921,N_14308,N_13708);
nor UO_922 (O_922,N_14559,N_14025);
nand UO_923 (O_923,N_14332,N_14840);
nor UO_924 (O_924,N_13580,N_13765);
or UO_925 (O_925,N_14203,N_13570);
nand UO_926 (O_926,N_14924,N_14444);
xor UO_927 (O_927,N_14925,N_14547);
and UO_928 (O_928,N_13745,N_14202);
and UO_929 (O_929,N_13862,N_13600);
and UO_930 (O_930,N_14493,N_14217);
nand UO_931 (O_931,N_14151,N_13843);
nand UO_932 (O_932,N_14383,N_13698);
or UO_933 (O_933,N_13526,N_13727);
nor UO_934 (O_934,N_14278,N_14001);
nor UO_935 (O_935,N_14291,N_14729);
nand UO_936 (O_936,N_14488,N_13578);
and UO_937 (O_937,N_13523,N_14350);
and UO_938 (O_938,N_14839,N_14768);
nand UO_939 (O_939,N_14886,N_14856);
nand UO_940 (O_940,N_14407,N_14348);
xor UO_941 (O_941,N_14197,N_14125);
and UO_942 (O_942,N_14211,N_14769);
nand UO_943 (O_943,N_13828,N_14617);
nor UO_944 (O_944,N_14482,N_13853);
nor UO_945 (O_945,N_14543,N_14150);
nor UO_946 (O_946,N_14309,N_14325);
nor UO_947 (O_947,N_13687,N_13793);
or UO_948 (O_948,N_14723,N_14626);
xnor UO_949 (O_949,N_14377,N_14876);
nand UO_950 (O_950,N_13785,N_14681);
or UO_951 (O_951,N_13961,N_13715);
nand UO_952 (O_952,N_14178,N_14388);
nor UO_953 (O_953,N_14854,N_14335);
xnor UO_954 (O_954,N_14005,N_13723);
nand UO_955 (O_955,N_13707,N_14067);
nand UO_956 (O_956,N_14701,N_14200);
and UO_957 (O_957,N_14308,N_13857);
and UO_958 (O_958,N_13791,N_14101);
xnor UO_959 (O_959,N_14591,N_14084);
nor UO_960 (O_960,N_14234,N_14426);
xor UO_961 (O_961,N_14349,N_14256);
or UO_962 (O_962,N_14347,N_14559);
nand UO_963 (O_963,N_13881,N_13822);
nor UO_964 (O_964,N_14890,N_14190);
xnor UO_965 (O_965,N_14338,N_14842);
nor UO_966 (O_966,N_14013,N_13576);
xor UO_967 (O_967,N_13589,N_14027);
nor UO_968 (O_968,N_13520,N_14059);
nor UO_969 (O_969,N_14974,N_14719);
nand UO_970 (O_970,N_14972,N_14664);
nor UO_971 (O_971,N_13717,N_13802);
or UO_972 (O_972,N_14552,N_14615);
nor UO_973 (O_973,N_13924,N_14638);
nand UO_974 (O_974,N_13532,N_14575);
nor UO_975 (O_975,N_14288,N_14368);
nand UO_976 (O_976,N_13781,N_13615);
nand UO_977 (O_977,N_13822,N_14804);
xnor UO_978 (O_978,N_13826,N_14585);
nor UO_979 (O_979,N_14703,N_13584);
and UO_980 (O_980,N_13998,N_13558);
or UO_981 (O_981,N_14228,N_14610);
xor UO_982 (O_982,N_13987,N_14312);
xor UO_983 (O_983,N_14747,N_14888);
nor UO_984 (O_984,N_14335,N_13508);
nand UO_985 (O_985,N_14782,N_14801);
nand UO_986 (O_986,N_13898,N_14670);
and UO_987 (O_987,N_14938,N_14787);
and UO_988 (O_988,N_13829,N_13931);
nor UO_989 (O_989,N_14465,N_14214);
and UO_990 (O_990,N_14218,N_14453);
nand UO_991 (O_991,N_14087,N_13690);
nand UO_992 (O_992,N_14822,N_14109);
nand UO_993 (O_993,N_14125,N_13583);
nor UO_994 (O_994,N_14346,N_13764);
or UO_995 (O_995,N_14159,N_14980);
or UO_996 (O_996,N_13835,N_14248);
and UO_997 (O_997,N_14913,N_14389);
and UO_998 (O_998,N_13566,N_14338);
nand UO_999 (O_999,N_14428,N_13570);
nor UO_1000 (O_1000,N_13689,N_13720);
or UO_1001 (O_1001,N_14823,N_14320);
xnor UO_1002 (O_1002,N_14282,N_13888);
xor UO_1003 (O_1003,N_14196,N_14401);
xnor UO_1004 (O_1004,N_14301,N_13699);
xnor UO_1005 (O_1005,N_14433,N_14286);
xnor UO_1006 (O_1006,N_13803,N_14768);
and UO_1007 (O_1007,N_14821,N_13536);
or UO_1008 (O_1008,N_13604,N_13821);
and UO_1009 (O_1009,N_13682,N_14722);
nand UO_1010 (O_1010,N_14828,N_14224);
xnor UO_1011 (O_1011,N_13985,N_14219);
xor UO_1012 (O_1012,N_13768,N_13857);
and UO_1013 (O_1013,N_14131,N_14327);
or UO_1014 (O_1014,N_13540,N_14326);
and UO_1015 (O_1015,N_14663,N_13722);
xnor UO_1016 (O_1016,N_13727,N_14319);
xor UO_1017 (O_1017,N_13602,N_14365);
nor UO_1018 (O_1018,N_14218,N_13712);
and UO_1019 (O_1019,N_14539,N_14582);
nor UO_1020 (O_1020,N_14016,N_13521);
or UO_1021 (O_1021,N_14565,N_14423);
xnor UO_1022 (O_1022,N_14173,N_13714);
xor UO_1023 (O_1023,N_13853,N_14843);
nand UO_1024 (O_1024,N_14934,N_13757);
nor UO_1025 (O_1025,N_14056,N_14089);
xor UO_1026 (O_1026,N_14700,N_13559);
xor UO_1027 (O_1027,N_14820,N_14071);
nand UO_1028 (O_1028,N_13763,N_14307);
nand UO_1029 (O_1029,N_14387,N_14092);
nor UO_1030 (O_1030,N_13806,N_14785);
and UO_1031 (O_1031,N_14440,N_13655);
xnor UO_1032 (O_1032,N_13809,N_14948);
or UO_1033 (O_1033,N_13540,N_13544);
xor UO_1034 (O_1034,N_14465,N_14750);
nor UO_1035 (O_1035,N_14311,N_14598);
and UO_1036 (O_1036,N_14453,N_14562);
or UO_1037 (O_1037,N_13842,N_13882);
xnor UO_1038 (O_1038,N_14326,N_14383);
and UO_1039 (O_1039,N_13883,N_13905);
or UO_1040 (O_1040,N_13582,N_13729);
nor UO_1041 (O_1041,N_13744,N_13624);
xor UO_1042 (O_1042,N_13779,N_14556);
and UO_1043 (O_1043,N_13795,N_14346);
nor UO_1044 (O_1044,N_14199,N_14195);
and UO_1045 (O_1045,N_14911,N_13903);
and UO_1046 (O_1046,N_14806,N_14499);
and UO_1047 (O_1047,N_14962,N_14026);
nand UO_1048 (O_1048,N_13859,N_14930);
nand UO_1049 (O_1049,N_13880,N_14809);
nand UO_1050 (O_1050,N_14399,N_13607);
and UO_1051 (O_1051,N_13677,N_13509);
or UO_1052 (O_1052,N_14339,N_14203);
and UO_1053 (O_1053,N_14389,N_14280);
nor UO_1054 (O_1054,N_14316,N_14579);
nand UO_1055 (O_1055,N_14644,N_13663);
xnor UO_1056 (O_1056,N_14972,N_14556);
or UO_1057 (O_1057,N_13952,N_14499);
or UO_1058 (O_1058,N_14497,N_14194);
and UO_1059 (O_1059,N_14595,N_14588);
or UO_1060 (O_1060,N_14560,N_13568);
and UO_1061 (O_1061,N_13671,N_14374);
nor UO_1062 (O_1062,N_14270,N_13728);
nor UO_1063 (O_1063,N_14334,N_14738);
xnor UO_1064 (O_1064,N_13539,N_14757);
nor UO_1065 (O_1065,N_13928,N_13575);
nand UO_1066 (O_1066,N_14368,N_14303);
xnor UO_1067 (O_1067,N_13972,N_14415);
nor UO_1068 (O_1068,N_14691,N_13664);
nor UO_1069 (O_1069,N_13917,N_14918);
or UO_1070 (O_1070,N_13932,N_13625);
xnor UO_1071 (O_1071,N_14742,N_13995);
nor UO_1072 (O_1072,N_14058,N_13833);
xor UO_1073 (O_1073,N_13905,N_13899);
nor UO_1074 (O_1074,N_14968,N_14658);
or UO_1075 (O_1075,N_14009,N_14398);
xnor UO_1076 (O_1076,N_14082,N_14167);
or UO_1077 (O_1077,N_13558,N_14186);
or UO_1078 (O_1078,N_14016,N_14381);
nand UO_1079 (O_1079,N_14060,N_14541);
or UO_1080 (O_1080,N_13704,N_14475);
and UO_1081 (O_1081,N_14977,N_14366);
xor UO_1082 (O_1082,N_14686,N_14550);
nand UO_1083 (O_1083,N_13500,N_14125);
and UO_1084 (O_1084,N_14262,N_14224);
xor UO_1085 (O_1085,N_14555,N_13592);
and UO_1086 (O_1086,N_13548,N_13573);
and UO_1087 (O_1087,N_14834,N_14255);
and UO_1088 (O_1088,N_13960,N_14979);
or UO_1089 (O_1089,N_14018,N_14727);
and UO_1090 (O_1090,N_14255,N_14618);
or UO_1091 (O_1091,N_14067,N_14005);
or UO_1092 (O_1092,N_13539,N_14753);
or UO_1093 (O_1093,N_14615,N_14644);
and UO_1094 (O_1094,N_14169,N_13685);
and UO_1095 (O_1095,N_14260,N_14006);
and UO_1096 (O_1096,N_14651,N_13809);
or UO_1097 (O_1097,N_14317,N_14957);
xnor UO_1098 (O_1098,N_13865,N_13988);
or UO_1099 (O_1099,N_13852,N_14529);
xnor UO_1100 (O_1100,N_14333,N_14094);
xor UO_1101 (O_1101,N_13816,N_14568);
nand UO_1102 (O_1102,N_14426,N_14461);
or UO_1103 (O_1103,N_13577,N_13613);
xor UO_1104 (O_1104,N_13511,N_14604);
nand UO_1105 (O_1105,N_13661,N_14527);
nor UO_1106 (O_1106,N_14283,N_14015);
xnor UO_1107 (O_1107,N_14101,N_14618);
and UO_1108 (O_1108,N_14829,N_14307);
or UO_1109 (O_1109,N_14228,N_14105);
or UO_1110 (O_1110,N_14015,N_13926);
xnor UO_1111 (O_1111,N_14972,N_14291);
nor UO_1112 (O_1112,N_14936,N_14202);
and UO_1113 (O_1113,N_13892,N_14053);
or UO_1114 (O_1114,N_14660,N_14399);
xnor UO_1115 (O_1115,N_14909,N_14205);
and UO_1116 (O_1116,N_14292,N_14501);
nor UO_1117 (O_1117,N_14180,N_14991);
nand UO_1118 (O_1118,N_14359,N_13688);
or UO_1119 (O_1119,N_13869,N_14747);
nor UO_1120 (O_1120,N_13837,N_14521);
and UO_1121 (O_1121,N_14061,N_14650);
nor UO_1122 (O_1122,N_14389,N_14151);
xnor UO_1123 (O_1123,N_14356,N_14528);
nand UO_1124 (O_1124,N_14026,N_13874);
or UO_1125 (O_1125,N_13785,N_13560);
or UO_1126 (O_1126,N_13585,N_14444);
xor UO_1127 (O_1127,N_14337,N_13884);
or UO_1128 (O_1128,N_13900,N_13573);
nand UO_1129 (O_1129,N_14033,N_13644);
and UO_1130 (O_1130,N_14354,N_13716);
or UO_1131 (O_1131,N_14746,N_14842);
nand UO_1132 (O_1132,N_14888,N_14696);
or UO_1133 (O_1133,N_14722,N_14100);
nor UO_1134 (O_1134,N_13652,N_14335);
and UO_1135 (O_1135,N_14527,N_13631);
xnor UO_1136 (O_1136,N_13547,N_14767);
nand UO_1137 (O_1137,N_14246,N_13807);
and UO_1138 (O_1138,N_14925,N_14596);
nor UO_1139 (O_1139,N_14476,N_14054);
and UO_1140 (O_1140,N_14551,N_14697);
nand UO_1141 (O_1141,N_14837,N_14745);
nor UO_1142 (O_1142,N_14160,N_14138);
nor UO_1143 (O_1143,N_14355,N_13600);
xnor UO_1144 (O_1144,N_13537,N_14346);
and UO_1145 (O_1145,N_14272,N_14353);
or UO_1146 (O_1146,N_13873,N_13811);
and UO_1147 (O_1147,N_14426,N_14154);
and UO_1148 (O_1148,N_14662,N_14363);
and UO_1149 (O_1149,N_14264,N_13684);
or UO_1150 (O_1150,N_14843,N_13786);
and UO_1151 (O_1151,N_14945,N_14920);
and UO_1152 (O_1152,N_14653,N_13638);
or UO_1153 (O_1153,N_14290,N_14786);
or UO_1154 (O_1154,N_14709,N_14235);
nor UO_1155 (O_1155,N_14790,N_13835);
or UO_1156 (O_1156,N_13805,N_13687);
nand UO_1157 (O_1157,N_14389,N_13756);
nand UO_1158 (O_1158,N_14666,N_14976);
xor UO_1159 (O_1159,N_14212,N_13578);
xor UO_1160 (O_1160,N_14804,N_14280);
and UO_1161 (O_1161,N_14342,N_14594);
xor UO_1162 (O_1162,N_13531,N_13761);
or UO_1163 (O_1163,N_14736,N_14312);
nand UO_1164 (O_1164,N_14442,N_14193);
or UO_1165 (O_1165,N_14105,N_14132);
or UO_1166 (O_1166,N_14689,N_13690);
or UO_1167 (O_1167,N_13882,N_14682);
nor UO_1168 (O_1168,N_13720,N_14745);
nor UO_1169 (O_1169,N_13849,N_13951);
nand UO_1170 (O_1170,N_14577,N_13885);
nand UO_1171 (O_1171,N_14780,N_13906);
xnor UO_1172 (O_1172,N_13999,N_14472);
xor UO_1173 (O_1173,N_14608,N_14091);
xor UO_1174 (O_1174,N_13512,N_14435);
nand UO_1175 (O_1175,N_13797,N_14834);
xnor UO_1176 (O_1176,N_13867,N_13965);
nor UO_1177 (O_1177,N_14738,N_14190);
or UO_1178 (O_1178,N_13546,N_14538);
and UO_1179 (O_1179,N_14096,N_14774);
nor UO_1180 (O_1180,N_13570,N_13732);
and UO_1181 (O_1181,N_13600,N_14169);
or UO_1182 (O_1182,N_14207,N_13684);
or UO_1183 (O_1183,N_14761,N_13994);
nor UO_1184 (O_1184,N_14360,N_14643);
nand UO_1185 (O_1185,N_13640,N_14546);
or UO_1186 (O_1186,N_14060,N_14644);
nor UO_1187 (O_1187,N_13598,N_14905);
nor UO_1188 (O_1188,N_14874,N_13562);
xor UO_1189 (O_1189,N_14811,N_13946);
nand UO_1190 (O_1190,N_14864,N_14383);
nor UO_1191 (O_1191,N_14333,N_14168);
or UO_1192 (O_1192,N_14706,N_14938);
xnor UO_1193 (O_1193,N_14771,N_13892);
nand UO_1194 (O_1194,N_14757,N_13853);
nand UO_1195 (O_1195,N_13864,N_14632);
xnor UO_1196 (O_1196,N_14596,N_14556);
nand UO_1197 (O_1197,N_14696,N_14325);
nand UO_1198 (O_1198,N_14379,N_14098);
xnor UO_1199 (O_1199,N_13772,N_13952);
or UO_1200 (O_1200,N_13589,N_14893);
nand UO_1201 (O_1201,N_14921,N_13736);
and UO_1202 (O_1202,N_14937,N_14518);
or UO_1203 (O_1203,N_14755,N_13793);
nand UO_1204 (O_1204,N_14439,N_14452);
nand UO_1205 (O_1205,N_13670,N_14205);
xnor UO_1206 (O_1206,N_14721,N_14634);
or UO_1207 (O_1207,N_14152,N_14081);
nor UO_1208 (O_1208,N_14921,N_14261);
xnor UO_1209 (O_1209,N_14131,N_13916);
or UO_1210 (O_1210,N_14503,N_14198);
nor UO_1211 (O_1211,N_13588,N_14390);
or UO_1212 (O_1212,N_14944,N_14575);
or UO_1213 (O_1213,N_14637,N_13853);
nand UO_1214 (O_1214,N_14550,N_14459);
xnor UO_1215 (O_1215,N_13604,N_14219);
and UO_1216 (O_1216,N_14938,N_14874);
nor UO_1217 (O_1217,N_13666,N_14240);
or UO_1218 (O_1218,N_13942,N_13529);
nand UO_1219 (O_1219,N_13708,N_14592);
nor UO_1220 (O_1220,N_14870,N_13758);
nor UO_1221 (O_1221,N_13967,N_13798);
xnor UO_1222 (O_1222,N_13846,N_14703);
nand UO_1223 (O_1223,N_14093,N_14834);
nand UO_1224 (O_1224,N_13909,N_13719);
nor UO_1225 (O_1225,N_14495,N_14931);
nor UO_1226 (O_1226,N_14274,N_14079);
or UO_1227 (O_1227,N_13714,N_13892);
nor UO_1228 (O_1228,N_13501,N_14757);
xnor UO_1229 (O_1229,N_14904,N_14886);
nor UO_1230 (O_1230,N_14563,N_13883);
nand UO_1231 (O_1231,N_13978,N_14484);
xnor UO_1232 (O_1232,N_13690,N_14912);
nand UO_1233 (O_1233,N_14791,N_14572);
xor UO_1234 (O_1234,N_14570,N_13828);
nor UO_1235 (O_1235,N_14629,N_13782);
or UO_1236 (O_1236,N_14051,N_14819);
or UO_1237 (O_1237,N_13888,N_13812);
and UO_1238 (O_1238,N_14708,N_13859);
nand UO_1239 (O_1239,N_14163,N_14674);
or UO_1240 (O_1240,N_14793,N_14361);
xnor UO_1241 (O_1241,N_14016,N_14416);
or UO_1242 (O_1242,N_14461,N_13775);
nor UO_1243 (O_1243,N_14840,N_14194);
xor UO_1244 (O_1244,N_14317,N_14431);
nor UO_1245 (O_1245,N_13817,N_14308);
or UO_1246 (O_1246,N_14791,N_14926);
nand UO_1247 (O_1247,N_14538,N_14471);
nand UO_1248 (O_1248,N_14462,N_14953);
xnor UO_1249 (O_1249,N_14839,N_14897);
xnor UO_1250 (O_1250,N_14154,N_14112);
nand UO_1251 (O_1251,N_14313,N_14359);
nand UO_1252 (O_1252,N_14975,N_14123);
xor UO_1253 (O_1253,N_14220,N_13634);
and UO_1254 (O_1254,N_13665,N_13866);
and UO_1255 (O_1255,N_14589,N_13718);
or UO_1256 (O_1256,N_14642,N_13843);
nor UO_1257 (O_1257,N_14125,N_13710);
or UO_1258 (O_1258,N_14592,N_14195);
nor UO_1259 (O_1259,N_13825,N_13606);
xor UO_1260 (O_1260,N_13693,N_13895);
nand UO_1261 (O_1261,N_13709,N_14144);
and UO_1262 (O_1262,N_13951,N_14653);
or UO_1263 (O_1263,N_14464,N_14870);
xnor UO_1264 (O_1264,N_14914,N_13630);
nor UO_1265 (O_1265,N_14808,N_13651);
xor UO_1266 (O_1266,N_13786,N_13547);
xnor UO_1267 (O_1267,N_13929,N_13593);
or UO_1268 (O_1268,N_14874,N_13572);
xnor UO_1269 (O_1269,N_14485,N_14075);
nor UO_1270 (O_1270,N_13839,N_13943);
nand UO_1271 (O_1271,N_13784,N_14441);
or UO_1272 (O_1272,N_14018,N_13805);
or UO_1273 (O_1273,N_14942,N_14015);
nor UO_1274 (O_1274,N_14206,N_14051);
xnor UO_1275 (O_1275,N_13631,N_14569);
and UO_1276 (O_1276,N_14786,N_14824);
nor UO_1277 (O_1277,N_14368,N_14668);
nor UO_1278 (O_1278,N_14251,N_14160);
or UO_1279 (O_1279,N_14703,N_14331);
xnor UO_1280 (O_1280,N_14829,N_14845);
and UO_1281 (O_1281,N_14799,N_13704);
xor UO_1282 (O_1282,N_14266,N_14465);
and UO_1283 (O_1283,N_13513,N_14768);
nor UO_1284 (O_1284,N_14853,N_13539);
nand UO_1285 (O_1285,N_14944,N_14203);
and UO_1286 (O_1286,N_14442,N_14197);
nor UO_1287 (O_1287,N_14733,N_13957);
xnor UO_1288 (O_1288,N_13937,N_14531);
nor UO_1289 (O_1289,N_14140,N_14687);
nand UO_1290 (O_1290,N_14293,N_14930);
nor UO_1291 (O_1291,N_14545,N_13554);
nand UO_1292 (O_1292,N_14851,N_13584);
nand UO_1293 (O_1293,N_13939,N_13905);
nor UO_1294 (O_1294,N_13854,N_14586);
xnor UO_1295 (O_1295,N_14297,N_13795);
xor UO_1296 (O_1296,N_14426,N_13547);
nor UO_1297 (O_1297,N_13775,N_14780);
nor UO_1298 (O_1298,N_14004,N_13761);
nand UO_1299 (O_1299,N_14842,N_13556);
nor UO_1300 (O_1300,N_14071,N_14994);
xor UO_1301 (O_1301,N_14236,N_13583);
and UO_1302 (O_1302,N_14167,N_14030);
or UO_1303 (O_1303,N_14571,N_13888);
or UO_1304 (O_1304,N_14821,N_13886);
and UO_1305 (O_1305,N_14757,N_13650);
nand UO_1306 (O_1306,N_14977,N_14131);
xor UO_1307 (O_1307,N_14259,N_13889);
or UO_1308 (O_1308,N_14540,N_14297);
and UO_1309 (O_1309,N_13820,N_14413);
and UO_1310 (O_1310,N_14199,N_13813);
nand UO_1311 (O_1311,N_14750,N_14843);
or UO_1312 (O_1312,N_13941,N_14594);
or UO_1313 (O_1313,N_14164,N_14784);
nor UO_1314 (O_1314,N_14374,N_14982);
nand UO_1315 (O_1315,N_13884,N_13714);
nor UO_1316 (O_1316,N_13546,N_14514);
nor UO_1317 (O_1317,N_14252,N_13983);
nor UO_1318 (O_1318,N_14022,N_14228);
nor UO_1319 (O_1319,N_14082,N_13511);
and UO_1320 (O_1320,N_13821,N_13687);
nand UO_1321 (O_1321,N_13666,N_13941);
or UO_1322 (O_1322,N_13831,N_14353);
nor UO_1323 (O_1323,N_14878,N_14574);
or UO_1324 (O_1324,N_13969,N_13593);
nor UO_1325 (O_1325,N_13935,N_13595);
or UO_1326 (O_1326,N_14280,N_14189);
nand UO_1327 (O_1327,N_14204,N_13813);
xor UO_1328 (O_1328,N_13878,N_14377);
and UO_1329 (O_1329,N_14107,N_14631);
or UO_1330 (O_1330,N_14498,N_14280);
and UO_1331 (O_1331,N_13706,N_13940);
xnor UO_1332 (O_1332,N_13965,N_14197);
xnor UO_1333 (O_1333,N_14895,N_14789);
nand UO_1334 (O_1334,N_14036,N_14071);
nor UO_1335 (O_1335,N_14254,N_13740);
xnor UO_1336 (O_1336,N_14884,N_14319);
or UO_1337 (O_1337,N_14036,N_14709);
nand UO_1338 (O_1338,N_14169,N_13975);
xnor UO_1339 (O_1339,N_13782,N_14095);
and UO_1340 (O_1340,N_14796,N_14246);
xnor UO_1341 (O_1341,N_14787,N_13972);
or UO_1342 (O_1342,N_14642,N_14808);
or UO_1343 (O_1343,N_14968,N_14905);
nand UO_1344 (O_1344,N_13982,N_14484);
nor UO_1345 (O_1345,N_14107,N_14389);
and UO_1346 (O_1346,N_13818,N_14456);
nand UO_1347 (O_1347,N_14589,N_13883);
nand UO_1348 (O_1348,N_14408,N_14407);
nor UO_1349 (O_1349,N_13930,N_14581);
xor UO_1350 (O_1350,N_14694,N_13925);
nor UO_1351 (O_1351,N_13552,N_14634);
nor UO_1352 (O_1352,N_13620,N_14223);
and UO_1353 (O_1353,N_13841,N_13922);
xnor UO_1354 (O_1354,N_14219,N_13679);
and UO_1355 (O_1355,N_14259,N_14193);
xnor UO_1356 (O_1356,N_14552,N_14234);
nand UO_1357 (O_1357,N_14701,N_13703);
nor UO_1358 (O_1358,N_14594,N_14697);
nor UO_1359 (O_1359,N_13698,N_13872);
nand UO_1360 (O_1360,N_14449,N_13909);
xnor UO_1361 (O_1361,N_14238,N_14613);
and UO_1362 (O_1362,N_13933,N_13936);
nand UO_1363 (O_1363,N_13950,N_14495);
nor UO_1364 (O_1364,N_14807,N_13854);
or UO_1365 (O_1365,N_13607,N_14769);
and UO_1366 (O_1366,N_14213,N_14429);
and UO_1367 (O_1367,N_14903,N_14506);
nand UO_1368 (O_1368,N_14162,N_14755);
and UO_1369 (O_1369,N_14105,N_14748);
xor UO_1370 (O_1370,N_13956,N_14322);
or UO_1371 (O_1371,N_14088,N_13736);
nor UO_1372 (O_1372,N_14666,N_14916);
and UO_1373 (O_1373,N_13706,N_14414);
nand UO_1374 (O_1374,N_14207,N_14264);
xor UO_1375 (O_1375,N_13827,N_13717);
and UO_1376 (O_1376,N_14662,N_14232);
nand UO_1377 (O_1377,N_14091,N_13711);
nor UO_1378 (O_1378,N_13592,N_14808);
nand UO_1379 (O_1379,N_14560,N_14201);
nor UO_1380 (O_1380,N_13835,N_14750);
nor UO_1381 (O_1381,N_13734,N_14456);
and UO_1382 (O_1382,N_13757,N_14498);
xor UO_1383 (O_1383,N_14149,N_13654);
nand UO_1384 (O_1384,N_14747,N_14478);
nand UO_1385 (O_1385,N_14078,N_13752);
or UO_1386 (O_1386,N_14171,N_13654);
and UO_1387 (O_1387,N_14918,N_14180);
nor UO_1388 (O_1388,N_14698,N_13678);
xor UO_1389 (O_1389,N_14867,N_14872);
nand UO_1390 (O_1390,N_13972,N_13690);
nor UO_1391 (O_1391,N_14959,N_13969);
nor UO_1392 (O_1392,N_13542,N_14697);
xor UO_1393 (O_1393,N_14542,N_14928);
and UO_1394 (O_1394,N_13986,N_13644);
xor UO_1395 (O_1395,N_14856,N_14153);
nor UO_1396 (O_1396,N_13908,N_14276);
xor UO_1397 (O_1397,N_14697,N_13787);
nor UO_1398 (O_1398,N_14274,N_14289);
nand UO_1399 (O_1399,N_14821,N_13518);
nor UO_1400 (O_1400,N_13931,N_14345);
xnor UO_1401 (O_1401,N_14424,N_14085);
nor UO_1402 (O_1402,N_14457,N_13657);
or UO_1403 (O_1403,N_13972,N_14303);
or UO_1404 (O_1404,N_13728,N_14137);
and UO_1405 (O_1405,N_13738,N_14942);
xnor UO_1406 (O_1406,N_13919,N_14178);
and UO_1407 (O_1407,N_14263,N_14476);
and UO_1408 (O_1408,N_14158,N_13888);
or UO_1409 (O_1409,N_13715,N_14279);
or UO_1410 (O_1410,N_14631,N_14626);
and UO_1411 (O_1411,N_14584,N_14058);
or UO_1412 (O_1412,N_13850,N_14155);
and UO_1413 (O_1413,N_14146,N_13817);
or UO_1414 (O_1414,N_14988,N_14526);
nor UO_1415 (O_1415,N_14173,N_13804);
xor UO_1416 (O_1416,N_14746,N_13510);
and UO_1417 (O_1417,N_14588,N_14069);
or UO_1418 (O_1418,N_14295,N_14843);
and UO_1419 (O_1419,N_14402,N_13701);
nand UO_1420 (O_1420,N_14384,N_13543);
nand UO_1421 (O_1421,N_14440,N_14707);
nand UO_1422 (O_1422,N_13506,N_14484);
and UO_1423 (O_1423,N_14703,N_14661);
nand UO_1424 (O_1424,N_14392,N_14719);
and UO_1425 (O_1425,N_14363,N_13590);
and UO_1426 (O_1426,N_13729,N_14991);
nor UO_1427 (O_1427,N_14210,N_14153);
nand UO_1428 (O_1428,N_14014,N_14008);
xnor UO_1429 (O_1429,N_14581,N_13886);
and UO_1430 (O_1430,N_14732,N_14655);
or UO_1431 (O_1431,N_13649,N_14510);
xnor UO_1432 (O_1432,N_14236,N_13813);
and UO_1433 (O_1433,N_14771,N_14662);
and UO_1434 (O_1434,N_14990,N_14118);
xor UO_1435 (O_1435,N_14645,N_14076);
nor UO_1436 (O_1436,N_14320,N_14854);
xnor UO_1437 (O_1437,N_14742,N_14202);
and UO_1438 (O_1438,N_14677,N_14859);
and UO_1439 (O_1439,N_14908,N_13943);
and UO_1440 (O_1440,N_14311,N_14326);
nand UO_1441 (O_1441,N_13992,N_13630);
nor UO_1442 (O_1442,N_13735,N_14565);
or UO_1443 (O_1443,N_14731,N_14627);
nor UO_1444 (O_1444,N_13761,N_13833);
xor UO_1445 (O_1445,N_14141,N_14304);
nand UO_1446 (O_1446,N_13519,N_13903);
or UO_1447 (O_1447,N_14898,N_14834);
xor UO_1448 (O_1448,N_14210,N_13807);
xor UO_1449 (O_1449,N_13929,N_14836);
nand UO_1450 (O_1450,N_14865,N_14550);
and UO_1451 (O_1451,N_14056,N_14217);
or UO_1452 (O_1452,N_14108,N_14319);
nand UO_1453 (O_1453,N_14749,N_14200);
nand UO_1454 (O_1454,N_14698,N_14270);
xnor UO_1455 (O_1455,N_14745,N_14540);
or UO_1456 (O_1456,N_14876,N_14836);
nor UO_1457 (O_1457,N_14898,N_13828);
nand UO_1458 (O_1458,N_13848,N_14552);
nand UO_1459 (O_1459,N_14553,N_14675);
nor UO_1460 (O_1460,N_13832,N_13837);
nor UO_1461 (O_1461,N_13977,N_14915);
or UO_1462 (O_1462,N_14618,N_14405);
nand UO_1463 (O_1463,N_14056,N_14740);
nand UO_1464 (O_1464,N_14750,N_13880);
nand UO_1465 (O_1465,N_14734,N_14731);
xnor UO_1466 (O_1466,N_14977,N_14650);
or UO_1467 (O_1467,N_14038,N_13847);
and UO_1468 (O_1468,N_14621,N_14908);
or UO_1469 (O_1469,N_14831,N_13676);
or UO_1470 (O_1470,N_14863,N_14512);
nor UO_1471 (O_1471,N_13952,N_14964);
nor UO_1472 (O_1472,N_13543,N_13981);
nand UO_1473 (O_1473,N_14144,N_13941);
nor UO_1474 (O_1474,N_13582,N_14283);
xor UO_1475 (O_1475,N_14931,N_14655);
nor UO_1476 (O_1476,N_14655,N_14386);
and UO_1477 (O_1477,N_14611,N_13645);
and UO_1478 (O_1478,N_13909,N_13774);
or UO_1479 (O_1479,N_14483,N_14501);
xor UO_1480 (O_1480,N_14889,N_14354);
xor UO_1481 (O_1481,N_13581,N_14383);
nand UO_1482 (O_1482,N_14043,N_14460);
and UO_1483 (O_1483,N_14157,N_14476);
nor UO_1484 (O_1484,N_14125,N_13751);
nor UO_1485 (O_1485,N_14690,N_13537);
nand UO_1486 (O_1486,N_14929,N_14265);
nand UO_1487 (O_1487,N_14344,N_14165);
nor UO_1488 (O_1488,N_14669,N_13642);
nand UO_1489 (O_1489,N_13502,N_14790);
xnor UO_1490 (O_1490,N_14122,N_14490);
or UO_1491 (O_1491,N_13505,N_13869);
and UO_1492 (O_1492,N_13817,N_14444);
and UO_1493 (O_1493,N_14634,N_14730);
nand UO_1494 (O_1494,N_14957,N_14729);
nand UO_1495 (O_1495,N_13549,N_14269);
xnor UO_1496 (O_1496,N_14611,N_14012);
or UO_1497 (O_1497,N_14850,N_14846);
nand UO_1498 (O_1498,N_14296,N_14581);
and UO_1499 (O_1499,N_13718,N_14685);
nand UO_1500 (O_1500,N_14397,N_14861);
or UO_1501 (O_1501,N_14587,N_14961);
and UO_1502 (O_1502,N_14059,N_13723);
nand UO_1503 (O_1503,N_14114,N_13701);
nor UO_1504 (O_1504,N_14816,N_13581);
and UO_1505 (O_1505,N_14736,N_13815);
and UO_1506 (O_1506,N_14275,N_14385);
and UO_1507 (O_1507,N_14930,N_14546);
xnor UO_1508 (O_1508,N_14910,N_13773);
nor UO_1509 (O_1509,N_14181,N_14375);
nor UO_1510 (O_1510,N_14912,N_14910);
nand UO_1511 (O_1511,N_14836,N_14067);
and UO_1512 (O_1512,N_14693,N_14625);
xor UO_1513 (O_1513,N_14326,N_13918);
or UO_1514 (O_1514,N_13730,N_13965);
nor UO_1515 (O_1515,N_14230,N_13910);
and UO_1516 (O_1516,N_14463,N_14937);
and UO_1517 (O_1517,N_13539,N_13577);
or UO_1518 (O_1518,N_14461,N_13676);
or UO_1519 (O_1519,N_14885,N_13618);
nor UO_1520 (O_1520,N_14524,N_14023);
xnor UO_1521 (O_1521,N_14326,N_14732);
and UO_1522 (O_1522,N_14729,N_14726);
xor UO_1523 (O_1523,N_13551,N_14446);
xor UO_1524 (O_1524,N_14710,N_14731);
nor UO_1525 (O_1525,N_14847,N_14701);
nand UO_1526 (O_1526,N_14128,N_14731);
nand UO_1527 (O_1527,N_14410,N_14843);
and UO_1528 (O_1528,N_13942,N_14172);
nand UO_1529 (O_1529,N_14290,N_13981);
and UO_1530 (O_1530,N_14351,N_14601);
nor UO_1531 (O_1531,N_13808,N_14998);
nand UO_1532 (O_1532,N_14004,N_14671);
xnor UO_1533 (O_1533,N_14373,N_14510);
nand UO_1534 (O_1534,N_14224,N_14031);
nand UO_1535 (O_1535,N_14532,N_14168);
or UO_1536 (O_1536,N_13871,N_13524);
and UO_1537 (O_1537,N_13768,N_14812);
xnor UO_1538 (O_1538,N_13550,N_14878);
or UO_1539 (O_1539,N_13717,N_13617);
nor UO_1540 (O_1540,N_14201,N_13786);
and UO_1541 (O_1541,N_14266,N_13823);
and UO_1542 (O_1542,N_14605,N_13755);
xor UO_1543 (O_1543,N_14423,N_14799);
or UO_1544 (O_1544,N_13883,N_14486);
nand UO_1545 (O_1545,N_14017,N_13749);
nor UO_1546 (O_1546,N_14236,N_14389);
nor UO_1547 (O_1547,N_14237,N_14293);
and UO_1548 (O_1548,N_14310,N_14328);
xnor UO_1549 (O_1549,N_14886,N_14050);
nand UO_1550 (O_1550,N_13610,N_14526);
xnor UO_1551 (O_1551,N_14090,N_14763);
nand UO_1552 (O_1552,N_14783,N_14725);
or UO_1553 (O_1553,N_13682,N_13506);
nor UO_1554 (O_1554,N_14403,N_14555);
nor UO_1555 (O_1555,N_14213,N_13575);
nor UO_1556 (O_1556,N_14436,N_14936);
nand UO_1557 (O_1557,N_14358,N_14405);
xnor UO_1558 (O_1558,N_14041,N_14683);
nor UO_1559 (O_1559,N_14967,N_14600);
and UO_1560 (O_1560,N_13525,N_14253);
xnor UO_1561 (O_1561,N_14831,N_14697);
nand UO_1562 (O_1562,N_14479,N_13539);
nor UO_1563 (O_1563,N_13617,N_14385);
or UO_1564 (O_1564,N_13681,N_14126);
and UO_1565 (O_1565,N_13520,N_14284);
or UO_1566 (O_1566,N_13716,N_13564);
nand UO_1567 (O_1567,N_14099,N_14689);
and UO_1568 (O_1568,N_14197,N_13621);
and UO_1569 (O_1569,N_14247,N_14227);
and UO_1570 (O_1570,N_13629,N_14219);
or UO_1571 (O_1571,N_13799,N_14770);
and UO_1572 (O_1572,N_13918,N_13763);
nor UO_1573 (O_1573,N_14186,N_14972);
and UO_1574 (O_1574,N_13874,N_14965);
or UO_1575 (O_1575,N_13881,N_14071);
xnor UO_1576 (O_1576,N_14989,N_13669);
nor UO_1577 (O_1577,N_14377,N_13987);
nand UO_1578 (O_1578,N_14481,N_14962);
nand UO_1579 (O_1579,N_14550,N_14694);
or UO_1580 (O_1580,N_14611,N_14679);
and UO_1581 (O_1581,N_14815,N_13625);
xor UO_1582 (O_1582,N_14423,N_13759);
and UO_1583 (O_1583,N_13996,N_14368);
or UO_1584 (O_1584,N_14425,N_14377);
nor UO_1585 (O_1585,N_14130,N_14168);
nand UO_1586 (O_1586,N_14207,N_14981);
nor UO_1587 (O_1587,N_14061,N_14029);
nand UO_1588 (O_1588,N_13781,N_14950);
and UO_1589 (O_1589,N_14464,N_14471);
nand UO_1590 (O_1590,N_14674,N_13810);
nand UO_1591 (O_1591,N_14906,N_14598);
or UO_1592 (O_1592,N_14028,N_13851);
nor UO_1593 (O_1593,N_14426,N_14656);
or UO_1594 (O_1594,N_13988,N_14730);
nor UO_1595 (O_1595,N_13784,N_13909);
or UO_1596 (O_1596,N_14130,N_14065);
xnor UO_1597 (O_1597,N_14820,N_14094);
nor UO_1598 (O_1598,N_13718,N_14509);
nand UO_1599 (O_1599,N_14904,N_13842);
and UO_1600 (O_1600,N_14441,N_14861);
nor UO_1601 (O_1601,N_13984,N_14643);
nand UO_1602 (O_1602,N_13926,N_13968);
nor UO_1603 (O_1603,N_14091,N_14663);
or UO_1604 (O_1604,N_13550,N_14935);
and UO_1605 (O_1605,N_14261,N_14703);
or UO_1606 (O_1606,N_14106,N_13659);
nand UO_1607 (O_1607,N_14923,N_14122);
xor UO_1608 (O_1608,N_14311,N_14802);
nand UO_1609 (O_1609,N_14114,N_14488);
and UO_1610 (O_1610,N_14519,N_14762);
and UO_1611 (O_1611,N_13727,N_14166);
nand UO_1612 (O_1612,N_13865,N_13983);
xor UO_1613 (O_1613,N_14619,N_13726);
and UO_1614 (O_1614,N_14687,N_13512);
and UO_1615 (O_1615,N_14568,N_14454);
and UO_1616 (O_1616,N_14664,N_14922);
nand UO_1617 (O_1617,N_13638,N_14736);
and UO_1618 (O_1618,N_13549,N_13906);
xor UO_1619 (O_1619,N_14867,N_13533);
nand UO_1620 (O_1620,N_14724,N_14738);
xor UO_1621 (O_1621,N_14695,N_14423);
nand UO_1622 (O_1622,N_14946,N_14178);
nor UO_1623 (O_1623,N_13695,N_14195);
nor UO_1624 (O_1624,N_14691,N_14869);
nand UO_1625 (O_1625,N_14371,N_14391);
nor UO_1626 (O_1626,N_14385,N_14947);
nand UO_1627 (O_1627,N_13574,N_14504);
nor UO_1628 (O_1628,N_13520,N_14596);
or UO_1629 (O_1629,N_14913,N_14672);
or UO_1630 (O_1630,N_14875,N_13603);
and UO_1631 (O_1631,N_14249,N_13821);
xor UO_1632 (O_1632,N_13924,N_13630);
nand UO_1633 (O_1633,N_13698,N_14457);
xor UO_1634 (O_1634,N_14980,N_13972);
or UO_1635 (O_1635,N_14562,N_13997);
and UO_1636 (O_1636,N_14187,N_13640);
and UO_1637 (O_1637,N_14923,N_14557);
nor UO_1638 (O_1638,N_13755,N_14293);
or UO_1639 (O_1639,N_14222,N_13754);
xor UO_1640 (O_1640,N_14056,N_13594);
and UO_1641 (O_1641,N_14389,N_14562);
xor UO_1642 (O_1642,N_14178,N_14847);
or UO_1643 (O_1643,N_14898,N_14587);
and UO_1644 (O_1644,N_14530,N_14186);
xor UO_1645 (O_1645,N_14214,N_14885);
nand UO_1646 (O_1646,N_14225,N_14044);
or UO_1647 (O_1647,N_14168,N_13754);
nand UO_1648 (O_1648,N_13688,N_14883);
nor UO_1649 (O_1649,N_14295,N_13845);
and UO_1650 (O_1650,N_14691,N_14548);
xnor UO_1651 (O_1651,N_14617,N_13836);
nand UO_1652 (O_1652,N_14609,N_13681);
nor UO_1653 (O_1653,N_14753,N_14521);
nand UO_1654 (O_1654,N_13990,N_14324);
nand UO_1655 (O_1655,N_14826,N_13875);
nand UO_1656 (O_1656,N_13887,N_14575);
or UO_1657 (O_1657,N_13576,N_13975);
nand UO_1658 (O_1658,N_14018,N_14391);
nand UO_1659 (O_1659,N_14440,N_14783);
nand UO_1660 (O_1660,N_13960,N_14440);
nor UO_1661 (O_1661,N_14105,N_14754);
xor UO_1662 (O_1662,N_14318,N_14580);
and UO_1663 (O_1663,N_14963,N_14891);
or UO_1664 (O_1664,N_13709,N_14482);
and UO_1665 (O_1665,N_13664,N_13520);
nor UO_1666 (O_1666,N_14883,N_14487);
and UO_1667 (O_1667,N_13517,N_14183);
nor UO_1668 (O_1668,N_13724,N_13728);
nor UO_1669 (O_1669,N_14666,N_13971);
nor UO_1670 (O_1670,N_14569,N_14775);
xnor UO_1671 (O_1671,N_14713,N_14579);
and UO_1672 (O_1672,N_14158,N_14889);
or UO_1673 (O_1673,N_14079,N_14385);
nand UO_1674 (O_1674,N_14977,N_14162);
nand UO_1675 (O_1675,N_13808,N_13665);
nand UO_1676 (O_1676,N_13814,N_14339);
nor UO_1677 (O_1677,N_13666,N_13530);
nand UO_1678 (O_1678,N_13722,N_13841);
and UO_1679 (O_1679,N_14312,N_14366);
and UO_1680 (O_1680,N_14747,N_13577);
or UO_1681 (O_1681,N_13929,N_13522);
nor UO_1682 (O_1682,N_14348,N_14183);
nand UO_1683 (O_1683,N_14848,N_14788);
and UO_1684 (O_1684,N_13578,N_14044);
and UO_1685 (O_1685,N_13776,N_14629);
nor UO_1686 (O_1686,N_13556,N_14097);
xor UO_1687 (O_1687,N_13714,N_13976);
nor UO_1688 (O_1688,N_14600,N_14253);
xnor UO_1689 (O_1689,N_14972,N_14618);
nor UO_1690 (O_1690,N_14930,N_13582);
nor UO_1691 (O_1691,N_14060,N_14763);
and UO_1692 (O_1692,N_14072,N_14734);
nand UO_1693 (O_1693,N_13722,N_14541);
and UO_1694 (O_1694,N_14806,N_14954);
nand UO_1695 (O_1695,N_14314,N_14866);
xnor UO_1696 (O_1696,N_14141,N_13859);
nand UO_1697 (O_1697,N_13706,N_14504);
or UO_1698 (O_1698,N_13635,N_13742);
xnor UO_1699 (O_1699,N_13754,N_13692);
nor UO_1700 (O_1700,N_14078,N_14988);
or UO_1701 (O_1701,N_14739,N_14340);
xnor UO_1702 (O_1702,N_13878,N_14558);
nor UO_1703 (O_1703,N_13795,N_14865);
nor UO_1704 (O_1704,N_14828,N_14172);
nand UO_1705 (O_1705,N_14706,N_14798);
and UO_1706 (O_1706,N_14771,N_14586);
nor UO_1707 (O_1707,N_14557,N_13582);
or UO_1708 (O_1708,N_14699,N_14174);
and UO_1709 (O_1709,N_14081,N_14912);
nor UO_1710 (O_1710,N_14989,N_14169);
xnor UO_1711 (O_1711,N_13545,N_13960);
nor UO_1712 (O_1712,N_13729,N_13703);
or UO_1713 (O_1713,N_13890,N_13556);
nand UO_1714 (O_1714,N_14124,N_14446);
nand UO_1715 (O_1715,N_13883,N_13530);
and UO_1716 (O_1716,N_14512,N_14454);
nor UO_1717 (O_1717,N_14046,N_13956);
nor UO_1718 (O_1718,N_13932,N_14269);
nand UO_1719 (O_1719,N_14673,N_14795);
nor UO_1720 (O_1720,N_14284,N_14763);
nand UO_1721 (O_1721,N_14918,N_14329);
xor UO_1722 (O_1722,N_14213,N_13709);
and UO_1723 (O_1723,N_13518,N_14862);
xor UO_1724 (O_1724,N_13560,N_13886);
and UO_1725 (O_1725,N_13524,N_14934);
xnor UO_1726 (O_1726,N_13700,N_14887);
nand UO_1727 (O_1727,N_14134,N_14507);
xor UO_1728 (O_1728,N_13827,N_14791);
or UO_1729 (O_1729,N_14676,N_14138);
or UO_1730 (O_1730,N_14130,N_14624);
xor UO_1731 (O_1731,N_14694,N_13812);
and UO_1732 (O_1732,N_13949,N_13647);
nand UO_1733 (O_1733,N_14897,N_13740);
xor UO_1734 (O_1734,N_13915,N_14475);
xnor UO_1735 (O_1735,N_13751,N_14304);
nand UO_1736 (O_1736,N_14546,N_14011);
and UO_1737 (O_1737,N_14968,N_14026);
and UO_1738 (O_1738,N_14656,N_14400);
nand UO_1739 (O_1739,N_13585,N_14651);
or UO_1740 (O_1740,N_13864,N_14198);
nor UO_1741 (O_1741,N_13695,N_13787);
or UO_1742 (O_1742,N_14539,N_14190);
nand UO_1743 (O_1743,N_14354,N_14443);
and UO_1744 (O_1744,N_14695,N_14099);
and UO_1745 (O_1745,N_14248,N_14059);
nor UO_1746 (O_1746,N_14635,N_14489);
and UO_1747 (O_1747,N_13800,N_14768);
and UO_1748 (O_1748,N_14621,N_14486);
nand UO_1749 (O_1749,N_14613,N_13838);
and UO_1750 (O_1750,N_13926,N_14066);
nand UO_1751 (O_1751,N_14042,N_14267);
nor UO_1752 (O_1752,N_14186,N_14700);
xor UO_1753 (O_1753,N_13878,N_13768);
nor UO_1754 (O_1754,N_14360,N_13783);
xnor UO_1755 (O_1755,N_14304,N_13834);
or UO_1756 (O_1756,N_14404,N_14177);
nor UO_1757 (O_1757,N_14286,N_14436);
or UO_1758 (O_1758,N_14926,N_14138);
xor UO_1759 (O_1759,N_14026,N_13917);
nand UO_1760 (O_1760,N_14597,N_13902);
nor UO_1761 (O_1761,N_13930,N_14065);
nand UO_1762 (O_1762,N_14921,N_14969);
nor UO_1763 (O_1763,N_14202,N_13844);
nand UO_1764 (O_1764,N_14751,N_14762);
and UO_1765 (O_1765,N_14818,N_14212);
nor UO_1766 (O_1766,N_13852,N_13538);
or UO_1767 (O_1767,N_14404,N_13978);
and UO_1768 (O_1768,N_13927,N_14915);
nand UO_1769 (O_1769,N_14749,N_14845);
or UO_1770 (O_1770,N_14888,N_14770);
nor UO_1771 (O_1771,N_14119,N_14754);
and UO_1772 (O_1772,N_13819,N_14578);
nand UO_1773 (O_1773,N_14304,N_13729);
or UO_1774 (O_1774,N_13858,N_14700);
xnor UO_1775 (O_1775,N_14136,N_14342);
nand UO_1776 (O_1776,N_13996,N_13752);
nand UO_1777 (O_1777,N_14899,N_14384);
nor UO_1778 (O_1778,N_14244,N_14816);
and UO_1779 (O_1779,N_14955,N_13866);
and UO_1780 (O_1780,N_13558,N_14665);
nor UO_1781 (O_1781,N_14030,N_14083);
nand UO_1782 (O_1782,N_14559,N_13515);
and UO_1783 (O_1783,N_14760,N_14564);
xnor UO_1784 (O_1784,N_14507,N_13580);
or UO_1785 (O_1785,N_14853,N_14764);
or UO_1786 (O_1786,N_14860,N_14711);
nand UO_1787 (O_1787,N_14577,N_14287);
nand UO_1788 (O_1788,N_14818,N_14656);
xor UO_1789 (O_1789,N_13831,N_14804);
or UO_1790 (O_1790,N_13769,N_14993);
nor UO_1791 (O_1791,N_13790,N_13501);
nand UO_1792 (O_1792,N_14539,N_13586);
or UO_1793 (O_1793,N_13560,N_14698);
and UO_1794 (O_1794,N_14596,N_13779);
nor UO_1795 (O_1795,N_13981,N_13690);
xor UO_1796 (O_1796,N_14374,N_14569);
or UO_1797 (O_1797,N_14541,N_14265);
nor UO_1798 (O_1798,N_14790,N_14326);
or UO_1799 (O_1799,N_14963,N_14607);
nor UO_1800 (O_1800,N_14529,N_14575);
or UO_1801 (O_1801,N_14867,N_14941);
and UO_1802 (O_1802,N_13715,N_13560);
nand UO_1803 (O_1803,N_13605,N_14701);
nand UO_1804 (O_1804,N_14364,N_14729);
or UO_1805 (O_1805,N_14850,N_13546);
xor UO_1806 (O_1806,N_14944,N_13962);
and UO_1807 (O_1807,N_13685,N_14031);
nor UO_1808 (O_1808,N_13834,N_14348);
nor UO_1809 (O_1809,N_13574,N_14245);
xor UO_1810 (O_1810,N_14815,N_13754);
or UO_1811 (O_1811,N_13700,N_14796);
xor UO_1812 (O_1812,N_13613,N_13615);
xnor UO_1813 (O_1813,N_13602,N_14260);
or UO_1814 (O_1814,N_14909,N_13597);
xor UO_1815 (O_1815,N_14741,N_13808);
and UO_1816 (O_1816,N_14663,N_13730);
and UO_1817 (O_1817,N_14055,N_13600);
and UO_1818 (O_1818,N_14787,N_13902);
and UO_1819 (O_1819,N_14106,N_14480);
nand UO_1820 (O_1820,N_14633,N_13581);
xnor UO_1821 (O_1821,N_14582,N_14799);
nor UO_1822 (O_1822,N_14803,N_14658);
nor UO_1823 (O_1823,N_14972,N_14543);
or UO_1824 (O_1824,N_14180,N_14775);
or UO_1825 (O_1825,N_13916,N_14912);
xnor UO_1826 (O_1826,N_13649,N_13736);
or UO_1827 (O_1827,N_14942,N_14460);
and UO_1828 (O_1828,N_14945,N_14030);
nor UO_1829 (O_1829,N_13689,N_13838);
nand UO_1830 (O_1830,N_13953,N_14782);
nor UO_1831 (O_1831,N_13854,N_14508);
nand UO_1832 (O_1832,N_14727,N_14194);
nand UO_1833 (O_1833,N_13727,N_14084);
xor UO_1834 (O_1834,N_14397,N_14959);
or UO_1835 (O_1835,N_13941,N_14754);
xor UO_1836 (O_1836,N_14172,N_14344);
nand UO_1837 (O_1837,N_14645,N_14385);
nand UO_1838 (O_1838,N_13796,N_14445);
nor UO_1839 (O_1839,N_14102,N_14513);
nor UO_1840 (O_1840,N_14240,N_13508);
nor UO_1841 (O_1841,N_13645,N_14921);
or UO_1842 (O_1842,N_14283,N_14007);
or UO_1843 (O_1843,N_14415,N_14324);
or UO_1844 (O_1844,N_13666,N_14814);
xor UO_1845 (O_1845,N_13894,N_14291);
nor UO_1846 (O_1846,N_14132,N_14437);
or UO_1847 (O_1847,N_14147,N_14855);
and UO_1848 (O_1848,N_13849,N_14443);
nand UO_1849 (O_1849,N_14128,N_14908);
or UO_1850 (O_1850,N_13796,N_13854);
and UO_1851 (O_1851,N_13751,N_14888);
or UO_1852 (O_1852,N_13525,N_14314);
or UO_1853 (O_1853,N_13967,N_14693);
xor UO_1854 (O_1854,N_14001,N_14228);
and UO_1855 (O_1855,N_14494,N_14141);
or UO_1856 (O_1856,N_14309,N_14177);
nor UO_1857 (O_1857,N_13776,N_14017);
and UO_1858 (O_1858,N_14498,N_14631);
nand UO_1859 (O_1859,N_14969,N_14279);
xnor UO_1860 (O_1860,N_14469,N_13552);
nor UO_1861 (O_1861,N_14673,N_14507);
or UO_1862 (O_1862,N_13852,N_14176);
nand UO_1863 (O_1863,N_14291,N_14514);
or UO_1864 (O_1864,N_14386,N_14475);
nor UO_1865 (O_1865,N_14160,N_14041);
nand UO_1866 (O_1866,N_13845,N_13666);
nand UO_1867 (O_1867,N_14790,N_14009);
xor UO_1868 (O_1868,N_13695,N_13811);
xnor UO_1869 (O_1869,N_14676,N_14931);
xor UO_1870 (O_1870,N_14516,N_14612);
nand UO_1871 (O_1871,N_13725,N_14826);
and UO_1872 (O_1872,N_14642,N_13705);
xnor UO_1873 (O_1873,N_13547,N_14752);
nand UO_1874 (O_1874,N_13519,N_14392);
nor UO_1875 (O_1875,N_14233,N_13889);
or UO_1876 (O_1876,N_13735,N_14059);
or UO_1877 (O_1877,N_13575,N_14182);
or UO_1878 (O_1878,N_14838,N_14502);
and UO_1879 (O_1879,N_14592,N_13937);
nand UO_1880 (O_1880,N_14805,N_14763);
nand UO_1881 (O_1881,N_14660,N_14221);
nand UO_1882 (O_1882,N_14675,N_14732);
nor UO_1883 (O_1883,N_14961,N_14365);
nand UO_1884 (O_1884,N_14015,N_14333);
xnor UO_1885 (O_1885,N_14293,N_14624);
or UO_1886 (O_1886,N_14762,N_13788);
and UO_1887 (O_1887,N_14380,N_14387);
or UO_1888 (O_1888,N_14772,N_14783);
nand UO_1889 (O_1889,N_14643,N_14063);
or UO_1890 (O_1890,N_13512,N_14995);
nor UO_1891 (O_1891,N_14506,N_13574);
or UO_1892 (O_1892,N_14929,N_13766);
and UO_1893 (O_1893,N_14592,N_13573);
xnor UO_1894 (O_1894,N_13985,N_13803);
nor UO_1895 (O_1895,N_14417,N_14559);
nor UO_1896 (O_1896,N_13825,N_13733);
xnor UO_1897 (O_1897,N_14846,N_14550);
or UO_1898 (O_1898,N_13942,N_14215);
and UO_1899 (O_1899,N_13738,N_13636);
and UO_1900 (O_1900,N_14581,N_14900);
xnor UO_1901 (O_1901,N_13535,N_14829);
nand UO_1902 (O_1902,N_14358,N_13739);
nand UO_1903 (O_1903,N_13737,N_14275);
nand UO_1904 (O_1904,N_14538,N_13895);
or UO_1905 (O_1905,N_13702,N_13984);
xnor UO_1906 (O_1906,N_14699,N_14424);
nor UO_1907 (O_1907,N_14061,N_14871);
nand UO_1908 (O_1908,N_14720,N_13822);
xnor UO_1909 (O_1909,N_14646,N_14062);
nand UO_1910 (O_1910,N_14426,N_14187);
and UO_1911 (O_1911,N_14188,N_14852);
and UO_1912 (O_1912,N_14255,N_13855);
nand UO_1913 (O_1913,N_14836,N_14627);
xnor UO_1914 (O_1914,N_14648,N_14267);
or UO_1915 (O_1915,N_14246,N_13744);
nand UO_1916 (O_1916,N_14084,N_14739);
nand UO_1917 (O_1917,N_13846,N_14008);
nand UO_1918 (O_1918,N_13786,N_14916);
nand UO_1919 (O_1919,N_14716,N_14993);
or UO_1920 (O_1920,N_13949,N_14935);
and UO_1921 (O_1921,N_14976,N_13969);
and UO_1922 (O_1922,N_13933,N_14419);
nand UO_1923 (O_1923,N_14570,N_14263);
xor UO_1924 (O_1924,N_14943,N_14897);
nand UO_1925 (O_1925,N_14376,N_14339);
nand UO_1926 (O_1926,N_14259,N_13984);
or UO_1927 (O_1927,N_14594,N_13956);
nor UO_1928 (O_1928,N_14408,N_14533);
or UO_1929 (O_1929,N_14250,N_13883);
nor UO_1930 (O_1930,N_13715,N_14769);
nor UO_1931 (O_1931,N_13811,N_14214);
nor UO_1932 (O_1932,N_14744,N_14911);
or UO_1933 (O_1933,N_13646,N_14273);
nor UO_1934 (O_1934,N_13691,N_13638);
and UO_1935 (O_1935,N_14091,N_14243);
nand UO_1936 (O_1936,N_13627,N_14303);
nor UO_1937 (O_1937,N_13638,N_13692);
xor UO_1938 (O_1938,N_13500,N_13897);
nor UO_1939 (O_1939,N_14725,N_14599);
and UO_1940 (O_1940,N_14857,N_14955);
or UO_1941 (O_1941,N_13912,N_14475);
nor UO_1942 (O_1942,N_13992,N_13807);
and UO_1943 (O_1943,N_14490,N_14946);
xor UO_1944 (O_1944,N_13692,N_14118);
or UO_1945 (O_1945,N_14589,N_13941);
or UO_1946 (O_1946,N_13932,N_14991);
nand UO_1947 (O_1947,N_14853,N_13630);
xnor UO_1948 (O_1948,N_14018,N_13550);
nand UO_1949 (O_1949,N_14400,N_14628);
or UO_1950 (O_1950,N_13765,N_13572);
nand UO_1951 (O_1951,N_14164,N_14944);
nand UO_1952 (O_1952,N_13523,N_13857);
or UO_1953 (O_1953,N_14154,N_14196);
and UO_1954 (O_1954,N_14515,N_13588);
or UO_1955 (O_1955,N_13611,N_13778);
xnor UO_1956 (O_1956,N_14586,N_13790);
xor UO_1957 (O_1957,N_14881,N_13608);
nor UO_1958 (O_1958,N_13871,N_13930);
nor UO_1959 (O_1959,N_13793,N_13573);
xor UO_1960 (O_1960,N_14972,N_13965);
nor UO_1961 (O_1961,N_14412,N_13756);
nor UO_1962 (O_1962,N_14910,N_14985);
or UO_1963 (O_1963,N_13787,N_14596);
or UO_1964 (O_1964,N_14213,N_14911);
nand UO_1965 (O_1965,N_13726,N_14677);
or UO_1966 (O_1966,N_14119,N_13961);
nor UO_1967 (O_1967,N_13930,N_14034);
nor UO_1968 (O_1968,N_14000,N_14504);
xnor UO_1969 (O_1969,N_14461,N_14599);
xnor UO_1970 (O_1970,N_14987,N_14550);
nand UO_1971 (O_1971,N_14847,N_14000);
or UO_1972 (O_1972,N_13986,N_14300);
nor UO_1973 (O_1973,N_13751,N_14771);
nor UO_1974 (O_1974,N_14030,N_14704);
or UO_1975 (O_1975,N_14914,N_14072);
xor UO_1976 (O_1976,N_13853,N_14343);
xnor UO_1977 (O_1977,N_13741,N_13981);
nand UO_1978 (O_1978,N_14138,N_14509);
xor UO_1979 (O_1979,N_14093,N_14285);
or UO_1980 (O_1980,N_13523,N_13878);
xnor UO_1981 (O_1981,N_14039,N_14411);
and UO_1982 (O_1982,N_13596,N_13856);
nand UO_1983 (O_1983,N_14620,N_14602);
or UO_1984 (O_1984,N_14625,N_13870);
or UO_1985 (O_1985,N_13975,N_13741);
and UO_1986 (O_1986,N_14526,N_14382);
or UO_1987 (O_1987,N_14440,N_13504);
nor UO_1988 (O_1988,N_14010,N_14894);
or UO_1989 (O_1989,N_14700,N_14618);
or UO_1990 (O_1990,N_14420,N_13917);
nor UO_1991 (O_1991,N_14507,N_14777);
nand UO_1992 (O_1992,N_13843,N_13918);
nand UO_1993 (O_1993,N_13950,N_14635);
and UO_1994 (O_1994,N_13951,N_13748);
nand UO_1995 (O_1995,N_14696,N_13512);
xor UO_1996 (O_1996,N_14727,N_14884);
or UO_1997 (O_1997,N_13537,N_14585);
or UO_1998 (O_1998,N_14479,N_13641);
and UO_1999 (O_1999,N_14034,N_13558);
endmodule