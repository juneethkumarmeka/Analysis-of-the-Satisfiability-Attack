module basic_500_3000_500_6_levels_1xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_24,In_2);
nand U1 (N_1,In_421,In_99);
nor U2 (N_2,In_388,In_380);
nor U3 (N_3,In_453,In_191);
or U4 (N_4,In_32,In_349);
nor U5 (N_5,In_247,In_493);
nor U6 (N_6,In_298,In_224);
nand U7 (N_7,In_381,In_141);
or U8 (N_8,In_294,In_261);
nor U9 (N_9,In_74,In_184);
or U10 (N_10,In_179,In_375);
or U11 (N_11,In_254,In_389);
nand U12 (N_12,In_445,In_334);
or U13 (N_13,In_473,In_50);
nand U14 (N_14,In_277,In_156);
nand U15 (N_15,In_393,In_483);
and U16 (N_16,In_499,In_414);
nor U17 (N_17,In_171,In_409);
and U18 (N_18,In_283,In_237);
and U19 (N_19,In_385,In_5);
nor U20 (N_20,In_206,In_82);
or U21 (N_21,In_85,In_299);
nor U22 (N_22,In_96,In_29);
and U23 (N_23,In_266,In_244);
nor U24 (N_24,In_450,In_459);
or U25 (N_25,In_210,In_291);
nand U26 (N_26,In_316,In_371);
nor U27 (N_27,In_347,In_154);
nor U28 (N_28,In_423,In_91);
nor U29 (N_29,In_178,In_480);
and U30 (N_30,In_357,In_387);
nor U31 (N_31,In_458,In_286);
nor U32 (N_32,In_406,In_170);
or U33 (N_33,In_114,In_278);
nor U34 (N_34,In_489,In_163);
xnor U35 (N_35,In_331,In_84);
nand U36 (N_36,In_362,In_152);
or U37 (N_37,In_369,In_70);
and U38 (N_38,In_185,In_364);
nor U39 (N_39,In_255,In_465);
or U40 (N_40,In_494,In_83);
nor U41 (N_41,In_177,In_345);
and U42 (N_42,In_344,In_295);
and U43 (N_43,In_263,In_147);
or U44 (N_44,In_63,In_384);
nor U45 (N_45,In_399,In_352);
nand U46 (N_46,In_451,In_328);
and U47 (N_47,In_468,In_167);
and U48 (N_48,In_164,In_333);
nand U49 (N_49,In_319,In_322);
nand U50 (N_50,In_361,In_284);
nor U51 (N_51,In_73,In_422);
nor U52 (N_52,In_75,In_484);
nor U53 (N_53,In_72,In_78);
or U54 (N_54,In_300,In_466);
or U55 (N_55,In_27,In_95);
or U56 (N_56,In_7,In_123);
or U57 (N_57,In_208,In_374);
nand U58 (N_58,In_222,In_146);
nor U59 (N_59,In_281,In_241);
nand U60 (N_60,In_497,In_166);
or U61 (N_61,In_290,In_253);
and U62 (N_62,In_320,In_350);
nor U63 (N_63,In_193,In_6);
nand U64 (N_64,In_402,In_176);
or U65 (N_65,In_126,In_128);
and U66 (N_66,In_233,In_416);
nor U67 (N_67,In_348,In_418);
and U68 (N_68,In_61,In_228);
nor U69 (N_69,In_332,In_62);
nor U70 (N_70,In_94,In_80);
or U71 (N_71,In_410,In_433);
nand U72 (N_72,In_215,In_446);
and U73 (N_73,In_106,In_127);
or U74 (N_74,In_209,In_135);
nand U75 (N_75,In_77,In_205);
or U76 (N_76,In_162,In_113);
or U77 (N_77,In_47,In_4);
nand U78 (N_78,In_137,In_10);
nand U79 (N_79,In_59,In_462);
and U80 (N_80,In_153,In_190);
or U81 (N_81,In_330,In_150);
or U82 (N_82,In_377,In_46);
xor U83 (N_83,In_186,In_230);
nand U84 (N_84,In_432,In_67);
nand U85 (N_85,In_396,In_54);
nand U86 (N_86,In_58,In_256);
nor U87 (N_87,In_45,In_51);
or U88 (N_88,In_57,In_325);
nand U89 (N_89,In_76,In_492);
nand U90 (N_90,In_487,In_485);
and U91 (N_91,In_175,In_30);
nor U92 (N_92,In_33,In_340);
nor U93 (N_93,In_315,In_182);
nor U94 (N_94,In_417,In_69);
nand U95 (N_95,In_472,In_66);
nand U96 (N_96,In_274,In_343);
nor U97 (N_97,In_265,In_238);
or U98 (N_98,In_155,In_239);
nor U99 (N_99,In_460,In_216);
and U100 (N_100,In_447,In_86);
nand U101 (N_101,In_285,In_88);
nand U102 (N_102,In_207,In_194);
nor U103 (N_103,In_20,In_201);
or U104 (N_104,In_144,In_133);
or U105 (N_105,In_108,In_48);
or U106 (N_106,In_329,In_243);
nor U107 (N_107,In_313,In_386);
nand U108 (N_108,In_192,In_415);
and U109 (N_109,In_424,In_467);
or U110 (N_110,In_197,In_309);
nand U111 (N_111,In_165,In_49);
nor U112 (N_112,In_169,In_26);
or U113 (N_113,In_264,In_105);
or U114 (N_114,In_401,In_279);
nand U115 (N_115,In_246,In_172);
and U116 (N_116,In_41,In_436);
or U117 (N_117,In_488,In_0);
nand U118 (N_118,In_428,In_323);
nor U119 (N_119,In_435,In_9);
nor U120 (N_120,In_405,In_273);
and U121 (N_121,In_231,In_110);
and U122 (N_122,In_79,In_482);
and U123 (N_123,In_434,In_232);
xnor U124 (N_124,In_440,In_426);
and U125 (N_125,In_37,In_303);
nand U126 (N_126,In_287,In_275);
nand U127 (N_127,In_363,In_173);
or U128 (N_128,In_395,In_118);
and U129 (N_129,In_262,In_35);
or U130 (N_130,In_336,In_214);
nand U131 (N_131,In_203,In_109);
nor U132 (N_132,In_14,In_307);
and U133 (N_133,In_81,In_324);
nand U134 (N_134,In_202,In_36);
or U135 (N_135,In_317,In_444);
or U136 (N_136,In_71,In_431);
or U137 (N_137,In_200,In_370);
nor U138 (N_138,In_139,In_151);
nand U139 (N_139,In_116,In_55);
nand U140 (N_140,In_136,In_327);
nand U141 (N_141,In_65,In_93);
nand U142 (N_142,In_249,In_411);
and U143 (N_143,In_142,In_217);
and U144 (N_144,In_271,In_412);
nand U145 (N_145,In_476,In_188);
and U146 (N_146,In_21,In_270);
nor U147 (N_147,In_124,In_259);
nand U148 (N_148,In_251,In_280);
and U149 (N_149,In_8,In_293);
or U150 (N_150,In_353,In_227);
nor U151 (N_151,In_159,In_211);
nor U152 (N_152,In_23,In_22);
nand U153 (N_153,In_276,In_252);
or U154 (N_154,In_351,In_145);
and U155 (N_155,In_104,In_456);
nand U156 (N_156,In_408,In_15);
and U157 (N_157,In_3,In_346);
nor U158 (N_158,In_366,In_437);
nor U159 (N_159,In_143,In_360);
or U160 (N_160,In_398,In_103);
nor U161 (N_161,In_168,In_121);
and U162 (N_162,In_486,In_269);
nand U163 (N_163,In_111,In_199);
or U164 (N_164,In_394,In_301);
nor U165 (N_165,In_469,In_305);
or U166 (N_166,In_282,In_212);
nor U167 (N_167,In_187,In_52);
nand U168 (N_168,In_157,In_365);
nand U169 (N_169,In_267,In_454);
nand U170 (N_170,In_356,In_438);
or U171 (N_171,In_102,In_31);
nor U172 (N_172,In_314,In_268);
nor U173 (N_173,In_359,In_335);
nand U174 (N_174,In_318,In_220);
nand U175 (N_175,In_90,In_89);
or U176 (N_176,In_470,In_439);
or U177 (N_177,In_400,In_326);
nand U178 (N_178,In_260,In_1);
or U179 (N_179,In_463,In_296);
or U180 (N_180,In_443,In_373);
or U181 (N_181,In_478,In_97);
nor U182 (N_182,In_240,In_92);
nor U183 (N_183,In_180,In_42);
nor U184 (N_184,In_391,In_337);
and U185 (N_185,In_425,In_367);
nor U186 (N_186,In_310,In_496);
nand U187 (N_187,In_101,In_455);
and U188 (N_188,In_229,In_464);
or U189 (N_189,In_43,In_308);
nor U190 (N_190,In_196,In_429);
nand U191 (N_191,In_53,In_390);
or U192 (N_192,In_181,In_60);
or U193 (N_193,In_120,In_38);
and U194 (N_194,In_403,In_481);
or U195 (N_195,In_119,In_491);
and U196 (N_196,In_64,In_413);
nand U197 (N_197,In_297,In_132);
nand U198 (N_198,In_420,In_339);
and U199 (N_199,In_342,In_302);
nand U200 (N_200,In_183,In_131);
nor U201 (N_201,In_219,In_235);
nand U202 (N_202,In_248,In_404);
and U203 (N_203,In_321,In_204);
or U204 (N_204,In_148,In_441);
nor U205 (N_205,In_160,In_311);
or U206 (N_206,In_174,In_34);
or U207 (N_207,In_39,In_19);
or U208 (N_208,In_245,In_382);
or U209 (N_209,In_130,In_407);
nor U210 (N_210,In_461,In_448);
and U211 (N_211,In_198,In_213);
and U212 (N_212,In_258,In_475);
nor U213 (N_213,In_379,In_392);
nor U214 (N_214,In_18,In_419);
nor U215 (N_215,In_87,In_25);
nor U216 (N_216,In_122,In_16);
and U217 (N_217,In_479,In_355);
or U218 (N_218,In_341,In_138);
and U219 (N_219,In_13,In_44);
nand U220 (N_220,In_195,In_115);
and U221 (N_221,In_107,In_312);
or U222 (N_222,In_338,In_221);
or U223 (N_223,In_292,In_68);
or U224 (N_224,In_289,In_56);
nor U225 (N_225,In_452,In_189);
and U226 (N_226,In_140,In_223);
nand U227 (N_227,In_383,In_474);
xor U228 (N_228,In_112,In_218);
nand U229 (N_229,In_158,In_288);
or U230 (N_230,In_490,In_236);
or U231 (N_231,In_28,In_477);
and U232 (N_232,In_129,In_457);
nor U233 (N_233,In_134,In_354);
nor U234 (N_234,In_272,In_125);
and U235 (N_235,In_430,In_98);
and U236 (N_236,In_471,In_257);
and U237 (N_237,In_225,In_40);
and U238 (N_238,In_117,In_306);
or U239 (N_239,In_11,In_304);
or U240 (N_240,In_376,In_234);
nor U241 (N_241,In_397,In_226);
and U242 (N_242,In_149,In_250);
and U243 (N_243,In_161,In_449);
nand U244 (N_244,In_498,In_368);
or U245 (N_245,In_100,In_372);
nand U246 (N_246,In_242,In_12);
nand U247 (N_247,In_427,In_442);
and U248 (N_248,In_495,In_378);
and U249 (N_249,In_17,In_358);
nor U250 (N_250,In_35,In_213);
nand U251 (N_251,In_186,In_490);
and U252 (N_252,In_50,In_153);
and U253 (N_253,In_275,In_288);
nand U254 (N_254,In_413,In_183);
or U255 (N_255,In_117,In_497);
nor U256 (N_256,In_376,In_278);
nand U257 (N_257,In_111,In_243);
or U258 (N_258,In_426,In_200);
and U259 (N_259,In_391,In_388);
nor U260 (N_260,In_359,In_20);
or U261 (N_261,In_482,In_120);
nand U262 (N_262,In_312,In_369);
or U263 (N_263,In_383,In_305);
nand U264 (N_264,In_136,In_268);
nor U265 (N_265,In_399,In_453);
and U266 (N_266,In_381,In_53);
or U267 (N_267,In_198,In_104);
nor U268 (N_268,In_61,In_12);
nand U269 (N_269,In_315,In_265);
xor U270 (N_270,In_50,In_308);
or U271 (N_271,In_96,In_492);
nand U272 (N_272,In_109,In_23);
nor U273 (N_273,In_471,In_62);
nand U274 (N_274,In_431,In_362);
nand U275 (N_275,In_370,In_5);
nand U276 (N_276,In_411,In_5);
nor U277 (N_277,In_289,In_443);
or U278 (N_278,In_305,In_32);
or U279 (N_279,In_361,In_75);
or U280 (N_280,In_484,In_112);
or U281 (N_281,In_190,In_148);
and U282 (N_282,In_408,In_457);
or U283 (N_283,In_227,In_84);
and U284 (N_284,In_109,In_134);
and U285 (N_285,In_49,In_309);
nor U286 (N_286,In_443,In_211);
nand U287 (N_287,In_209,In_246);
nor U288 (N_288,In_195,In_78);
nor U289 (N_289,In_213,In_186);
nand U290 (N_290,In_238,In_140);
or U291 (N_291,In_244,In_415);
or U292 (N_292,In_57,In_338);
nand U293 (N_293,In_474,In_484);
and U294 (N_294,In_302,In_127);
nand U295 (N_295,In_293,In_378);
or U296 (N_296,In_154,In_255);
nand U297 (N_297,In_421,In_295);
or U298 (N_298,In_40,In_170);
nand U299 (N_299,In_8,In_339);
or U300 (N_300,In_143,In_98);
nand U301 (N_301,In_36,In_494);
nand U302 (N_302,In_444,In_311);
nand U303 (N_303,In_413,In_345);
nand U304 (N_304,In_165,In_352);
nand U305 (N_305,In_494,In_401);
or U306 (N_306,In_68,In_219);
nor U307 (N_307,In_324,In_208);
and U308 (N_308,In_223,In_389);
nor U309 (N_309,In_160,In_31);
nand U310 (N_310,In_356,In_465);
nand U311 (N_311,In_440,In_474);
nand U312 (N_312,In_261,In_484);
or U313 (N_313,In_445,In_122);
nor U314 (N_314,In_484,In_342);
and U315 (N_315,In_456,In_12);
nand U316 (N_316,In_62,In_321);
nand U317 (N_317,In_345,In_212);
and U318 (N_318,In_428,In_89);
nand U319 (N_319,In_16,In_314);
and U320 (N_320,In_444,In_275);
nand U321 (N_321,In_41,In_300);
nor U322 (N_322,In_92,In_32);
nand U323 (N_323,In_111,In_47);
or U324 (N_324,In_32,In_149);
and U325 (N_325,In_343,In_494);
and U326 (N_326,In_380,In_252);
nand U327 (N_327,In_452,In_77);
and U328 (N_328,In_247,In_8);
nor U329 (N_329,In_424,In_212);
and U330 (N_330,In_32,In_77);
xnor U331 (N_331,In_168,In_252);
nand U332 (N_332,In_147,In_400);
and U333 (N_333,In_351,In_199);
nand U334 (N_334,In_214,In_325);
nor U335 (N_335,In_427,In_488);
and U336 (N_336,In_354,In_160);
or U337 (N_337,In_406,In_480);
or U338 (N_338,In_480,In_227);
xor U339 (N_339,In_129,In_233);
nor U340 (N_340,In_83,In_111);
nor U341 (N_341,In_305,In_253);
nand U342 (N_342,In_182,In_187);
and U343 (N_343,In_169,In_300);
nand U344 (N_344,In_369,In_26);
and U345 (N_345,In_398,In_233);
and U346 (N_346,In_387,In_42);
nor U347 (N_347,In_375,In_15);
and U348 (N_348,In_449,In_202);
or U349 (N_349,In_146,In_462);
and U350 (N_350,In_136,In_86);
nand U351 (N_351,In_346,In_142);
or U352 (N_352,In_383,In_48);
or U353 (N_353,In_344,In_481);
nand U354 (N_354,In_115,In_391);
nand U355 (N_355,In_420,In_310);
or U356 (N_356,In_366,In_328);
xnor U357 (N_357,In_110,In_401);
nor U358 (N_358,In_454,In_367);
nand U359 (N_359,In_147,In_488);
nor U360 (N_360,In_217,In_216);
nor U361 (N_361,In_371,In_298);
nor U362 (N_362,In_212,In_258);
nor U363 (N_363,In_68,In_277);
nand U364 (N_364,In_306,In_198);
nand U365 (N_365,In_239,In_266);
and U366 (N_366,In_206,In_210);
nor U367 (N_367,In_96,In_441);
nor U368 (N_368,In_93,In_113);
and U369 (N_369,In_105,In_294);
nor U370 (N_370,In_355,In_83);
nand U371 (N_371,In_54,In_271);
nor U372 (N_372,In_104,In_229);
or U373 (N_373,In_386,In_396);
and U374 (N_374,In_23,In_132);
and U375 (N_375,In_141,In_260);
and U376 (N_376,In_458,In_78);
and U377 (N_377,In_385,In_26);
and U378 (N_378,In_370,In_43);
nor U379 (N_379,In_407,In_422);
or U380 (N_380,In_305,In_218);
or U381 (N_381,In_492,In_386);
or U382 (N_382,In_117,In_447);
nor U383 (N_383,In_488,In_435);
and U384 (N_384,In_418,In_430);
nand U385 (N_385,In_29,In_98);
and U386 (N_386,In_350,In_367);
and U387 (N_387,In_114,In_439);
and U388 (N_388,In_77,In_34);
nor U389 (N_389,In_9,In_88);
or U390 (N_390,In_269,In_283);
and U391 (N_391,In_7,In_148);
and U392 (N_392,In_178,In_92);
nor U393 (N_393,In_339,In_35);
or U394 (N_394,In_419,In_398);
nand U395 (N_395,In_56,In_223);
nor U396 (N_396,In_323,In_38);
nand U397 (N_397,In_14,In_230);
nand U398 (N_398,In_171,In_213);
and U399 (N_399,In_296,In_492);
nand U400 (N_400,In_278,In_323);
or U401 (N_401,In_492,In_377);
or U402 (N_402,In_28,In_226);
nand U403 (N_403,In_346,In_286);
and U404 (N_404,In_236,In_212);
nand U405 (N_405,In_499,In_151);
nor U406 (N_406,In_487,In_441);
nor U407 (N_407,In_118,In_382);
or U408 (N_408,In_455,In_10);
nor U409 (N_409,In_196,In_460);
and U410 (N_410,In_35,In_449);
nor U411 (N_411,In_66,In_342);
and U412 (N_412,In_252,In_1);
or U413 (N_413,In_119,In_442);
nand U414 (N_414,In_433,In_301);
and U415 (N_415,In_90,In_123);
nand U416 (N_416,In_293,In_493);
and U417 (N_417,In_13,In_370);
and U418 (N_418,In_465,In_423);
nor U419 (N_419,In_162,In_98);
or U420 (N_420,In_102,In_154);
nor U421 (N_421,In_152,In_348);
nor U422 (N_422,In_61,In_128);
and U423 (N_423,In_206,In_43);
nor U424 (N_424,In_393,In_74);
or U425 (N_425,In_161,In_53);
nand U426 (N_426,In_237,In_443);
nand U427 (N_427,In_199,In_165);
or U428 (N_428,In_229,In_252);
or U429 (N_429,In_243,In_90);
and U430 (N_430,In_13,In_126);
or U431 (N_431,In_468,In_125);
nor U432 (N_432,In_334,In_473);
nor U433 (N_433,In_371,In_89);
nand U434 (N_434,In_236,In_58);
or U435 (N_435,In_248,In_205);
nand U436 (N_436,In_333,In_346);
or U437 (N_437,In_81,In_99);
nand U438 (N_438,In_469,In_89);
nand U439 (N_439,In_422,In_429);
or U440 (N_440,In_393,In_422);
nand U441 (N_441,In_209,In_219);
and U442 (N_442,In_185,In_164);
and U443 (N_443,In_171,In_149);
nand U444 (N_444,In_296,In_424);
or U445 (N_445,In_165,In_258);
xor U446 (N_446,In_128,In_165);
nor U447 (N_447,In_57,In_18);
nor U448 (N_448,In_388,In_444);
and U449 (N_449,In_42,In_102);
nand U450 (N_450,In_113,In_30);
and U451 (N_451,In_314,In_34);
and U452 (N_452,In_467,In_434);
or U453 (N_453,In_475,In_276);
and U454 (N_454,In_49,In_99);
nand U455 (N_455,In_152,In_262);
and U456 (N_456,In_406,In_257);
nand U457 (N_457,In_221,In_98);
nor U458 (N_458,In_9,In_322);
or U459 (N_459,In_182,In_87);
nor U460 (N_460,In_367,In_133);
nor U461 (N_461,In_108,In_409);
or U462 (N_462,In_58,In_311);
nand U463 (N_463,In_428,In_339);
or U464 (N_464,In_78,In_337);
and U465 (N_465,In_369,In_419);
nor U466 (N_466,In_288,In_411);
and U467 (N_467,In_72,In_315);
or U468 (N_468,In_42,In_435);
and U469 (N_469,In_402,In_364);
and U470 (N_470,In_473,In_398);
nand U471 (N_471,In_469,In_470);
nand U472 (N_472,In_226,In_387);
or U473 (N_473,In_385,In_470);
nand U474 (N_474,In_156,In_407);
nor U475 (N_475,In_416,In_487);
nor U476 (N_476,In_139,In_273);
nand U477 (N_477,In_43,In_400);
and U478 (N_478,In_235,In_61);
and U479 (N_479,In_63,In_453);
or U480 (N_480,In_430,In_366);
nand U481 (N_481,In_251,In_452);
nand U482 (N_482,In_92,In_438);
or U483 (N_483,In_256,In_356);
nor U484 (N_484,In_419,In_215);
and U485 (N_485,In_417,In_253);
or U486 (N_486,In_311,In_132);
and U487 (N_487,In_485,In_360);
nand U488 (N_488,In_133,In_243);
xor U489 (N_489,In_304,In_362);
or U490 (N_490,In_43,In_422);
and U491 (N_491,In_179,In_363);
nor U492 (N_492,In_223,In_217);
and U493 (N_493,In_228,In_452);
and U494 (N_494,In_69,In_461);
nand U495 (N_495,In_422,In_167);
and U496 (N_496,In_328,In_412);
and U497 (N_497,In_404,In_43);
and U498 (N_498,In_339,In_299);
nand U499 (N_499,In_186,In_454);
nand U500 (N_500,N_412,N_259);
nor U501 (N_501,N_206,N_253);
nand U502 (N_502,N_75,N_317);
and U503 (N_503,N_233,N_213);
or U504 (N_504,N_3,N_303);
and U505 (N_505,N_389,N_214);
and U506 (N_506,N_394,N_332);
nand U507 (N_507,N_322,N_383);
and U508 (N_508,N_321,N_67);
nor U509 (N_509,N_313,N_151);
or U510 (N_510,N_226,N_441);
nand U511 (N_511,N_436,N_431);
or U512 (N_512,N_299,N_438);
or U513 (N_513,N_451,N_315);
and U514 (N_514,N_103,N_170);
xnor U515 (N_515,N_480,N_168);
nor U516 (N_516,N_23,N_49);
or U517 (N_517,N_97,N_335);
or U518 (N_518,N_93,N_160);
nand U519 (N_519,N_138,N_297);
and U520 (N_520,N_489,N_15);
nand U521 (N_521,N_413,N_24);
or U522 (N_522,N_109,N_347);
nor U523 (N_523,N_471,N_84);
nand U524 (N_524,N_352,N_384);
nor U525 (N_525,N_342,N_224);
nor U526 (N_526,N_266,N_429);
nor U527 (N_527,N_368,N_498);
nor U528 (N_528,N_407,N_123);
nor U529 (N_529,N_55,N_418);
or U530 (N_530,N_27,N_387);
and U531 (N_531,N_33,N_296);
and U532 (N_532,N_222,N_346);
or U533 (N_533,N_126,N_153);
nor U534 (N_534,N_98,N_4);
or U535 (N_535,N_240,N_223);
and U536 (N_536,N_295,N_403);
nand U537 (N_537,N_300,N_369);
nand U538 (N_538,N_398,N_255);
nor U539 (N_539,N_38,N_22);
nand U540 (N_540,N_169,N_89);
or U541 (N_541,N_125,N_218);
nor U542 (N_542,N_78,N_385);
and U543 (N_543,N_179,N_204);
or U544 (N_544,N_172,N_69);
and U545 (N_545,N_435,N_478);
nand U546 (N_546,N_455,N_227);
and U547 (N_547,N_469,N_499);
nand U548 (N_548,N_34,N_280);
or U549 (N_549,N_21,N_12);
or U550 (N_550,N_154,N_470);
nand U551 (N_551,N_492,N_50);
and U552 (N_552,N_239,N_488);
nand U553 (N_553,N_175,N_219);
or U554 (N_554,N_460,N_445);
nor U555 (N_555,N_462,N_28);
nor U556 (N_556,N_70,N_302);
or U557 (N_557,N_35,N_472);
nand U558 (N_558,N_272,N_85);
and U559 (N_559,N_304,N_9);
nor U560 (N_560,N_31,N_359);
nand U561 (N_561,N_159,N_156);
nor U562 (N_562,N_446,N_444);
or U563 (N_563,N_421,N_428);
and U564 (N_564,N_130,N_54);
nor U565 (N_565,N_29,N_107);
nand U566 (N_566,N_173,N_254);
or U567 (N_567,N_60,N_399);
nand U568 (N_568,N_201,N_132);
and U569 (N_569,N_207,N_152);
nand U570 (N_570,N_289,N_59);
nand U571 (N_571,N_419,N_329);
nor U572 (N_572,N_250,N_264);
or U573 (N_573,N_185,N_217);
or U574 (N_574,N_330,N_192);
nor U575 (N_575,N_113,N_479);
or U576 (N_576,N_162,N_442);
and U577 (N_577,N_281,N_366);
and U578 (N_578,N_124,N_376);
xor U579 (N_579,N_432,N_120);
or U580 (N_580,N_465,N_390);
nand U581 (N_581,N_102,N_181);
nand U582 (N_582,N_112,N_95);
or U583 (N_583,N_288,N_326);
nor U584 (N_584,N_450,N_423);
and U585 (N_585,N_88,N_294);
nand U586 (N_586,N_458,N_2);
nand U587 (N_587,N_232,N_251);
nand U588 (N_588,N_47,N_482);
nor U589 (N_589,N_453,N_65);
nand U590 (N_590,N_215,N_5);
nand U591 (N_591,N_16,N_490);
nand U592 (N_592,N_205,N_230);
nor U593 (N_593,N_41,N_196);
and U594 (N_594,N_468,N_312);
and U595 (N_595,N_496,N_497);
nand U596 (N_596,N_358,N_178);
nand U597 (N_597,N_210,N_475);
nand U598 (N_598,N_81,N_186);
or U599 (N_599,N_249,N_51);
and U600 (N_600,N_354,N_360);
and U601 (N_601,N_56,N_106);
and U602 (N_602,N_61,N_426);
nor U603 (N_603,N_94,N_150);
nor U604 (N_604,N_145,N_379);
nand U605 (N_605,N_344,N_286);
nor U606 (N_606,N_43,N_209);
nand U607 (N_607,N_386,N_375);
or U608 (N_608,N_314,N_293);
or U609 (N_609,N_66,N_339);
or U610 (N_610,N_447,N_108);
nand U611 (N_611,N_64,N_118);
or U612 (N_612,N_319,N_440);
nor U613 (N_613,N_324,N_305);
and U614 (N_614,N_269,N_381);
or U615 (N_615,N_284,N_80);
nand U616 (N_616,N_275,N_448);
nand U617 (N_617,N_62,N_278);
and U618 (N_618,N_271,N_474);
or U619 (N_619,N_466,N_393);
nor U620 (N_620,N_199,N_268);
and U621 (N_621,N_63,N_72);
nor U622 (N_622,N_433,N_486);
or U623 (N_623,N_191,N_237);
and U624 (N_624,N_211,N_323);
or U625 (N_625,N_245,N_270);
or U626 (N_626,N_76,N_142);
or U627 (N_627,N_414,N_307);
nor U628 (N_628,N_252,N_7);
or U629 (N_629,N_104,N_36);
nand U630 (N_630,N_92,N_87);
and U631 (N_631,N_262,N_96);
nand U632 (N_632,N_42,N_37);
nor U633 (N_633,N_17,N_361);
and U634 (N_634,N_157,N_267);
nand U635 (N_635,N_260,N_0);
or U636 (N_636,N_74,N_427);
or U637 (N_637,N_135,N_190);
nand U638 (N_638,N_114,N_309);
nand U639 (N_639,N_221,N_100);
and U640 (N_640,N_476,N_134);
and U641 (N_641,N_340,N_400);
nand U642 (N_642,N_131,N_422);
xnor U643 (N_643,N_424,N_147);
nor U644 (N_644,N_174,N_337);
or U645 (N_645,N_82,N_461);
and U646 (N_646,N_99,N_391);
nand U647 (N_647,N_495,N_164);
nor U648 (N_648,N_473,N_242);
nor U649 (N_649,N_32,N_325);
nand U650 (N_650,N_149,N_316);
and U651 (N_651,N_57,N_378);
nand U652 (N_652,N_208,N_333);
and U653 (N_653,N_200,N_158);
nor U654 (N_654,N_127,N_243);
nor U655 (N_655,N_443,N_203);
and U656 (N_656,N_417,N_18);
nor U657 (N_657,N_30,N_290);
nor U658 (N_658,N_265,N_276);
nand U659 (N_659,N_115,N_225);
and U660 (N_660,N_68,N_404);
nand U661 (N_661,N_128,N_183);
nor U662 (N_662,N_277,N_6);
nand U663 (N_663,N_416,N_353);
and U664 (N_664,N_212,N_189);
or U665 (N_665,N_44,N_248);
or U666 (N_666,N_463,N_238);
or U667 (N_667,N_246,N_167);
nor U668 (N_668,N_247,N_166);
nor U669 (N_669,N_318,N_148);
nand U670 (N_670,N_405,N_161);
and U671 (N_671,N_464,N_234);
and U672 (N_672,N_140,N_48);
nor U673 (N_673,N_373,N_367);
nand U674 (N_674,N_111,N_420);
or U675 (N_675,N_121,N_198);
and U676 (N_676,N_351,N_348);
and U677 (N_677,N_311,N_338);
or U678 (N_678,N_220,N_485);
nand U679 (N_679,N_341,N_256);
or U680 (N_680,N_439,N_229);
nand U681 (N_681,N_202,N_122);
nor U682 (N_682,N_40,N_14);
or U683 (N_683,N_292,N_144);
or U684 (N_684,N_53,N_494);
nor U685 (N_685,N_356,N_241);
nor U686 (N_686,N_146,N_45);
nand U687 (N_687,N_477,N_343);
and U688 (N_688,N_371,N_388);
or U689 (N_689,N_408,N_491);
nor U690 (N_690,N_110,N_236);
or U691 (N_691,N_197,N_415);
and U692 (N_692,N_77,N_137);
or U693 (N_693,N_392,N_334);
and U694 (N_694,N_263,N_52);
and U695 (N_695,N_397,N_449);
nor U696 (N_696,N_401,N_184);
or U697 (N_697,N_91,N_298);
and U698 (N_698,N_119,N_182);
nor U699 (N_699,N_493,N_411);
or U700 (N_700,N_39,N_155);
nand U701 (N_701,N_328,N_116);
or U702 (N_702,N_410,N_430);
nor U703 (N_703,N_180,N_336);
nor U704 (N_704,N_402,N_406);
nor U705 (N_705,N_20,N_117);
nand U706 (N_706,N_484,N_357);
and U707 (N_707,N_231,N_327);
or U708 (N_708,N_467,N_258);
or U709 (N_709,N_71,N_101);
and U710 (N_710,N_350,N_73);
or U711 (N_711,N_345,N_363);
or U712 (N_712,N_380,N_409);
or U713 (N_713,N_396,N_291);
nand U714 (N_714,N_310,N_46);
nand U715 (N_715,N_58,N_1);
or U716 (N_716,N_26,N_11);
or U717 (N_717,N_454,N_425);
nand U718 (N_718,N_195,N_193);
and U719 (N_719,N_457,N_13);
nor U720 (N_720,N_372,N_355);
and U721 (N_721,N_188,N_133);
nor U722 (N_722,N_19,N_481);
or U723 (N_723,N_306,N_487);
or U724 (N_724,N_279,N_365);
and U725 (N_725,N_136,N_331);
nor U726 (N_726,N_235,N_187);
nand U727 (N_727,N_176,N_143);
nor U728 (N_728,N_165,N_194);
and U729 (N_729,N_257,N_285);
nor U730 (N_730,N_283,N_261);
and U731 (N_731,N_8,N_370);
or U732 (N_732,N_90,N_320);
and U733 (N_733,N_163,N_382);
nand U734 (N_734,N_25,N_10);
or U735 (N_735,N_244,N_377);
nand U736 (N_736,N_437,N_349);
nand U737 (N_737,N_301,N_141);
or U738 (N_738,N_282,N_216);
and U739 (N_739,N_308,N_459);
and U740 (N_740,N_79,N_139);
nand U741 (N_741,N_171,N_228);
nor U742 (N_742,N_362,N_83);
nand U743 (N_743,N_105,N_434);
or U744 (N_744,N_274,N_287);
or U745 (N_745,N_129,N_452);
nand U746 (N_746,N_86,N_364);
and U747 (N_747,N_374,N_456);
or U748 (N_748,N_177,N_273);
nand U749 (N_749,N_395,N_483);
nand U750 (N_750,N_123,N_421);
nor U751 (N_751,N_0,N_154);
and U752 (N_752,N_119,N_239);
and U753 (N_753,N_114,N_442);
or U754 (N_754,N_413,N_250);
or U755 (N_755,N_486,N_243);
nor U756 (N_756,N_221,N_87);
and U757 (N_757,N_372,N_494);
and U758 (N_758,N_335,N_482);
and U759 (N_759,N_492,N_395);
nand U760 (N_760,N_20,N_434);
and U761 (N_761,N_434,N_283);
nand U762 (N_762,N_12,N_58);
or U763 (N_763,N_109,N_232);
or U764 (N_764,N_46,N_102);
nand U765 (N_765,N_117,N_126);
nand U766 (N_766,N_365,N_403);
nand U767 (N_767,N_54,N_322);
nor U768 (N_768,N_215,N_198);
and U769 (N_769,N_319,N_11);
or U770 (N_770,N_362,N_293);
or U771 (N_771,N_128,N_282);
and U772 (N_772,N_319,N_67);
nor U773 (N_773,N_7,N_198);
nand U774 (N_774,N_424,N_108);
nand U775 (N_775,N_242,N_320);
nor U776 (N_776,N_279,N_478);
nor U777 (N_777,N_398,N_325);
or U778 (N_778,N_58,N_402);
nor U779 (N_779,N_36,N_221);
nand U780 (N_780,N_438,N_477);
and U781 (N_781,N_62,N_221);
nand U782 (N_782,N_364,N_23);
and U783 (N_783,N_209,N_483);
or U784 (N_784,N_299,N_31);
and U785 (N_785,N_491,N_8);
nor U786 (N_786,N_407,N_466);
nor U787 (N_787,N_204,N_353);
or U788 (N_788,N_253,N_111);
nor U789 (N_789,N_13,N_391);
or U790 (N_790,N_145,N_158);
or U791 (N_791,N_420,N_56);
nor U792 (N_792,N_108,N_202);
and U793 (N_793,N_392,N_196);
or U794 (N_794,N_303,N_49);
and U795 (N_795,N_245,N_84);
nand U796 (N_796,N_96,N_355);
or U797 (N_797,N_407,N_435);
nand U798 (N_798,N_412,N_485);
or U799 (N_799,N_319,N_389);
nand U800 (N_800,N_120,N_203);
and U801 (N_801,N_430,N_113);
nor U802 (N_802,N_405,N_264);
nor U803 (N_803,N_118,N_48);
nor U804 (N_804,N_302,N_258);
or U805 (N_805,N_64,N_256);
xnor U806 (N_806,N_143,N_46);
and U807 (N_807,N_447,N_25);
and U808 (N_808,N_331,N_472);
nor U809 (N_809,N_191,N_495);
nand U810 (N_810,N_138,N_203);
nor U811 (N_811,N_335,N_1);
or U812 (N_812,N_252,N_143);
nand U813 (N_813,N_194,N_274);
nand U814 (N_814,N_78,N_72);
nand U815 (N_815,N_230,N_420);
nor U816 (N_816,N_43,N_259);
nor U817 (N_817,N_233,N_219);
nand U818 (N_818,N_59,N_421);
or U819 (N_819,N_170,N_360);
nor U820 (N_820,N_7,N_223);
or U821 (N_821,N_326,N_201);
or U822 (N_822,N_305,N_385);
nand U823 (N_823,N_180,N_126);
nand U824 (N_824,N_415,N_379);
nor U825 (N_825,N_308,N_446);
and U826 (N_826,N_182,N_12);
xor U827 (N_827,N_357,N_0);
nor U828 (N_828,N_113,N_31);
nor U829 (N_829,N_395,N_436);
and U830 (N_830,N_243,N_138);
or U831 (N_831,N_112,N_230);
xor U832 (N_832,N_173,N_139);
nor U833 (N_833,N_60,N_249);
or U834 (N_834,N_170,N_443);
nand U835 (N_835,N_139,N_136);
nor U836 (N_836,N_378,N_7);
nand U837 (N_837,N_98,N_189);
nand U838 (N_838,N_452,N_487);
or U839 (N_839,N_242,N_54);
nor U840 (N_840,N_37,N_294);
nor U841 (N_841,N_336,N_148);
nand U842 (N_842,N_139,N_287);
nor U843 (N_843,N_453,N_235);
nor U844 (N_844,N_117,N_94);
nor U845 (N_845,N_263,N_218);
and U846 (N_846,N_138,N_334);
and U847 (N_847,N_282,N_385);
nor U848 (N_848,N_15,N_433);
nand U849 (N_849,N_321,N_466);
or U850 (N_850,N_470,N_185);
or U851 (N_851,N_126,N_261);
and U852 (N_852,N_13,N_236);
and U853 (N_853,N_445,N_454);
and U854 (N_854,N_239,N_398);
or U855 (N_855,N_418,N_259);
nor U856 (N_856,N_15,N_20);
nand U857 (N_857,N_186,N_141);
and U858 (N_858,N_465,N_23);
nand U859 (N_859,N_67,N_316);
and U860 (N_860,N_41,N_167);
nor U861 (N_861,N_23,N_60);
nor U862 (N_862,N_376,N_394);
and U863 (N_863,N_171,N_371);
nand U864 (N_864,N_213,N_479);
nand U865 (N_865,N_276,N_50);
or U866 (N_866,N_348,N_275);
or U867 (N_867,N_375,N_151);
and U868 (N_868,N_266,N_1);
nand U869 (N_869,N_203,N_262);
nor U870 (N_870,N_464,N_394);
nand U871 (N_871,N_129,N_369);
nor U872 (N_872,N_90,N_360);
nand U873 (N_873,N_208,N_62);
nor U874 (N_874,N_456,N_159);
nor U875 (N_875,N_468,N_87);
nor U876 (N_876,N_417,N_94);
nand U877 (N_877,N_176,N_18);
nand U878 (N_878,N_131,N_428);
nand U879 (N_879,N_296,N_328);
nor U880 (N_880,N_383,N_301);
and U881 (N_881,N_228,N_461);
nand U882 (N_882,N_402,N_300);
nor U883 (N_883,N_362,N_393);
nor U884 (N_884,N_42,N_344);
nand U885 (N_885,N_22,N_256);
or U886 (N_886,N_314,N_16);
and U887 (N_887,N_84,N_392);
nand U888 (N_888,N_171,N_301);
and U889 (N_889,N_293,N_226);
nand U890 (N_890,N_53,N_400);
nand U891 (N_891,N_405,N_21);
nor U892 (N_892,N_4,N_381);
nor U893 (N_893,N_53,N_274);
nor U894 (N_894,N_346,N_60);
nand U895 (N_895,N_409,N_279);
and U896 (N_896,N_331,N_485);
and U897 (N_897,N_316,N_25);
and U898 (N_898,N_103,N_403);
or U899 (N_899,N_25,N_458);
nand U900 (N_900,N_135,N_424);
nand U901 (N_901,N_383,N_302);
and U902 (N_902,N_12,N_163);
nand U903 (N_903,N_68,N_470);
nor U904 (N_904,N_400,N_13);
nand U905 (N_905,N_234,N_386);
nor U906 (N_906,N_376,N_24);
or U907 (N_907,N_288,N_166);
nor U908 (N_908,N_368,N_193);
nand U909 (N_909,N_303,N_181);
nand U910 (N_910,N_490,N_386);
nor U911 (N_911,N_298,N_144);
nand U912 (N_912,N_204,N_380);
or U913 (N_913,N_280,N_133);
nor U914 (N_914,N_222,N_176);
nor U915 (N_915,N_133,N_257);
and U916 (N_916,N_1,N_26);
or U917 (N_917,N_431,N_325);
or U918 (N_918,N_126,N_21);
nand U919 (N_919,N_389,N_56);
or U920 (N_920,N_343,N_498);
nand U921 (N_921,N_59,N_189);
and U922 (N_922,N_109,N_62);
nand U923 (N_923,N_446,N_313);
nor U924 (N_924,N_180,N_345);
nand U925 (N_925,N_57,N_139);
nand U926 (N_926,N_272,N_243);
and U927 (N_927,N_468,N_36);
nand U928 (N_928,N_175,N_333);
nor U929 (N_929,N_266,N_402);
nor U930 (N_930,N_188,N_454);
and U931 (N_931,N_296,N_300);
nor U932 (N_932,N_325,N_118);
or U933 (N_933,N_192,N_44);
or U934 (N_934,N_272,N_314);
nor U935 (N_935,N_128,N_95);
nor U936 (N_936,N_464,N_468);
and U937 (N_937,N_238,N_384);
or U938 (N_938,N_181,N_84);
nand U939 (N_939,N_147,N_101);
nor U940 (N_940,N_135,N_28);
or U941 (N_941,N_445,N_262);
nand U942 (N_942,N_278,N_351);
or U943 (N_943,N_199,N_67);
and U944 (N_944,N_169,N_76);
and U945 (N_945,N_118,N_84);
nand U946 (N_946,N_207,N_329);
and U947 (N_947,N_242,N_223);
and U948 (N_948,N_426,N_228);
or U949 (N_949,N_50,N_2);
or U950 (N_950,N_39,N_367);
nor U951 (N_951,N_367,N_98);
and U952 (N_952,N_201,N_212);
and U953 (N_953,N_388,N_73);
nand U954 (N_954,N_335,N_378);
and U955 (N_955,N_329,N_144);
and U956 (N_956,N_292,N_301);
nand U957 (N_957,N_129,N_159);
or U958 (N_958,N_139,N_405);
nand U959 (N_959,N_430,N_22);
and U960 (N_960,N_74,N_408);
nor U961 (N_961,N_153,N_384);
nor U962 (N_962,N_179,N_258);
or U963 (N_963,N_423,N_65);
nor U964 (N_964,N_214,N_165);
and U965 (N_965,N_131,N_363);
or U966 (N_966,N_268,N_459);
nand U967 (N_967,N_223,N_492);
nand U968 (N_968,N_289,N_238);
or U969 (N_969,N_40,N_358);
and U970 (N_970,N_372,N_292);
nor U971 (N_971,N_464,N_40);
nor U972 (N_972,N_129,N_167);
nor U973 (N_973,N_155,N_271);
nor U974 (N_974,N_147,N_198);
or U975 (N_975,N_371,N_32);
and U976 (N_976,N_2,N_101);
or U977 (N_977,N_66,N_465);
nand U978 (N_978,N_76,N_110);
and U979 (N_979,N_175,N_13);
nor U980 (N_980,N_289,N_75);
or U981 (N_981,N_456,N_189);
nand U982 (N_982,N_90,N_22);
and U983 (N_983,N_254,N_26);
and U984 (N_984,N_49,N_333);
nand U985 (N_985,N_395,N_259);
nor U986 (N_986,N_23,N_53);
or U987 (N_987,N_464,N_347);
nand U988 (N_988,N_152,N_494);
or U989 (N_989,N_338,N_27);
nor U990 (N_990,N_173,N_109);
and U991 (N_991,N_20,N_447);
and U992 (N_992,N_360,N_418);
or U993 (N_993,N_296,N_41);
and U994 (N_994,N_1,N_139);
and U995 (N_995,N_469,N_89);
xnor U996 (N_996,N_392,N_202);
nand U997 (N_997,N_318,N_434);
nor U998 (N_998,N_408,N_24);
and U999 (N_999,N_258,N_226);
or U1000 (N_1000,N_538,N_631);
nor U1001 (N_1001,N_574,N_627);
or U1002 (N_1002,N_589,N_825);
and U1003 (N_1003,N_852,N_885);
and U1004 (N_1004,N_646,N_670);
nor U1005 (N_1005,N_613,N_565);
nor U1006 (N_1006,N_692,N_686);
or U1007 (N_1007,N_751,N_626);
or U1008 (N_1008,N_653,N_941);
nand U1009 (N_1009,N_520,N_904);
nor U1010 (N_1010,N_521,N_654);
and U1011 (N_1011,N_771,N_749);
or U1012 (N_1012,N_702,N_615);
or U1013 (N_1013,N_839,N_788);
or U1014 (N_1014,N_933,N_802);
or U1015 (N_1015,N_843,N_801);
nand U1016 (N_1016,N_898,N_918);
or U1017 (N_1017,N_951,N_674);
nor U1018 (N_1018,N_945,N_656);
nand U1019 (N_1019,N_551,N_546);
nor U1020 (N_1020,N_972,N_769);
and U1021 (N_1021,N_806,N_792);
nor U1022 (N_1022,N_633,N_803);
nand U1023 (N_1023,N_726,N_937);
and U1024 (N_1024,N_557,N_582);
or U1025 (N_1025,N_794,N_580);
nor U1026 (N_1026,N_955,N_638);
and U1027 (N_1027,N_598,N_710);
xnor U1028 (N_1028,N_840,N_900);
nor U1029 (N_1029,N_929,N_824);
or U1030 (N_1030,N_970,N_616);
nor U1031 (N_1031,N_872,N_628);
nand U1032 (N_1032,N_962,N_677);
and U1033 (N_1033,N_690,N_691);
nor U1034 (N_1034,N_735,N_657);
and U1035 (N_1035,N_780,N_555);
or U1036 (N_1036,N_581,N_781);
or U1037 (N_1037,N_925,N_560);
and U1038 (N_1038,N_684,N_655);
nor U1039 (N_1039,N_965,N_787);
nand U1040 (N_1040,N_664,N_876);
and U1041 (N_1041,N_992,N_608);
nand U1042 (N_1042,N_881,N_832);
nor U1043 (N_1043,N_807,N_879);
and U1044 (N_1044,N_948,N_562);
or U1045 (N_1045,N_525,N_734);
and U1046 (N_1046,N_821,N_812);
and U1047 (N_1047,N_896,N_540);
or U1048 (N_1048,N_770,N_682);
nor U1049 (N_1049,N_609,N_725);
nor U1050 (N_1050,N_901,N_916);
nor U1051 (N_1051,N_587,N_561);
or U1052 (N_1052,N_575,N_985);
and U1053 (N_1053,N_963,N_571);
and U1054 (N_1054,N_903,N_997);
nand U1055 (N_1055,N_535,N_886);
nand U1056 (N_1056,N_584,N_563);
or U1057 (N_1057,N_813,N_665);
or U1058 (N_1058,N_579,N_978);
nor U1059 (N_1059,N_758,N_741);
nand U1060 (N_1060,N_795,N_549);
nand U1061 (N_1061,N_658,N_515);
and U1062 (N_1062,N_651,N_636);
nor U1063 (N_1063,N_531,N_967);
nor U1064 (N_1064,N_714,N_661);
and U1065 (N_1065,N_891,N_688);
and U1066 (N_1066,N_796,N_974);
nand U1067 (N_1067,N_632,N_863);
nand U1068 (N_1068,N_827,N_991);
nand U1069 (N_1069,N_995,N_829);
or U1070 (N_1070,N_745,N_981);
or U1071 (N_1071,N_849,N_620);
or U1072 (N_1072,N_854,N_659);
or U1073 (N_1073,N_695,N_811);
and U1074 (N_1074,N_754,N_694);
nor U1075 (N_1075,N_953,N_585);
nor U1076 (N_1076,N_610,N_765);
or U1077 (N_1077,N_836,N_764);
and U1078 (N_1078,N_950,N_591);
nor U1079 (N_1079,N_946,N_680);
nand U1080 (N_1080,N_760,N_973);
or U1081 (N_1081,N_833,N_819);
nand U1082 (N_1082,N_921,N_982);
and U1083 (N_1083,N_858,N_957);
nand U1084 (N_1084,N_880,N_910);
nor U1085 (N_1085,N_782,N_569);
or U1086 (N_1086,N_502,N_869);
nand U1087 (N_1087,N_867,N_537);
and U1088 (N_1088,N_570,N_828);
nor U1089 (N_1089,N_855,N_547);
and U1090 (N_1090,N_823,N_697);
and U1091 (N_1091,N_786,N_737);
and U1092 (N_1092,N_789,N_588);
nor U1093 (N_1093,N_720,N_975);
or U1094 (N_1094,N_662,N_968);
nor U1095 (N_1095,N_922,N_911);
and U1096 (N_1096,N_919,N_504);
nand U1097 (N_1097,N_532,N_623);
nor U1098 (N_1098,N_920,N_503);
nand U1099 (N_1099,N_740,N_722);
or U1100 (N_1100,N_889,N_660);
and U1101 (N_1101,N_606,N_614);
or U1102 (N_1102,N_630,N_830);
nor U1103 (N_1103,N_597,N_791);
or U1104 (N_1104,N_550,N_507);
nor U1105 (N_1105,N_790,N_966);
nand U1106 (N_1106,N_592,N_558);
or U1107 (N_1107,N_988,N_862);
and U1108 (N_1108,N_681,N_753);
and U1109 (N_1109,N_835,N_524);
or U1110 (N_1110,N_939,N_809);
and U1111 (N_1111,N_719,N_645);
nand U1112 (N_1112,N_599,N_712);
or U1113 (N_1113,N_923,N_942);
nand U1114 (N_1114,N_882,N_528);
or U1115 (N_1115,N_698,N_913);
and U1116 (N_1116,N_508,N_800);
or U1117 (N_1117,N_912,N_993);
and U1118 (N_1118,N_730,N_757);
nor U1119 (N_1119,N_964,N_715);
nor U1120 (N_1120,N_746,N_642);
nand U1121 (N_1121,N_831,N_944);
or U1122 (N_1122,N_940,N_706);
nand U1123 (N_1123,N_938,N_685);
or U1124 (N_1124,N_994,N_568);
nor U1125 (N_1125,N_534,N_637);
nand U1126 (N_1126,N_894,N_977);
and U1127 (N_1127,N_530,N_527);
nand U1128 (N_1128,N_878,N_837);
nand U1129 (N_1129,N_639,N_999);
nand U1130 (N_1130,N_905,N_721);
nor U1131 (N_1131,N_986,N_793);
nor U1132 (N_1132,N_513,N_776);
xnor U1133 (N_1133,N_666,N_778);
nor U1134 (N_1134,N_871,N_518);
and U1135 (N_1135,N_577,N_853);
or U1136 (N_1136,N_506,N_756);
and U1137 (N_1137,N_625,N_516);
or U1138 (N_1138,N_750,N_818);
nor U1139 (N_1139,N_783,N_762);
nor U1140 (N_1140,N_731,N_509);
nand U1141 (N_1141,N_844,N_874);
nand U1142 (N_1142,N_583,N_600);
nand U1143 (N_1143,N_667,N_576);
and U1144 (N_1144,N_775,N_851);
nor U1145 (N_1145,N_621,N_897);
nor U1146 (N_1146,N_696,N_602);
nor U1147 (N_1147,N_596,N_888);
nand U1148 (N_1148,N_611,N_961);
nand U1149 (N_1149,N_554,N_564);
nand U1150 (N_1150,N_603,N_747);
nand U1151 (N_1151,N_728,N_777);
nand U1152 (N_1152,N_989,N_675);
nand U1153 (N_1153,N_672,N_541);
nand U1154 (N_1154,N_960,N_522);
nor U1155 (N_1155,N_622,N_542);
nor U1156 (N_1156,N_716,N_932);
or U1157 (N_1157,N_709,N_959);
and U1158 (N_1158,N_604,N_887);
and U1159 (N_1159,N_718,N_772);
or U1160 (N_1160,N_629,N_573);
nor U1161 (N_1161,N_805,N_890);
nor U1162 (N_1162,N_984,N_934);
nand U1163 (N_1163,N_924,N_971);
nand U1164 (N_1164,N_644,N_877);
nor U1165 (N_1165,N_703,N_906);
and U1166 (N_1166,N_536,N_847);
or U1167 (N_1167,N_908,N_768);
and U1168 (N_1168,N_701,N_822);
nand U1169 (N_1169,N_643,N_761);
nand U1170 (N_1170,N_567,N_669);
nand U1171 (N_1171,N_748,N_779);
and U1172 (N_1172,N_752,N_641);
nand U1173 (N_1173,N_875,N_586);
or U1174 (N_1174,N_935,N_505);
and U1175 (N_1175,N_711,N_566);
or U1176 (N_1176,N_733,N_958);
or U1177 (N_1177,N_907,N_744);
or U1178 (N_1178,N_511,N_866);
or U1179 (N_1179,N_859,N_857);
nor U1180 (N_1180,N_526,N_815);
nor U1181 (N_1181,N_713,N_607);
or U1182 (N_1182,N_652,N_671);
nor U1183 (N_1183,N_539,N_766);
nor U1184 (N_1184,N_553,N_699);
nor U1185 (N_1185,N_848,N_724);
and U1186 (N_1186,N_552,N_902);
nand U1187 (N_1187,N_846,N_826);
and U1188 (N_1188,N_729,N_817);
nand U1189 (N_1189,N_742,N_892);
nor U1190 (N_1190,N_868,N_861);
and U1191 (N_1191,N_842,N_884);
nand U1192 (N_1192,N_593,N_899);
nor U1193 (N_1193,N_545,N_914);
or U1194 (N_1194,N_949,N_917);
and U1195 (N_1195,N_727,N_990);
and U1196 (N_1196,N_605,N_808);
or U1197 (N_1197,N_601,N_928);
nand U1198 (N_1198,N_648,N_612);
nor U1199 (N_1199,N_804,N_936);
nor U1200 (N_1200,N_865,N_578);
nand U1201 (N_1201,N_523,N_705);
nor U1202 (N_1202,N_909,N_943);
and U1203 (N_1203,N_860,N_931);
or U1204 (N_1204,N_723,N_954);
nand U1205 (N_1205,N_785,N_883);
nand U1206 (N_1206,N_980,N_930);
and U1207 (N_1207,N_850,N_704);
and U1208 (N_1208,N_510,N_683);
and U1209 (N_1209,N_864,N_947);
nor U1210 (N_1210,N_634,N_996);
and U1211 (N_1211,N_895,N_987);
and U1212 (N_1212,N_700,N_514);
nand U1213 (N_1213,N_798,N_717);
and U1214 (N_1214,N_820,N_556);
and U1215 (N_1215,N_678,N_647);
and U1216 (N_1216,N_926,N_998);
nor U1217 (N_1217,N_693,N_927);
or U1218 (N_1218,N_763,N_687);
and U1219 (N_1219,N_799,N_640);
and U1220 (N_1220,N_755,N_797);
nor U1221 (N_1221,N_673,N_773);
and U1222 (N_1222,N_635,N_533);
nand U1223 (N_1223,N_834,N_501);
nand U1224 (N_1224,N_617,N_814);
nand U1225 (N_1225,N_624,N_544);
nand U1226 (N_1226,N_618,N_548);
or U1227 (N_1227,N_979,N_893);
nand U1228 (N_1228,N_668,N_873);
or U1229 (N_1229,N_708,N_983);
nand U1230 (N_1230,N_969,N_838);
or U1231 (N_1231,N_559,N_956);
and U1232 (N_1232,N_707,N_870);
or U1233 (N_1233,N_512,N_676);
or U1234 (N_1234,N_845,N_841);
nand U1235 (N_1235,N_816,N_650);
and U1236 (N_1236,N_500,N_519);
or U1237 (N_1237,N_572,N_689);
nor U1238 (N_1238,N_543,N_649);
and U1239 (N_1239,N_595,N_679);
or U1240 (N_1240,N_774,N_736);
nor U1241 (N_1241,N_529,N_952);
nor U1242 (N_1242,N_810,N_784);
nor U1243 (N_1243,N_594,N_590);
nor U1244 (N_1244,N_517,N_759);
nor U1245 (N_1245,N_739,N_619);
or U1246 (N_1246,N_767,N_732);
nor U1247 (N_1247,N_738,N_856);
and U1248 (N_1248,N_976,N_663);
or U1249 (N_1249,N_743,N_915);
nor U1250 (N_1250,N_721,N_913);
and U1251 (N_1251,N_512,N_771);
and U1252 (N_1252,N_854,N_767);
or U1253 (N_1253,N_887,N_997);
or U1254 (N_1254,N_735,N_530);
and U1255 (N_1255,N_670,N_775);
or U1256 (N_1256,N_614,N_680);
or U1257 (N_1257,N_554,N_709);
nor U1258 (N_1258,N_772,N_929);
nor U1259 (N_1259,N_697,N_580);
and U1260 (N_1260,N_889,N_799);
nand U1261 (N_1261,N_562,N_668);
and U1262 (N_1262,N_864,N_890);
nor U1263 (N_1263,N_864,N_843);
nor U1264 (N_1264,N_644,N_849);
or U1265 (N_1265,N_835,N_921);
and U1266 (N_1266,N_812,N_744);
nor U1267 (N_1267,N_606,N_552);
or U1268 (N_1268,N_729,N_958);
nor U1269 (N_1269,N_531,N_627);
and U1270 (N_1270,N_744,N_974);
and U1271 (N_1271,N_802,N_782);
and U1272 (N_1272,N_894,N_772);
nor U1273 (N_1273,N_500,N_997);
or U1274 (N_1274,N_570,N_802);
nand U1275 (N_1275,N_995,N_914);
nor U1276 (N_1276,N_879,N_869);
nand U1277 (N_1277,N_530,N_808);
nor U1278 (N_1278,N_847,N_721);
and U1279 (N_1279,N_654,N_828);
nand U1280 (N_1280,N_780,N_849);
nor U1281 (N_1281,N_739,N_749);
nand U1282 (N_1282,N_791,N_986);
and U1283 (N_1283,N_575,N_849);
nand U1284 (N_1284,N_879,N_545);
or U1285 (N_1285,N_652,N_810);
nand U1286 (N_1286,N_756,N_901);
nand U1287 (N_1287,N_987,N_958);
and U1288 (N_1288,N_523,N_781);
or U1289 (N_1289,N_622,N_752);
nor U1290 (N_1290,N_873,N_504);
and U1291 (N_1291,N_670,N_808);
or U1292 (N_1292,N_776,N_980);
nand U1293 (N_1293,N_693,N_978);
and U1294 (N_1294,N_500,N_741);
and U1295 (N_1295,N_698,N_750);
or U1296 (N_1296,N_640,N_930);
nand U1297 (N_1297,N_896,N_803);
or U1298 (N_1298,N_938,N_738);
nand U1299 (N_1299,N_947,N_607);
or U1300 (N_1300,N_580,N_565);
and U1301 (N_1301,N_966,N_923);
nor U1302 (N_1302,N_985,N_799);
or U1303 (N_1303,N_590,N_835);
nand U1304 (N_1304,N_773,N_629);
nand U1305 (N_1305,N_841,N_901);
nand U1306 (N_1306,N_508,N_560);
nand U1307 (N_1307,N_666,N_881);
or U1308 (N_1308,N_768,N_592);
nand U1309 (N_1309,N_952,N_798);
nand U1310 (N_1310,N_595,N_579);
nor U1311 (N_1311,N_785,N_891);
nand U1312 (N_1312,N_616,N_661);
nand U1313 (N_1313,N_552,N_660);
nand U1314 (N_1314,N_970,N_657);
nand U1315 (N_1315,N_920,N_744);
xnor U1316 (N_1316,N_555,N_840);
nor U1317 (N_1317,N_871,N_670);
or U1318 (N_1318,N_948,N_752);
xnor U1319 (N_1319,N_725,N_692);
and U1320 (N_1320,N_695,N_879);
nand U1321 (N_1321,N_682,N_564);
nand U1322 (N_1322,N_892,N_509);
nor U1323 (N_1323,N_737,N_525);
nor U1324 (N_1324,N_662,N_890);
nand U1325 (N_1325,N_718,N_952);
or U1326 (N_1326,N_770,N_920);
nor U1327 (N_1327,N_528,N_960);
nand U1328 (N_1328,N_726,N_632);
nor U1329 (N_1329,N_616,N_696);
nand U1330 (N_1330,N_818,N_656);
or U1331 (N_1331,N_663,N_511);
nor U1332 (N_1332,N_784,N_812);
or U1333 (N_1333,N_538,N_685);
or U1334 (N_1334,N_859,N_878);
nand U1335 (N_1335,N_558,N_889);
nand U1336 (N_1336,N_960,N_968);
or U1337 (N_1337,N_906,N_870);
and U1338 (N_1338,N_984,N_715);
and U1339 (N_1339,N_515,N_575);
nor U1340 (N_1340,N_796,N_583);
nor U1341 (N_1341,N_804,N_868);
nor U1342 (N_1342,N_955,N_587);
xor U1343 (N_1343,N_539,N_899);
and U1344 (N_1344,N_990,N_689);
nor U1345 (N_1345,N_695,N_864);
nand U1346 (N_1346,N_627,N_687);
nand U1347 (N_1347,N_890,N_638);
or U1348 (N_1348,N_961,N_745);
nand U1349 (N_1349,N_701,N_853);
nand U1350 (N_1350,N_989,N_522);
and U1351 (N_1351,N_521,N_514);
nor U1352 (N_1352,N_515,N_888);
xnor U1353 (N_1353,N_629,N_848);
nand U1354 (N_1354,N_792,N_563);
or U1355 (N_1355,N_912,N_902);
nor U1356 (N_1356,N_889,N_821);
nand U1357 (N_1357,N_565,N_957);
or U1358 (N_1358,N_794,N_817);
nand U1359 (N_1359,N_971,N_500);
nor U1360 (N_1360,N_826,N_689);
nor U1361 (N_1361,N_614,N_612);
and U1362 (N_1362,N_873,N_508);
nand U1363 (N_1363,N_531,N_686);
nand U1364 (N_1364,N_741,N_690);
nand U1365 (N_1365,N_855,N_969);
nand U1366 (N_1366,N_631,N_563);
nor U1367 (N_1367,N_995,N_586);
nor U1368 (N_1368,N_554,N_844);
nor U1369 (N_1369,N_887,N_569);
or U1370 (N_1370,N_964,N_530);
and U1371 (N_1371,N_558,N_752);
and U1372 (N_1372,N_700,N_745);
and U1373 (N_1373,N_899,N_615);
or U1374 (N_1374,N_657,N_545);
nor U1375 (N_1375,N_921,N_843);
nand U1376 (N_1376,N_745,N_841);
or U1377 (N_1377,N_929,N_685);
or U1378 (N_1378,N_994,N_516);
nor U1379 (N_1379,N_681,N_507);
and U1380 (N_1380,N_620,N_896);
or U1381 (N_1381,N_831,N_744);
and U1382 (N_1382,N_739,N_589);
and U1383 (N_1383,N_684,N_722);
nor U1384 (N_1384,N_931,N_583);
nor U1385 (N_1385,N_766,N_826);
nand U1386 (N_1386,N_851,N_946);
or U1387 (N_1387,N_997,N_833);
and U1388 (N_1388,N_650,N_998);
nor U1389 (N_1389,N_528,N_702);
nand U1390 (N_1390,N_596,N_575);
nor U1391 (N_1391,N_930,N_939);
or U1392 (N_1392,N_836,N_951);
xor U1393 (N_1393,N_619,N_605);
nand U1394 (N_1394,N_545,N_688);
nand U1395 (N_1395,N_615,N_571);
or U1396 (N_1396,N_661,N_889);
and U1397 (N_1397,N_650,N_528);
or U1398 (N_1398,N_782,N_537);
nor U1399 (N_1399,N_993,N_835);
nand U1400 (N_1400,N_911,N_918);
nor U1401 (N_1401,N_663,N_796);
nor U1402 (N_1402,N_751,N_852);
or U1403 (N_1403,N_671,N_951);
nand U1404 (N_1404,N_604,N_771);
and U1405 (N_1405,N_662,N_738);
nand U1406 (N_1406,N_904,N_985);
nor U1407 (N_1407,N_776,N_827);
and U1408 (N_1408,N_937,N_565);
nand U1409 (N_1409,N_903,N_582);
and U1410 (N_1410,N_637,N_672);
nor U1411 (N_1411,N_709,N_763);
nand U1412 (N_1412,N_840,N_501);
and U1413 (N_1413,N_608,N_603);
and U1414 (N_1414,N_574,N_677);
or U1415 (N_1415,N_506,N_893);
nand U1416 (N_1416,N_810,N_858);
nand U1417 (N_1417,N_583,N_850);
and U1418 (N_1418,N_699,N_978);
nand U1419 (N_1419,N_705,N_635);
nor U1420 (N_1420,N_848,N_922);
or U1421 (N_1421,N_507,N_789);
nor U1422 (N_1422,N_861,N_581);
and U1423 (N_1423,N_668,N_912);
nand U1424 (N_1424,N_788,N_927);
nor U1425 (N_1425,N_725,N_645);
and U1426 (N_1426,N_502,N_787);
nor U1427 (N_1427,N_513,N_706);
and U1428 (N_1428,N_797,N_653);
or U1429 (N_1429,N_832,N_755);
nand U1430 (N_1430,N_988,N_716);
and U1431 (N_1431,N_519,N_742);
nor U1432 (N_1432,N_670,N_634);
nand U1433 (N_1433,N_956,N_576);
nand U1434 (N_1434,N_687,N_534);
nand U1435 (N_1435,N_968,N_714);
nor U1436 (N_1436,N_986,N_522);
and U1437 (N_1437,N_923,N_985);
nor U1438 (N_1438,N_553,N_638);
nand U1439 (N_1439,N_591,N_941);
nor U1440 (N_1440,N_988,N_904);
or U1441 (N_1441,N_990,N_658);
nand U1442 (N_1442,N_523,N_845);
or U1443 (N_1443,N_853,N_909);
and U1444 (N_1444,N_558,N_623);
or U1445 (N_1445,N_766,N_570);
nand U1446 (N_1446,N_896,N_765);
nand U1447 (N_1447,N_886,N_825);
or U1448 (N_1448,N_543,N_951);
and U1449 (N_1449,N_751,N_878);
nor U1450 (N_1450,N_983,N_558);
or U1451 (N_1451,N_600,N_683);
or U1452 (N_1452,N_818,N_809);
nand U1453 (N_1453,N_925,N_602);
or U1454 (N_1454,N_668,N_503);
nand U1455 (N_1455,N_936,N_861);
or U1456 (N_1456,N_669,N_697);
or U1457 (N_1457,N_811,N_810);
nand U1458 (N_1458,N_904,N_686);
nand U1459 (N_1459,N_541,N_989);
nand U1460 (N_1460,N_748,N_836);
and U1461 (N_1461,N_719,N_576);
or U1462 (N_1462,N_568,N_920);
and U1463 (N_1463,N_689,N_620);
nand U1464 (N_1464,N_645,N_957);
nand U1465 (N_1465,N_813,N_778);
nand U1466 (N_1466,N_802,N_704);
nand U1467 (N_1467,N_589,N_620);
nor U1468 (N_1468,N_857,N_955);
nor U1469 (N_1469,N_987,N_930);
or U1470 (N_1470,N_799,N_681);
or U1471 (N_1471,N_646,N_520);
and U1472 (N_1472,N_539,N_994);
nor U1473 (N_1473,N_608,N_956);
nand U1474 (N_1474,N_554,N_643);
nand U1475 (N_1475,N_935,N_636);
and U1476 (N_1476,N_663,N_507);
and U1477 (N_1477,N_895,N_573);
and U1478 (N_1478,N_907,N_632);
or U1479 (N_1479,N_902,N_707);
and U1480 (N_1480,N_545,N_768);
and U1481 (N_1481,N_704,N_833);
and U1482 (N_1482,N_709,N_985);
nand U1483 (N_1483,N_695,N_640);
and U1484 (N_1484,N_736,N_864);
nor U1485 (N_1485,N_886,N_533);
or U1486 (N_1486,N_518,N_742);
nor U1487 (N_1487,N_652,N_935);
or U1488 (N_1488,N_670,N_680);
or U1489 (N_1489,N_625,N_970);
nand U1490 (N_1490,N_504,N_975);
nor U1491 (N_1491,N_553,N_783);
and U1492 (N_1492,N_652,N_578);
or U1493 (N_1493,N_771,N_522);
and U1494 (N_1494,N_608,N_611);
or U1495 (N_1495,N_941,N_563);
nand U1496 (N_1496,N_678,N_729);
or U1497 (N_1497,N_649,N_961);
nand U1498 (N_1498,N_513,N_775);
nand U1499 (N_1499,N_747,N_569);
and U1500 (N_1500,N_1069,N_1206);
and U1501 (N_1501,N_1433,N_1055);
xnor U1502 (N_1502,N_1041,N_1226);
nor U1503 (N_1503,N_1151,N_1390);
nor U1504 (N_1504,N_1033,N_1266);
nand U1505 (N_1505,N_1378,N_1026);
and U1506 (N_1506,N_1110,N_1246);
nor U1507 (N_1507,N_1254,N_1007);
nor U1508 (N_1508,N_1376,N_1495);
nor U1509 (N_1509,N_1317,N_1114);
nand U1510 (N_1510,N_1072,N_1261);
nand U1511 (N_1511,N_1112,N_1292);
and U1512 (N_1512,N_1490,N_1385);
nor U1513 (N_1513,N_1172,N_1077);
and U1514 (N_1514,N_1263,N_1352);
nand U1515 (N_1515,N_1207,N_1182);
nand U1516 (N_1516,N_1109,N_1068);
or U1517 (N_1517,N_1075,N_1479);
nor U1518 (N_1518,N_1361,N_1125);
or U1519 (N_1519,N_1475,N_1160);
and U1520 (N_1520,N_1059,N_1157);
nor U1521 (N_1521,N_1304,N_1186);
nand U1522 (N_1522,N_1228,N_1078);
nand U1523 (N_1523,N_1379,N_1375);
or U1524 (N_1524,N_1211,N_1076);
or U1525 (N_1525,N_1045,N_1168);
nor U1526 (N_1526,N_1034,N_1435);
nand U1527 (N_1527,N_1346,N_1382);
or U1528 (N_1528,N_1279,N_1159);
nor U1529 (N_1529,N_1024,N_1147);
nand U1530 (N_1530,N_1418,N_1188);
nand U1531 (N_1531,N_1103,N_1311);
and U1532 (N_1532,N_1025,N_1129);
and U1533 (N_1533,N_1058,N_1499);
and U1534 (N_1534,N_1067,N_1101);
nor U1535 (N_1535,N_1128,N_1054);
or U1536 (N_1536,N_1307,N_1403);
nand U1537 (N_1537,N_1194,N_1264);
or U1538 (N_1538,N_1015,N_1323);
nor U1539 (N_1539,N_1428,N_1008);
and U1540 (N_1540,N_1169,N_1117);
or U1541 (N_1541,N_1487,N_1011);
and U1542 (N_1542,N_1044,N_1448);
nor U1543 (N_1543,N_1404,N_1465);
nor U1544 (N_1544,N_1452,N_1464);
or U1545 (N_1545,N_1038,N_1371);
xor U1546 (N_1546,N_1231,N_1020);
nand U1547 (N_1547,N_1407,N_1486);
and U1548 (N_1548,N_1306,N_1272);
and U1549 (N_1549,N_1039,N_1043);
nor U1550 (N_1550,N_1130,N_1167);
and U1551 (N_1551,N_1256,N_1285);
nor U1552 (N_1552,N_1133,N_1402);
nor U1553 (N_1553,N_1003,N_1444);
nor U1554 (N_1554,N_1494,N_1190);
nand U1555 (N_1555,N_1210,N_1019);
and U1556 (N_1556,N_1267,N_1293);
and U1557 (N_1557,N_1155,N_1489);
nor U1558 (N_1558,N_1217,N_1380);
nand U1559 (N_1559,N_1295,N_1153);
nor U1560 (N_1560,N_1421,N_1368);
nor U1561 (N_1561,N_1126,N_1351);
and U1562 (N_1562,N_1337,N_1191);
and U1563 (N_1563,N_1431,N_1095);
nand U1564 (N_1564,N_1362,N_1203);
and U1565 (N_1565,N_1284,N_1181);
or U1566 (N_1566,N_1050,N_1199);
nand U1567 (N_1567,N_1123,N_1436);
and U1568 (N_1568,N_1184,N_1392);
or U1569 (N_1569,N_1189,N_1163);
and U1570 (N_1570,N_1111,N_1106);
nand U1571 (N_1571,N_1061,N_1331);
and U1572 (N_1572,N_1012,N_1460);
nor U1573 (N_1573,N_1056,N_1328);
nand U1574 (N_1574,N_1276,N_1088);
or U1575 (N_1575,N_1297,N_1350);
or U1576 (N_1576,N_1273,N_1238);
and U1577 (N_1577,N_1296,N_1455);
nor U1578 (N_1578,N_1250,N_1491);
nand U1579 (N_1579,N_1209,N_1442);
and U1580 (N_1580,N_1286,N_1073);
and U1581 (N_1581,N_1218,N_1329);
nor U1582 (N_1582,N_1013,N_1144);
nand U1583 (N_1583,N_1174,N_1298);
and U1584 (N_1584,N_1035,N_1330);
or U1585 (N_1585,N_1409,N_1274);
nand U1586 (N_1586,N_1426,N_1320);
and U1587 (N_1587,N_1367,N_1429);
and U1588 (N_1588,N_1332,N_1283);
nand U1589 (N_1589,N_1224,N_1419);
and U1590 (N_1590,N_1493,N_1430);
nor U1591 (N_1591,N_1481,N_1185);
or U1592 (N_1592,N_1200,N_1303);
nand U1593 (N_1593,N_1021,N_1253);
and U1594 (N_1594,N_1221,N_1242);
and U1595 (N_1595,N_1372,N_1417);
nand U1596 (N_1596,N_1258,N_1064);
nor U1597 (N_1597,N_1454,N_1247);
nor U1598 (N_1598,N_1023,N_1192);
nor U1599 (N_1599,N_1136,N_1288);
nand U1600 (N_1600,N_1420,N_1387);
and U1601 (N_1601,N_1441,N_1463);
or U1602 (N_1602,N_1170,N_1270);
and U1603 (N_1603,N_1269,N_1471);
nor U1604 (N_1604,N_1116,N_1108);
nor U1605 (N_1605,N_1383,N_1062);
xnor U1606 (N_1606,N_1156,N_1301);
nand U1607 (N_1607,N_1363,N_1085);
nor U1608 (N_1608,N_1300,N_1289);
and U1609 (N_1609,N_1498,N_1422);
nor U1610 (N_1610,N_1316,N_1333);
and U1611 (N_1611,N_1102,N_1259);
xor U1612 (N_1612,N_1215,N_1060);
or U1613 (N_1613,N_1115,N_1016);
or U1614 (N_1614,N_1036,N_1347);
or U1615 (N_1615,N_1173,N_1208);
or U1616 (N_1616,N_1083,N_1121);
nor U1617 (N_1617,N_1308,N_1080);
and U1618 (N_1618,N_1353,N_1314);
nor U1619 (N_1619,N_1017,N_1462);
nand U1620 (N_1620,N_1183,N_1029);
nand U1621 (N_1621,N_1355,N_1251);
or U1622 (N_1622,N_1240,N_1482);
or U1623 (N_1623,N_1252,N_1492);
nor U1624 (N_1624,N_1282,N_1434);
nand U1625 (N_1625,N_1040,N_1214);
nand U1626 (N_1626,N_1066,N_1398);
nor U1627 (N_1627,N_1090,N_1213);
nand U1628 (N_1628,N_1358,N_1234);
and U1629 (N_1629,N_1177,N_1022);
and U1630 (N_1630,N_1229,N_1394);
nand U1631 (N_1631,N_1180,N_1152);
nand U1632 (N_1632,N_1104,N_1423);
xnor U1633 (N_1633,N_1411,N_1414);
or U1634 (N_1634,N_1139,N_1082);
or U1635 (N_1635,N_1443,N_1193);
nor U1636 (N_1636,N_1357,N_1137);
or U1637 (N_1637,N_1063,N_1027);
and U1638 (N_1638,N_1374,N_1459);
nor U1639 (N_1639,N_1236,N_1389);
nor U1640 (N_1640,N_1053,N_1446);
nor U1641 (N_1641,N_1142,N_1205);
and U1642 (N_1642,N_1466,N_1294);
and U1643 (N_1643,N_1166,N_1388);
or U1644 (N_1644,N_1119,N_1412);
and U1645 (N_1645,N_1230,N_1065);
or U1646 (N_1646,N_1335,N_1094);
or U1647 (N_1647,N_1470,N_1440);
and U1648 (N_1648,N_1149,N_1453);
nand U1649 (N_1649,N_1483,N_1354);
nor U1650 (N_1650,N_1439,N_1049);
nand U1651 (N_1651,N_1140,N_1042);
or U1652 (N_1652,N_1406,N_1132);
or U1653 (N_1653,N_1410,N_1290);
nor U1654 (N_1654,N_1322,N_1212);
or U1655 (N_1655,N_1037,N_1449);
nand U1656 (N_1656,N_1164,N_1239);
nor U1657 (N_1657,N_1081,N_1310);
and U1658 (N_1658,N_1338,N_1241);
and U1659 (N_1659,N_1079,N_1091);
nand U1660 (N_1660,N_1396,N_1009);
or U1661 (N_1661,N_1478,N_1324);
nand U1662 (N_1662,N_1334,N_1348);
or U1663 (N_1663,N_1496,N_1148);
nor U1664 (N_1664,N_1291,N_1124);
nand U1665 (N_1665,N_1405,N_1196);
nor U1666 (N_1666,N_1235,N_1154);
nand U1667 (N_1667,N_1287,N_1366);
and U1668 (N_1668,N_1048,N_1223);
or U1669 (N_1669,N_1018,N_1339);
and U1670 (N_1670,N_1000,N_1315);
or U1671 (N_1671,N_1087,N_1086);
nand U1672 (N_1672,N_1399,N_1145);
or U1673 (N_1673,N_1245,N_1474);
and U1674 (N_1674,N_1175,N_1179);
nor U1675 (N_1675,N_1312,N_1299);
nor U1676 (N_1676,N_1178,N_1244);
nor U1677 (N_1677,N_1386,N_1084);
or U1678 (N_1678,N_1359,N_1447);
nand U1679 (N_1679,N_1467,N_1002);
or U1680 (N_1680,N_1318,N_1381);
nand U1681 (N_1681,N_1134,N_1401);
nor U1682 (N_1682,N_1198,N_1201);
nand U1683 (N_1683,N_1100,N_1135);
nor U1684 (N_1684,N_1360,N_1395);
nor U1685 (N_1685,N_1451,N_1051);
nor U1686 (N_1686,N_1400,N_1098);
xor U1687 (N_1687,N_1006,N_1262);
and U1688 (N_1688,N_1099,N_1227);
or U1689 (N_1689,N_1369,N_1195);
xor U1690 (N_1690,N_1171,N_1344);
or U1691 (N_1691,N_1005,N_1438);
or U1692 (N_1692,N_1365,N_1001);
or U1693 (N_1693,N_1349,N_1010);
nand U1694 (N_1694,N_1437,N_1118);
or U1695 (N_1695,N_1032,N_1071);
nor U1696 (N_1696,N_1278,N_1485);
nand U1697 (N_1697,N_1014,N_1319);
or U1698 (N_1698,N_1089,N_1197);
nand U1699 (N_1699,N_1424,N_1127);
or U1700 (N_1700,N_1074,N_1327);
or U1701 (N_1701,N_1477,N_1187);
and U1702 (N_1702,N_1220,N_1141);
or U1703 (N_1703,N_1302,N_1384);
and U1704 (N_1704,N_1497,N_1326);
and U1705 (N_1705,N_1165,N_1393);
or U1706 (N_1706,N_1468,N_1105);
or U1707 (N_1707,N_1397,N_1281);
xnor U1708 (N_1708,N_1216,N_1484);
or U1709 (N_1709,N_1120,N_1162);
or U1710 (N_1710,N_1237,N_1280);
or U1711 (N_1711,N_1321,N_1373);
nand U1712 (N_1712,N_1408,N_1249);
nor U1713 (N_1713,N_1057,N_1277);
and U1714 (N_1714,N_1243,N_1313);
or U1715 (N_1715,N_1309,N_1030);
or U1716 (N_1716,N_1204,N_1047);
nor U1717 (N_1717,N_1265,N_1458);
and U1718 (N_1718,N_1416,N_1122);
or U1719 (N_1719,N_1222,N_1488);
nor U1720 (N_1720,N_1260,N_1342);
or U1721 (N_1721,N_1028,N_1031);
and U1722 (N_1722,N_1096,N_1143);
nand U1723 (N_1723,N_1425,N_1364);
nor U1724 (N_1724,N_1356,N_1131);
and U1725 (N_1725,N_1158,N_1255);
nor U1726 (N_1726,N_1092,N_1473);
nor U1727 (N_1727,N_1097,N_1138);
nor U1728 (N_1728,N_1268,N_1232);
or U1729 (N_1729,N_1248,N_1340);
and U1730 (N_1730,N_1219,N_1070);
nand U1731 (N_1731,N_1046,N_1341);
or U1732 (N_1732,N_1113,N_1325);
nand U1733 (N_1733,N_1052,N_1336);
and U1734 (N_1734,N_1432,N_1427);
nand U1735 (N_1735,N_1275,N_1107);
nor U1736 (N_1736,N_1461,N_1225);
or U1737 (N_1737,N_1233,N_1377);
nor U1738 (N_1738,N_1457,N_1472);
and U1739 (N_1739,N_1345,N_1161);
nand U1740 (N_1740,N_1343,N_1093);
nor U1741 (N_1741,N_1456,N_1391);
or U1742 (N_1742,N_1480,N_1415);
or U1743 (N_1743,N_1469,N_1176);
or U1744 (N_1744,N_1476,N_1257);
and U1745 (N_1745,N_1146,N_1202);
or U1746 (N_1746,N_1271,N_1450);
nor U1747 (N_1747,N_1445,N_1370);
nand U1748 (N_1748,N_1413,N_1305);
nor U1749 (N_1749,N_1004,N_1150);
nor U1750 (N_1750,N_1096,N_1146);
and U1751 (N_1751,N_1279,N_1014);
or U1752 (N_1752,N_1461,N_1380);
nand U1753 (N_1753,N_1193,N_1183);
or U1754 (N_1754,N_1321,N_1356);
nor U1755 (N_1755,N_1231,N_1274);
nor U1756 (N_1756,N_1358,N_1386);
nor U1757 (N_1757,N_1282,N_1152);
nand U1758 (N_1758,N_1427,N_1401);
nand U1759 (N_1759,N_1459,N_1277);
nor U1760 (N_1760,N_1349,N_1432);
and U1761 (N_1761,N_1487,N_1040);
nor U1762 (N_1762,N_1454,N_1134);
nand U1763 (N_1763,N_1179,N_1063);
and U1764 (N_1764,N_1131,N_1370);
or U1765 (N_1765,N_1280,N_1047);
and U1766 (N_1766,N_1462,N_1297);
xnor U1767 (N_1767,N_1451,N_1079);
nor U1768 (N_1768,N_1486,N_1441);
and U1769 (N_1769,N_1076,N_1074);
nand U1770 (N_1770,N_1320,N_1443);
or U1771 (N_1771,N_1014,N_1255);
nor U1772 (N_1772,N_1319,N_1189);
nor U1773 (N_1773,N_1059,N_1065);
nand U1774 (N_1774,N_1377,N_1022);
nand U1775 (N_1775,N_1450,N_1230);
nor U1776 (N_1776,N_1039,N_1410);
or U1777 (N_1777,N_1183,N_1496);
nand U1778 (N_1778,N_1433,N_1119);
or U1779 (N_1779,N_1317,N_1293);
or U1780 (N_1780,N_1395,N_1006);
nor U1781 (N_1781,N_1395,N_1199);
and U1782 (N_1782,N_1252,N_1222);
nor U1783 (N_1783,N_1346,N_1227);
or U1784 (N_1784,N_1497,N_1229);
nor U1785 (N_1785,N_1208,N_1261);
or U1786 (N_1786,N_1135,N_1349);
nor U1787 (N_1787,N_1433,N_1295);
nand U1788 (N_1788,N_1141,N_1310);
xnor U1789 (N_1789,N_1422,N_1141);
and U1790 (N_1790,N_1036,N_1056);
and U1791 (N_1791,N_1013,N_1217);
and U1792 (N_1792,N_1279,N_1224);
nand U1793 (N_1793,N_1444,N_1113);
nor U1794 (N_1794,N_1445,N_1336);
nor U1795 (N_1795,N_1499,N_1415);
and U1796 (N_1796,N_1462,N_1313);
or U1797 (N_1797,N_1173,N_1123);
nor U1798 (N_1798,N_1016,N_1333);
nor U1799 (N_1799,N_1187,N_1351);
or U1800 (N_1800,N_1003,N_1114);
and U1801 (N_1801,N_1486,N_1051);
or U1802 (N_1802,N_1382,N_1475);
nor U1803 (N_1803,N_1120,N_1292);
nand U1804 (N_1804,N_1037,N_1474);
and U1805 (N_1805,N_1231,N_1334);
nand U1806 (N_1806,N_1068,N_1465);
or U1807 (N_1807,N_1268,N_1306);
nor U1808 (N_1808,N_1145,N_1240);
nor U1809 (N_1809,N_1347,N_1356);
nand U1810 (N_1810,N_1088,N_1095);
nor U1811 (N_1811,N_1468,N_1483);
nand U1812 (N_1812,N_1432,N_1375);
and U1813 (N_1813,N_1304,N_1324);
nor U1814 (N_1814,N_1484,N_1387);
nand U1815 (N_1815,N_1102,N_1368);
or U1816 (N_1816,N_1233,N_1181);
and U1817 (N_1817,N_1469,N_1273);
or U1818 (N_1818,N_1368,N_1069);
or U1819 (N_1819,N_1071,N_1104);
or U1820 (N_1820,N_1436,N_1088);
xnor U1821 (N_1821,N_1397,N_1091);
or U1822 (N_1822,N_1274,N_1249);
nor U1823 (N_1823,N_1450,N_1231);
and U1824 (N_1824,N_1360,N_1312);
and U1825 (N_1825,N_1019,N_1141);
and U1826 (N_1826,N_1474,N_1000);
nor U1827 (N_1827,N_1459,N_1228);
and U1828 (N_1828,N_1217,N_1187);
nand U1829 (N_1829,N_1333,N_1023);
and U1830 (N_1830,N_1128,N_1175);
nor U1831 (N_1831,N_1395,N_1449);
nor U1832 (N_1832,N_1371,N_1114);
nand U1833 (N_1833,N_1330,N_1212);
and U1834 (N_1834,N_1472,N_1285);
or U1835 (N_1835,N_1287,N_1417);
nor U1836 (N_1836,N_1299,N_1446);
or U1837 (N_1837,N_1395,N_1466);
nor U1838 (N_1838,N_1355,N_1254);
nand U1839 (N_1839,N_1336,N_1205);
or U1840 (N_1840,N_1103,N_1336);
and U1841 (N_1841,N_1296,N_1168);
nand U1842 (N_1842,N_1426,N_1248);
nor U1843 (N_1843,N_1477,N_1339);
nand U1844 (N_1844,N_1485,N_1279);
nor U1845 (N_1845,N_1149,N_1106);
and U1846 (N_1846,N_1477,N_1176);
or U1847 (N_1847,N_1182,N_1226);
and U1848 (N_1848,N_1190,N_1390);
and U1849 (N_1849,N_1009,N_1203);
and U1850 (N_1850,N_1315,N_1150);
or U1851 (N_1851,N_1363,N_1047);
nand U1852 (N_1852,N_1285,N_1434);
nor U1853 (N_1853,N_1335,N_1136);
and U1854 (N_1854,N_1024,N_1446);
nand U1855 (N_1855,N_1109,N_1168);
or U1856 (N_1856,N_1311,N_1025);
nor U1857 (N_1857,N_1114,N_1089);
nor U1858 (N_1858,N_1252,N_1277);
or U1859 (N_1859,N_1497,N_1080);
and U1860 (N_1860,N_1368,N_1285);
or U1861 (N_1861,N_1443,N_1295);
nor U1862 (N_1862,N_1216,N_1344);
nand U1863 (N_1863,N_1487,N_1016);
nor U1864 (N_1864,N_1191,N_1127);
and U1865 (N_1865,N_1493,N_1414);
nand U1866 (N_1866,N_1386,N_1118);
or U1867 (N_1867,N_1317,N_1031);
xnor U1868 (N_1868,N_1081,N_1470);
and U1869 (N_1869,N_1289,N_1331);
or U1870 (N_1870,N_1363,N_1012);
and U1871 (N_1871,N_1339,N_1179);
nor U1872 (N_1872,N_1471,N_1167);
or U1873 (N_1873,N_1286,N_1065);
nand U1874 (N_1874,N_1093,N_1075);
nand U1875 (N_1875,N_1203,N_1134);
nor U1876 (N_1876,N_1344,N_1098);
xnor U1877 (N_1877,N_1145,N_1234);
or U1878 (N_1878,N_1385,N_1241);
nor U1879 (N_1879,N_1440,N_1116);
or U1880 (N_1880,N_1245,N_1156);
nor U1881 (N_1881,N_1337,N_1293);
or U1882 (N_1882,N_1306,N_1197);
and U1883 (N_1883,N_1194,N_1221);
or U1884 (N_1884,N_1241,N_1009);
and U1885 (N_1885,N_1314,N_1432);
and U1886 (N_1886,N_1496,N_1354);
nor U1887 (N_1887,N_1284,N_1267);
nor U1888 (N_1888,N_1005,N_1312);
nor U1889 (N_1889,N_1269,N_1235);
nand U1890 (N_1890,N_1140,N_1196);
and U1891 (N_1891,N_1194,N_1470);
nor U1892 (N_1892,N_1044,N_1498);
or U1893 (N_1893,N_1068,N_1334);
or U1894 (N_1894,N_1366,N_1100);
and U1895 (N_1895,N_1092,N_1399);
and U1896 (N_1896,N_1042,N_1341);
nor U1897 (N_1897,N_1191,N_1082);
nand U1898 (N_1898,N_1376,N_1087);
or U1899 (N_1899,N_1151,N_1303);
and U1900 (N_1900,N_1292,N_1295);
nor U1901 (N_1901,N_1047,N_1241);
or U1902 (N_1902,N_1130,N_1488);
or U1903 (N_1903,N_1221,N_1043);
nor U1904 (N_1904,N_1221,N_1029);
nor U1905 (N_1905,N_1328,N_1475);
nor U1906 (N_1906,N_1296,N_1480);
nand U1907 (N_1907,N_1218,N_1274);
or U1908 (N_1908,N_1030,N_1148);
nor U1909 (N_1909,N_1047,N_1136);
or U1910 (N_1910,N_1250,N_1160);
or U1911 (N_1911,N_1000,N_1326);
or U1912 (N_1912,N_1325,N_1309);
nor U1913 (N_1913,N_1491,N_1270);
nand U1914 (N_1914,N_1317,N_1464);
and U1915 (N_1915,N_1169,N_1061);
nand U1916 (N_1916,N_1344,N_1470);
or U1917 (N_1917,N_1199,N_1056);
nand U1918 (N_1918,N_1474,N_1460);
nand U1919 (N_1919,N_1108,N_1237);
nor U1920 (N_1920,N_1001,N_1236);
or U1921 (N_1921,N_1041,N_1322);
or U1922 (N_1922,N_1110,N_1268);
and U1923 (N_1923,N_1080,N_1037);
or U1924 (N_1924,N_1366,N_1036);
nand U1925 (N_1925,N_1433,N_1471);
nand U1926 (N_1926,N_1219,N_1491);
nor U1927 (N_1927,N_1122,N_1196);
nand U1928 (N_1928,N_1110,N_1417);
nand U1929 (N_1929,N_1321,N_1000);
or U1930 (N_1930,N_1086,N_1100);
or U1931 (N_1931,N_1456,N_1367);
or U1932 (N_1932,N_1298,N_1067);
and U1933 (N_1933,N_1357,N_1314);
and U1934 (N_1934,N_1397,N_1015);
nor U1935 (N_1935,N_1407,N_1225);
nand U1936 (N_1936,N_1010,N_1205);
nor U1937 (N_1937,N_1425,N_1322);
and U1938 (N_1938,N_1065,N_1217);
and U1939 (N_1939,N_1027,N_1337);
nand U1940 (N_1940,N_1160,N_1418);
nor U1941 (N_1941,N_1067,N_1378);
or U1942 (N_1942,N_1016,N_1239);
nor U1943 (N_1943,N_1006,N_1056);
nor U1944 (N_1944,N_1151,N_1165);
nand U1945 (N_1945,N_1212,N_1148);
and U1946 (N_1946,N_1326,N_1306);
nand U1947 (N_1947,N_1177,N_1039);
nand U1948 (N_1948,N_1145,N_1418);
or U1949 (N_1949,N_1031,N_1318);
and U1950 (N_1950,N_1050,N_1114);
nor U1951 (N_1951,N_1080,N_1374);
nand U1952 (N_1952,N_1024,N_1436);
nand U1953 (N_1953,N_1383,N_1495);
or U1954 (N_1954,N_1297,N_1135);
nor U1955 (N_1955,N_1469,N_1244);
or U1956 (N_1956,N_1406,N_1465);
and U1957 (N_1957,N_1309,N_1110);
and U1958 (N_1958,N_1105,N_1195);
nand U1959 (N_1959,N_1231,N_1373);
nand U1960 (N_1960,N_1080,N_1315);
xnor U1961 (N_1961,N_1244,N_1197);
xnor U1962 (N_1962,N_1185,N_1028);
or U1963 (N_1963,N_1057,N_1005);
nand U1964 (N_1964,N_1247,N_1457);
nand U1965 (N_1965,N_1263,N_1197);
and U1966 (N_1966,N_1132,N_1464);
xor U1967 (N_1967,N_1294,N_1107);
and U1968 (N_1968,N_1056,N_1456);
or U1969 (N_1969,N_1021,N_1364);
and U1970 (N_1970,N_1083,N_1145);
nor U1971 (N_1971,N_1121,N_1210);
nand U1972 (N_1972,N_1028,N_1025);
or U1973 (N_1973,N_1312,N_1488);
nand U1974 (N_1974,N_1013,N_1353);
and U1975 (N_1975,N_1290,N_1251);
nand U1976 (N_1976,N_1339,N_1080);
nor U1977 (N_1977,N_1373,N_1214);
xor U1978 (N_1978,N_1042,N_1423);
or U1979 (N_1979,N_1415,N_1173);
and U1980 (N_1980,N_1308,N_1263);
nand U1981 (N_1981,N_1364,N_1485);
and U1982 (N_1982,N_1065,N_1341);
xnor U1983 (N_1983,N_1458,N_1254);
and U1984 (N_1984,N_1129,N_1313);
nor U1985 (N_1985,N_1153,N_1362);
and U1986 (N_1986,N_1141,N_1379);
xnor U1987 (N_1987,N_1422,N_1023);
nand U1988 (N_1988,N_1152,N_1284);
and U1989 (N_1989,N_1127,N_1115);
and U1990 (N_1990,N_1248,N_1018);
nor U1991 (N_1991,N_1087,N_1252);
nand U1992 (N_1992,N_1071,N_1251);
xnor U1993 (N_1993,N_1390,N_1166);
nand U1994 (N_1994,N_1254,N_1077);
xnor U1995 (N_1995,N_1107,N_1068);
or U1996 (N_1996,N_1316,N_1012);
nor U1997 (N_1997,N_1205,N_1399);
or U1998 (N_1998,N_1287,N_1091);
and U1999 (N_1999,N_1187,N_1058);
or U2000 (N_2000,N_1949,N_1995);
and U2001 (N_2001,N_1842,N_1585);
or U2002 (N_2002,N_1718,N_1727);
and U2003 (N_2003,N_1890,N_1942);
or U2004 (N_2004,N_1661,N_1969);
nand U2005 (N_2005,N_1647,N_1902);
and U2006 (N_2006,N_1705,N_1852);
nor U2007 (N_2007,N_1572,N_1556);
nand U2008 (N_2008,N_1671,N_1526);
nand U2009 (N_2009,N_1606,N_1965);
nand U2010 (N_2010,N_1927,N_1602);
or U2011 (N_2011,N_1525,N_1990);
or U2012 (N_2012,N_1800,N_1924);
and U2013 (N_2013,N_1638,N_1695);
and U2014 (N_2014,N_1519,N_1713);
and U2015 (N_2015,N_1929,N_1825);
and U2016 (N_2016,N_1848,N_1616);
and U2017 (N_2017,N_1697,N_1684);
nand U2018 (N_2018,N_1515,N_1704);
nand U2019 (N_2019,N_1918,N_1652);
or U2020 (N_2020,N_1797,N_1945);
and U2021 (N_2021,N_1625,N_1829);
or U2022 (N_2022,N_1610,N_1617);
and U2023 (N_2023,N_1985,N_1845);
or U2024 (N_2024,N_1936,N_1582);
nor U2025 (N_2025,N_1916,N_1524);
or U2026 (N_2026,N_1788,N_1867);
and U2027 (N_2027,N_1898,N_1957);
nor U2028 (N_2028,N_1991,N_1590);
and U2029 (N_2029,N_1741,N_1812);
nand U2030 (N_2030,N_1873,N_1795);
nand U2031 (N_2031,N_1686,N_1874);
and U2032 (N_2032,N_1966,N_1931);
or U2033 (N_2033,N_1559,N_1920);
nand U2034 (N_2034,N_1939,N_1834);
nand U2035 (N_2035,N_1620,N_1659);
nor U2036 (N_2036,N_1921,N_1557);
and U2037 (N_2037,N_1553,N_1783);
and U2038 (N_2038,N_1778,N_1805);
and U2039 (N_2039,N_1643,N_1760);
nand U2040 (N_2040,N_1658,N_1635);
and U2041 (N_2041,N_1726,N_1640);
nand U2042 (N_2042,N_1978,N_1622);
or U2043 (N_2043,N_1974,N_1547);
nor U2044 (N_2044,N_1567,N_1979);
or U2045 (N_2045,N_1678,N_1598);
nor U2046 (N_2046,N_1619,N_1710);
or U2047 (N_2047,N_1782,N_1937);
and U2048 (N_2048,N_1796,N_1822);
nor U2049 (N_2049,N_1528,N_1709);
nand U2050 (N_2050,N_1993,N_1780);
and U2051 (N_2051,N_1531,N_1668);
and U2052 (N_2052,N_1592,N_1768);
and U2053 (N_2053,N_1802,N_1673);
or U2054 (N_2054,N_1753,N_1608);
and U2055 (N_2055,N_1880,N_1577);
or U2056 (N_2056,N_1779,N_1615);
nand U2057 (N_2057,N_1613,N_1910);
nor U2058 (N_2058,N_1682,N_1548);
or U2059 (N_2059,N_1892,N_1846);
or U2060 (N_2060,N_1561,N_1793);
nand U2061 (N_2061,N_1767,N_1500);
nor U2062 (N_2062,N_1715,N_1551);
nand U2063 (N_2063,N_1813,N_1792);
and U2064 (N_2064,N_1747,N_1568);
nor U2065 (N_2065,N_1830,N_1881);
nand U2066 (N_2066,N_1891,N_1909);
nor U2067 (N_2067,N_1955,N_1576);
or U2068 (N_2068,N_1662,N_1765);
nand U2069 (N_2069,N_1535,N_1807);
nand U2070 (N_2070,N_1972,N_1735);
or U2071 (N_2071,N_1683,N_1664);
and U2072 (N_2072,N_1959,N_1749);
nand U2073 (N_2073,N_1688,N_1968);
nand U2074 (N_2074,N_1850,N_1787);
nand U2075 (N_2075,N_1947,N_1626);
nand U2076 (N_2076,N_1511,N_1691);
or U2077 (N_2077,N_1772,N_1507);
and U2078 (N_2078,N_1893,N_1605);
nand U2079 (N_2079,N_1600,N_1611);
nor U2080 (N_2080,N_1895,N_1919);
nor U2081 (N_2081,N_1532,N_1948);
or U2082 (N_2082,N_1721,N_1984);
or U2083 (N_2083,N_1522,N_1998);
nor U2084 (N_2084,N_1618,N_1579);
nand U2085 (N_2085,N_1786,N_1657);
nor U2086 (N_2086,N_1868,N_1843);
and U2087 (N_2087,N_1630,N_1954);
and U2088 (N_2088,N_1733,N_1523);
and U2089 (N_2089,N_1756,N_1773);
nor U2090 (N_2090,N_1722,N_1975);
and U2091 (N_2091,N_1841,N_1837);
or U2092 (N_2092,N_1855,N_1856);
nand U2093 (N_2093,N_1963,N_1546);
or U2094 (N_2094,N_1899,N_1663);
nor U2095 (N_2095,N_1550,N_1989);
nor U2096 (N_2096,N_1934,N_1632);
and U2097 (N_2097,N_1903,N_1828);
nand U2098 (N_2098,N_1870,N_1791);
nor U2099 (N_2099,N_1516,N_1573);
nor U2100 (N_2100,N_1628,N_1708);
nand U2101 (N_2101,N_1701,N_1518);
or U2102 (N_2102,N_1588,N_1593);
and U2103 (N_2103,N_1956,N_1666);
nand U2104 (N_2104,N_1544,N_1723);
nor U2105 (N_2105,N_1700,N_1513);
and U2106 (N_2106,N_1818,N_1912);
and U2107 (N_2107,N_1575,N_1680);
and U2108 (N_2108,N_1614,N_1563);
nor U2109 (N_2109,N_1543,N_1504);
or U2110 (N_2110,N_1789,N_1992);
or U2111 (N_2111,N_1946,N_1997);
or U2112 (N_2112,N_1840,N_1816);
nand U2113 (N_2113,N_1521,N_1827);
and U2114 (N_2114,N_1624,N_1777);
and U2115 (N_2115,N_1871,N_1994);
or U2116 (N_2116,N_1764,N_1865);
nand U2117 (N_2117,N_1869,N_1915);
nor U2118 (N_2118,N_1886,N_1958);
and U2119 (N_2119,N_1669,N_1717);
nand U2120 (N_2120,N_1670,N_1694);
nor U2121 (N_2121,N_1542,N_1962);
and U2122 (N_2122,N_1970,N_1986);
nand U2123 (N_2123,N_1720,N_1569);
or U2124 (N_2124,N_1603,N_1736);
nor U2125 (N_2125,N_1923,N_1629);
or U2126 (N_2126,N_1784,N_1878);
nor U2127 (N_2127,N_1646,N_1885);
nand U2128 (N_2128,N_1862,N_1555);
nand U2129 (N_2129,N_1961,N_1739);
nor U2130 (N_2130,N_1501,N_1755);
nand U2131 (N_2131,N_1913,N_1766);
and U2132 (N_2132,N_1607,N_1505);
nand U2133 (N_2133,N_1545,N_1594);
nor U2134 (N_2134,N_1742,N_1861);
and U2135 (N_2135,N_1520,N_1960);
or U2136 (N_2136,N_1627,N_1687);
nand U2137 (N_2137,N_1637,N_1967);
or U2138 (N_2138,N_1982,N_1811);
and U2139 (N_2139,N_1769,N_1914);
or U2140 (N_2140,N_1716,N_1930);
or U2141 (N_2141,N_1844,N_1702);
or U2142 (N_2142,N_1552,N_1654);
nand U2143 (N_2143,N_1808,N_1571);
and U2144 (N_2144,N_1817,N_1771);
and U2145 (N_2145,N_1838,N_1774);
and U2146 (N_2146,N_1754,N_1743);
and U2147 (N_2147,N_1996,N_1884);
or U2148 (N_2148,N_1706,N_1578);
and U2149 (N_2149,N_1835,N_1847);
and U2150 (N_2150,N_1599,N_1584);
nand U2151 (N_2151,N_1724,N_1512);
nor U2152 (N_2152,N_1509,N_1536);
and U2153 (N_2153,N_1826,N_1514);
and U2154 (N_2154,N_1876,N_1656);
nand U2155 (N_2155,N_1679,N_1589);
or U2156 (N_2156,N_1751,N_1731);
nand U2157 (N_2157,N_1746,N_1650);
and U2158 (N_2158,N_1801,N_1866);
or U2159 (N_2159,N_1596,N_1888);
and U2160 (N_2160,N_1655,N_1860);
and U2161 (N_2161,N_1554,N_1950);
and U2162 (N_2162,N_1748,N_1623);
nand U2163 (N_2163,N_1642,N_1648);
and U2164 (N_2164,N_1824,N_1941);
nand U2165 (N_2165,N_1911,N_1908);
and U2166 (N_2166,N_1549,N_1570);
nor U2167 (N_2167,N_1711,N_1541);
nand U2168 (N_2168,N_1858,N_1758);
and U2169 (N_2169,N_1785,N_1665);
nor U2170 (N_2170,N_1639,N_1562);
and U2171 (N_2171,N_1601,N_1631);
nor U2172 (N_2172,N_1538,N_1904);
nand U2173 (N_2173,N_1539,N_1649);
nor U2174 (N_2174,N_1675,N_1667);
and U2175 (N_2175,N_1740,N_1566);
nor U2176 (N_2176,N_1759,N_1744);
nand U2177 (N_2177,N_1644,N_1928);
and U2178 (N_2178,N_1703,N_1879);
nand U2179 (N_2179,N_1776,N_1714);
and U2180 (N_2180,N_1988,N_1530);
or U2181 (N_2181,N_1728,N_1854);
nor U2182 (N_2182,N_1940,N_1853);
or U2183 (N_2183,N_1770,N_1636);
or U2184 (N_2184,N_1804,N_1537);
nor U2185 (N_2185,N_1732,N_1699);
nand U2186 (N_2186,N_1925,N_1729);
or U2187 (N_2187,N_1999,N_1690);
nand U2188 (N_2188,N_1534,N_1580);
or U2189 (N_2189,N_1897,N_1790);
nor U2190 (N_2190,N_1745,N_1685);
nor U2191 (N_2191,N_1973,N_1712);
nand U2192 (N_2192,N_1823,N_1604);
or U2193 (N_2193,N_1757,N_1612);
nand U2194 (N_2194,N_1595,N_1836);
and U2195 (N_2195,N_1815,N_1689);
and U2196 (N_2196,N_1810,N_1693);
nor U2197 (N_2197,N_1883,N_1952);
or U2198 (N_2198,N_1833,N_1634);
and U2199 (N_2199,N_1591,N_1981);
and U2200 (N_2200,N_1725,N_1849);
nand U2201 (N_2201,N_1574,N_1803);
and U2202 (N_2202,N_1506,N_1750);
nor U2203 (N_2203,N_1781,N_1763);
xnor U2204 (N_2204,N_1872,N_1877);
nor U2205 (N_2205,N_1887,N_1894);
nor U2206 (N_2206,N_1761,N_1560);
xor U2207 (N_2207,N_1677,N_1794);
nor U2208 (N_2208,N_1953,N_1660);
nand U2209 (N_2209,N_1583,N_1558);
nand U2210 (N_2210,N_1864,N_1889);
nand U2211 (N_2211,N_1821,N_1738);
or U2212 (N_2212,N_1900,N_1951);
nor U2213 (N_2213,N_1875,N_1932);
nor U2214 (N_2214,N_1933,N_1863);
or U2215 (N_2215,N_1653,N_1964);
or U2216 (N_2216,N_1737,N_1609);
nand U2217 (N_2217,N_1983,N_1882);
and U2218 (N_2218,N_1814,N_1674);
nor U2219 (N_2219,N_1806,N_1587);
nor U2220 (N_2220,N_1672,N_1832);
or U2221 (N_2221,N_1944,N_1819);
nor U2222 (N_2222,N_1859,N_1799);
or U2223 (N_2223,N_1633,N_1851);
nor U2224 (N_2224,N_1529,N_1935);
nand U2225 (N_2225,N_1676,N_1692);
and U2226 (N_2226,N_1831,N_1734);
or U2227 (N_2227,N_1762,N_1621);
or U2228 (N_2228,N_1540,N_1896);
nand U2229 (N_2229,N_1922,N_1752);
or U2230 (N_2230,N_1906,N_1597);
or U2231 (N_2231,N_1901,N_1820);
or U2232 (N_2232,N_1938,N_1508);
or U2233 (N_2233,N_1971,N_1839);
and U2234 (N_2234,N_1917,N_1926);
and U2235 (N_2235,N_1775,N_1586);
nand U2236 (N_2236,N_1581,N_1645);
and U2237 (N_2237,N_1527,N_1641);
nor U2238 (N_2238,N_1564,N_1707);
or U2239 (N_2239,N_1980,N_1510);
nor U2240 (N_2240,N_1976,N_1651);
and U2241 (N_2241,N_1905,N_1798);
nand U2242 (N_2242,N_1907,N_1696);
nand U2243 (N_2243,N_1987,N_1517);
nor U2244 (N_2244,N_1503,N_1681);
nand U2245 (N_2245,N_1533,N_1698);
nand U2246 (N_2246,N_1809,N_1977);
and U2247 (N_2247,N_1730,N_1857);
and U2248 (N_2248,N_1719,N_1565);
nor U2249 (N_2249,N_1943,N_1502);
and U2250 (N_2250,N_1871,N_1799);
nor U2251 (N_2251,N_1845,N_1930);
or U2252 (N_2252,N_1849,N_1966);
nand U2253 (N_2253,N_1667,N_1856);
and U2254 (N_2254,N_1756,N_1569);
xnor U2255 (N_2255,N_1646,N_1769);
and U2256 (N_2256,N_1856,N_1799);
and U2257 (N_2257,N_1606,N_1541);
nand U2258 (N_2258,N_1553,N_1704);
or U2259 (N_2259,N_1656,N_1811);
or U2260 (N_2260,N_1879,N_1914);
nand U2261 (N_2261,N_1606,N_1688);
and U2262 (N_2262,N_1517,N_1639);
nor U2263 (N_2263,N_1864,N_1986);
nand U2264 (N_2264,N_1887,N_1724);
and U2265 (N_2265,N_1804,N_1888);
nor U2266 (N_2266,N_1833,N_1803);
and U2267 (N_2267,N_1573,N_1813);
nor U2268 (N_2268,N_1670,N_1721);
and U2269 (N_2269,N_1951,N_1922);
and U2270 (N_2270,N_1848,N_1677);
or U2271 (N_2271,N_1586,N_1690);
or U2272 (N_2272,N_1982,N_1813);
and U2273 (N_2273,N_1745,N_1961);
nor U2274 (N_2274,N_1890,N_1651);
nor U2275 (N_2275,N_1989,N_1576);
and U2276 (N_2276,N_1859,N_1730);
nor U2277 (N_2277,N_1761,N_1996);
or U2278 (N_2278,N_1533,N_1977);
nor U2279 (N_2279,N_1996,N_1737);
nor U2280 (N_2280,N_1988,N_1979);
nand U2281 (N_2281,N_1514,N_1620);
nand U2282 (N_2282,N_1704,N_1919);
nor U2283 (N_2283,N_1692,N_1916);
and U2284 (N_2284,N_1838,N_1575);
nor U2285 (N_2285,N_1595,N_1715);
and U2286 (N_2286,N_1955,N_1919);
nor U2287 (N_2287,N_1654,N_1571);
nand U2288 (N_2288,N_1520,N_1915);
and U2289 (N_2289,N_1612,N_1762);
nor U2290 (N_2290,N_1783,N_1738);
nor U2291 (N_2291,N_1740,N_1730);
xor U2292 (N_2292,N_1697,N_1872);
xor U2293 (N_2293,N_1749,N_1619);
nand U2294 (N_2294,N_1895,N_1750);
and U2295 (N_2295,N_1969,N_1576);
or U2296 (N_2296,N_1880,N_1718);
nand U2297 (N_2297,N_1814,N_1955);
and U2298 (N_2298,N_1885,N_1903);
nand U2299 (N_2299,N_1918,N_1949);
or U2300 (N_2300,N_1850,N_1525);
nand U2301 (N_2301,N_1673,N_1773);
and U2302 (N_2302,N_1901,N_1571);
nand U2303 (N_2303,N_1891,N_1598);
or U2304 (N_2304,N_1855,N_1565);
or U2305 (N_2305,N_1896,N_1870);
or U2306 (N_2306,N_1932,N_1588);
and U2307 (N_2307,N_1818,N_1802);
or U2308 (N_2308,N_1537,N_1649);
or U2309 (N_2309,N_1923,N_1875);
and U2310 (N_2310,N_1633,N_1764);
nor U2311 (N_2311,N_1559,N_1911);
and U2312 (N_2312,N_1924,N_1755);
or U2313 (N_2313,N_1792,N_1509);
and U2314 (N_2314,N_1943,N_1566);
nor U2315 (N_2315,N_1633,N_1808);
or U2316 (N_2316,N_1817,N_1928);
and U2317 (N_2317,N_1768,N_1804);
nor U2318 (N_2318,N_1588,N_1918);
or U2319 (N_2319,N_1998,N_1699);
nor U2320 (N_2320,N_1907,N_1539);
nor U2321 (N_2321,N_1875,N_1950);
nand U2322 (N_2322,N_1729,N_1826);
nand U2323 (N_2323,N_1630,N_1846);
and U2324 (N_2324,N_1983,N_1979);
or U2325 (N_2325,N_1977,N_1872);
and U2326 (N_2326,N_1950,N_1881);
or U2327 (N_2327,N_1515,N_1936);
nand U2328 (N_2328,N_1548,N_1973);
and U2329 (N_2329,N_1591,N_1567);
nor U2330 (N_2330,N_1504,N_1861);
or U2331 (N_2331,N_1675,N_1746);
and U2332 (N_2332,N_1972,N_1503);
or U2333 (N_2333,N_1849,N_1964);
xor U2334 (N_2334,N_1598,N_1778);
or U2335 (N_2335,N_1529,N_1986);
nand U2336 (N_2336,N_1909,N_1847);
nand U2337 (N_2337,N_1897,N_1533);
or U2338 (N_2338,N_1670,N_1880);
and U2339 (N_2339,N_1942,N_1743);
nand U2340 (N_2340,N_1904,N_1719);
or U2341 (N_2341,N_1627,N_1729);
nand U2342 (N_2342,N_1591,N_1984);
nand U2343 (N_2343,N_1588,N_1727);
nand U2344 (N_2344,N_1858,N_1697);
nand U2345 (N_2345,N_1827,N_1804);
nor U2346 (N_2346,N_1695,N_1854);
nor U2347 (N_2347,N_1880,N_1743);
or U2348 (N_2348,N_1741,N_1717);
nand U2349 (N_2349,N_1972,N_1968);
nand U2350 (N_2350,N_1778,N_1737);
and U2351 (N_2351,N_1685,N_1833);
nor U2352 (N_2352,N_1744,N_1979);
and U2353 (N_2353,N_1711,N_1803);
nor U2354 (N_2354,N_1853,N_1609);
nand U2355 (N_2355,N_1694,N_1947);
and U2356 (N_2356,N_1974,N_1896);
or U2357 (N_2357,N_1655,N_1593);
and U2358 (N_2358,N_1765,N_1507);
nor U2359 (N_2359,N_1934,N_1534);
nor U2360 (N_2360,N_1515,N_1758);
nor U2361 (N_2361,N_1709,N_1574);
nand U2362 (N_2362,N_1638,N_1944);
nand U2363 (N_2363,N_1508,N_1681);
and U2364 (N_2364,N_1979,N_1616);
or U2365 (N_2365,N_1658,N_1962);
and U2366 (N_2366,N_1882,N_1832);
nor U2367 (N_2367,N_1845,N_1509);
nand U2368 (N_2368,N_1903,N_1510);
or U2369 (N_2369,N_1988,N_1852);
and U2370 (N_2370,N_1780,N_1532);
and U2371 (N_2371,N_1861,N_1751);
and U2372 (N_2372,N_1723,N_1787);
and U2373 (N_2373,N_1713,N_1628);
nor U2374 (N_2374,N_1613,N_1750);
nand U2375 (N_2375,N_1922,N_1717);
or U2376 (N_2376,N_1732,N_1709);
and U2377 (N_2377,N_1606,N_1801);
and U2378 (N_2378,N_1536,N_1797);
nand U2379 (N_2379,N_1969,N_1512);
and U2380 (N_2380,N_1762,N_1857);
nand U2381 (N_2381,N_1966,N_1583);
nand U2382 (N_2382,N_1883,N_1980);
xnor U2383 (N_2383,N_1759,N_1552);
and U2384 (N_2384,N_1568,N_1652);
and U2385 (N_2385,N_1820,N_1822);
nand U2386 (N_2386,N_1964,N_1837);
nor U2387 (N_2387,N_1790,N_1814);
and U2388 (N_2388,N_1573,N_1948);
nand U2389 (N_2389,N_1762,N_1707);
and U2390 (N_2390,N_1854,N_1963);
and U2391 (N_2391,N_1773,N_1914);
and U2392 (N_2392,N_1816,N_1617);
nand U2393 (N_2393,N_1768,N_1607);
or U2394 (N_2394,N_1743,N_1611);
nand U2395 (N_2395,N_1921,N_1722);
and U2396 (N_2396,N_1924,N_1571);
nand U2397 (N_2397,N_1655,N_1734);
nand U2398 (N_2398,N_1717,N_1543);
nand U2399 (N_2399,N_1501,N_1820);
nor U2400 (N_2400,N_1704,N_1702);
nand U2401 (N_2401,N_1702,N_1985);
or U2402 (N_2402,N_1695,N_1556);
xor U2403 (N_2403,N_1620,N_1959);
or U2404 (N_2404,N_1682,N_1629);
nor U2405 (N_2405,N_1890,N_1617);
or U2406 (N_2406,N_1911,N_1590);
or U2407 (N_2407,N_1757,N_1736);
or U2408 (N_2408,N_1879,N_1695);
nor U2409 (N_2409,N_1996,N_1785);
and U2410 (N_2410,N_1712,N_1904);
nor U2411 (N_2411,N_1533,N_1991);
and U2412 (N_2412,N_1777,N_1503);
and U2413 (N_2413,N_1694,N_1942);
and U2414 (N_2414,N_1510,N_1720);
nand U2415 (N_2415,N_1939,N_1723);
nor U2416 (N_2416,N_1608,N_1574);
nand U2417 (N_2417,N_1682,N_1551);
or U2418 (N_2418,N_1573,N_1601);
nor U2419 (N_2419,N_1934,N_1753);
nor U2420 (N_2420,N_1581,N_1509);
and U2421 (N_2421,N_1931,N_1911);
and U2422 (N_2422,N_1645,N_1858);
and U2423 (N_2423,N_1802,N_1900);
and U2424 (N_2424,N_1894,N_1598);
or U2425 (N_2425,N_1767,N_1606);
or U2426 (N_2426,N_1812,N_1839);
and U2427 (N_2427,N_1877,N_1559);
nand U2428 (N_2428,N_1768,N_1658);
and U2429 (N_2429,N_1980,N_1997);
nor U2430 (N_2430,N_1523,N_1824);
nor U2431 (N_2431,N_1611,N_1943);
and U2432 (N_2432,N_1655,N_1873);
and U2433 (N_2433,N_1958,N_1769);
nand U2434 (N_2434,N_1826,N_1946);
nand U2435 (N_2435,N_1761,N_1858);
nand U2436 (N_2436,N_1804,N_1998);
nor U2437 (N_2437,N_1885,N_1580);
and U2438 (N_2438,N_1964,N_1858);
nand U2439 (N_2439,N_1689,N_1842);
xnor U2440 (N_2440,N_1919,N_1775);
nand U2441 (N_2441,N_1917,N_1991);
nor U2442 (N_2442,N_1607,N_1954);
nor U2443 (N_2443,N_1792,N_1825);
nand U2444 (N_2444,N_1650,N_1532);
nor U2445 (N_2445,N_1962,N_1514);
nor U2446 (N_2446,N_1973,N_1578);
or U2447 (N_2447,N_1811,N_1864);
or U2448 (N_2448,N_1799,N_1782);
and U2449 (N_2449,N_1832,N_1913);
nor U2450 (N_2450,N_1862,N_1661);
and U2451 (N_2451,N_1953,N_1779);
or U2452 (N_2452,N_1958,N_1923);
nor U2453 (N_2453,N_1839,N_1728);
and U2454 (N_2454,N_1994,N_1978);
or U2455 (N_2455,N_1932,N_1505);
nand U2456 (N_2456,N_1636,N_1821);
or U2457 (N_2457,N_1665,N_1536);
nor U2458 (N_2458,N_1670,N_1734);
or U2459 (N_2459,N_1822,N_1737);
nand U2460 (N_2460,N_1822,N_1718);
nor U2461 (N_2461,N_1962,N_1583);
nand U2462 (N_2462,N_1505,N_1622);
nor U2463 (N_2463,N_1764,N_1833);
or U2464 (N_2464,N_1925,N_1870);
and U2465 (N_2465,N_1992,N_1761);
and U2466 (N_2466,N_1789,N_1936);
and U2467 (N_2467,N_1775,N_1650);
or U2468 (N_2468,N_1752,N_1877);
or U2469 (N_2469,N_1793,N_1754);
nand U2470 (N_2470,N_1869,N_1516);
nor U2471 (N_2471,N_1502,N_1588);
nand U2472 (N_2472,N_1757,N_1523);
nor U2473 (N_2473,N_1893,N_1946);
and U2474 (N_2474,N_1856,N_1947);
or U2475 (N_2475,N_1617,N_1712);
and U2476 (N_2476,N_1568,N_1660);
nor U2477 (N_2477,N_1846,N_1809);
or U2478 (N_2478,N_1778,N_1919);
nand U2479 (N_2479,N_1843,N_1819);
or U2480 (N_2480,N_1502,N_1959);
and U2481 (N_2481,N_1633,N_1992);
or U2482 (N_2482,N_1570,N_1824);
or U2483 (N_2483,N_1653,N_1640);
or U2484 (N_2484,N_1924,N_1592);
nand U2485 (N_2485,N_1732,N_1801);
or U2486 (N_2486,N_1838,N_1900);
or U2487 (N_2487,N_1852,N_1817);
or U2488 (N_2488,N_1901,N_1741);
and U2489 (N_2489,N_1916,N_1871);
and U2490 (N_2490,N_1629,N_1796);
or U2491 (N_2491,N_1762,N_1634);
nand U2492 (N_2492,N_1616,N_1698);
nor U2493 (N_2493,N_1635,N_1912);
and U2494 (N_2494,N_1717,N_1605);
and U2495 (N_2495,N_1774,N_1862);
nand U2496 (N_2496,N_1851,N_1950);
or U2497 (N_2497,N_1995,N_1924);
and U2498 (N_2498,N_1968,N_1949);
nand U2499 (N_2499,N_1642,N_1982);
nand U2500 (N_2500,N_2423,N_2127);
or U2501 (N_2501,N_2447,N_2422);
or U2502 (N_2502,N_2365,N_2151);
or U2503 (N_2503,N_2290,N_2246);
and U2504 (N_2504,N_2405,N_2400);
nor U2505 (N_2505,N_2213,N_2148);
and U2506 (N_2506,N_2368,N_2410);
and U2507 (N_2507,N_2175,N_2289);
nor U2508 (N_2508,N_2272,N_2321);
nor U2509 (N_2509,N_2179,N_2048);
and U2510 (N_2510,N_2444,N_2182);
or U2511 (N_2511,N_2378,N_2491);
nand U2512 (N_2512,N_2156,N_2011);
or U2513 (N_2513,N_2114,N_2055);
nor U2514 (N_2514,N_2295,N_2363);
or U2515 (N_2515,N_2432,N_2224);
or U2516 (N_2516,N_2379,N_2357);
and U2517 (N_2517,N_2210,N_2351);
and U2518 (N_2518,N_2040,N_2235);
nor U2519 (N_2519,N_2331,N_2384);
nand U2520 (N_2520,N_2307,N_2305);
and U2521 (N_2521,N_2031,N_2497);
nor U2522 (N_2522,N_2061,N_2406);
nor U2523 (N_2523,N_2338,N_2071);
nor U2524 (N_2524,N_2342,N_2292);
or U2525 (N_2525,N_2013,N_2177);
or U2526 (N_2526,N_2167,N_2471);
nor U2527 (N_2527,N_2385,N_2376);
nor U2528 (N_2528,N_2233,N_2125);
nand U2529 (N_2529,N_2395,N_2485);
and U2530 (N_2530,N_2077,N_2001);
or U2531 (N_2531,N_2032,N_2415);
or U2532 (N_2532,N_2117,N_2336);
and U2533 (N_2533,N_2064,N_2214);
nor U2534 (N_2534,N_2397,N_2411);
or U2535 (N_2535,N_2248,N_2195);
or U2536 (N_2536,N_2237,N_2147);
nand U2537 (N_2537,N_2154,N_2050);
nor U2538 (N_2538,N_2285,N_2204);
nor U2539 (N_2539,N_2129,N_2022);
or U2540 (N_2540,N_2315,N_2473);
and U2541 (N_2541,N_2312,N_2062);
and U2542 (N_2542,N_2468,N_2180);
nand U2543 (N_2543,N_2025,N_2197);
nor U2544 (N_2544,N_2058,N_2003);
or U2545 (N_2545,N_2329,N_2019);
and U2546 (N_2546,N_2082,N_2460);
nor U2547 (N_2547,N_2461,N_2344);
and U2548 (N_2548,N_2045,N_2449);
and U2549 (N_2549,N_2333,N_2222);
nand U2550 (N_2550,N_2486,N_2074);
nand U2551 (N_2551,N_2399,N_2206);
or U2552 (N_2552,N_2245,N_2083);
or U2553 (N_2553,N_2418,N_2260);
nor U2554 (N_2554,N_2402,N_2089);
nand U2555 (N_2555,N_2489,N_2115);
nor U2556 (N_2556,N_2116,N_2049);
nand U2557 (N_2557,N_2317,N_2421);
or U2558 (N_2558,N_2316,N_2067);
and U2559 (N_2559,N_2254,N_2106);
and U2560 (N_2560,N_2038,N_2141);
or U2561 (N_2561,N_2145,N_2030);
nand U2562 (N_2562,N_2036,N_2232);
nor U2563 (N_2563,N_2483,N_2161);
and U2564 (N_2564,N_2478,N_2476);
and U2565 (N_2565,N_2293,N_2322);
xor U2566 (N_2566,N_2092,N_2056);
nand U2567 (N_2567,N_2297,N_2446);
and U2568 (N_2568,N_2028,N_2269);
or U2569 (N_2569,N_2234,N_2466);
nor U2570 (N_2570,N_2018,N_2270);
and U2571 (N_2571,N_2291,N_2076);
nor U2572 (N_2572,N_2133,N_2226);
or U2573 (N_2573,N_2453,N_2169);
or U2574 (N_2574,N_2268,N_2079);
and U2575 (N_2575,N_2403,N_2173);
xnor U2576 (N_2576,N_2455,N_2241);
or U2577 (N_2577,N_2209,N_2371);
nor U2578 (N_2578,N_2484,N_2454);
nor U2579 (N_2579,N_2208,N_2300);
nor U2580 (N_2580,N_2251,N_2435);
or U2581 (N_2581,N_2345,N_2479);
or U2582 (N_2582,N_2252,N_2280);
and U2583 (N_2583,N_2080,N_2012);
nand U2584 (N_2584,N_2063,N_2093);
or U2585 (N_2585,N_2266,N_2009);
and U2586 (N_2586,N_2257,N_2166);
or U2587 (N_2587,N_2428,N_2296);
and U2588 (N_2588,N_2199,N_2218);
and U2589 (N_2589,N_2374,N_2457);
or U2590 (N_2590,N_2360,N_2355);
and U2591 (N_2591,N_2417,N_2301);
or U2592 (N_2592,N_2164,N_2034);
nor U2593 (N_2593,N_2382,N_2110);
nand U2594 (N_2594,N_2108,N_2035);
nor U2595 (N_2595,N_2361,N_2215);
and U2596 (N_2596,N_2383,N_2350);
or U2597 (N_2597,N_2230,N_2372);
and U2598 (N_2598,N_2440,N_2450);
and U2599 (N_2599,N_2118,N_2020);
and U2600 (N_2600,N_2111,N_2107);
nor U2601 (N_2601,N_2265,N_2391);
or U2602 (N_2602,N_2198,N_2352);
nand U2603 (N_2603,N_2276,N_2392);
nor U2604 (N_2604,N_2200,N_2467);
nor U2605 (N_2605,N_2472,N_2309);
and U2606 (N_2606,N_2323,N_2441);
nand U2607 (N_2607,N_2160,N_2263);
and U2608 (N_2608,N_2498,N_2103);
or U2609 (N_2609,N_2216,N_2404);
and U2610 (N_2610,N_2481,N_2119);
or U2611 (N_2611,N_2366,N_2330);
nand U2612 (N_2612,N_2217,N_2375);
or U2613 (N_2613,N_2088,N_2086);
nand U2614 (N_2614,N_2273,N_2097);
nor U2615 (N_2615,N_2016,N_2123);
or U2616 (N_2616,N_2277,N_2286);
or U2617 (N_2617,N_2475,N_2112);
nand U2618 (N_2618,N_2332,N_2135);
or U2619 (N_2619,N_2429,N_2349);
or U2620 (N_2620,N_2004,N_2303);
or U2621 (N_2621,N_2144,N_2168);
nor U2622 (N_2622,N_2101,N_2412);
and U2623 (N_2623,N_2462,N_2302);
or U2624 (N_2624,N_2370,N_2186);
or U2625 (N_2625,N_2059,N_2023);
nand U2626 (N_2626,N_2433,N_2424);
nor U2627 (N_2627,N_2319,N_2488);
nor U2628 (N_2628,N_2142,N_2126);
and U2629 (N_2629,N_2201,N_2452);
or U2630 (N_2630,N_2459,N_2027);
and U2631 (N_2631,N_2313,N_2121);
nand U2632 (N_2632,N_2493,N_2090);
and U2633 (N_2633,N_2387,N_2278);
nor U2634 (N_2634,N_2211,N_2024);
and U2635 (N_2635,N_2304,N_2369);
and U2636 (N_2636,N_2196,N_2044);
or U2637 (N_2637,N_2084,N_2487);
or U2638 (N_2638,N_2482,N_2174);
nor U2639 (N_2639,N_2436,N_2456);
nand U2640 (N_2640,N_2223,N_2311);
nor U2641 (N_2641,N_2253,N_2492);
nand U2642 (N_2642,N_2353,N_2068);
and U2643 (N_2643,N_2396,N_2026);
nor U2644 (N_2644,N_2124,N_2334);
nor U2645 (N_2645,N_2495,N_2364);
nand U2646 (N_2646,N_2343,N_2499);
nor U2647 (N_2647,N_2439,N_2137);
and U2648 (N_2648,N_2075,N_2202);
or U2649 (N_2649,N_2434,N_2178);
or U2650 (N_2650,N_2095,N_2078);
and U2651 (N_2651,N_2393,N_2037);
and U2652 (N_2652,N_2367,N_2132);
nand U2653 (N_2653,N_2212,N_2005);
or U2654 (N_2654,N_2041,N_2389);
and U2655 (N_2655,N_2072,N_2007);
nor U2656 (N_2656,N_2138,N_2427);
or U2657 (N_2657,N_2244,N_2134);
or U2658 (N_2658,N_2053,N_2231);
or U2659 (N_2659,N_2390,N_2425);
nand U2660 (N_2660,N_2170,N_2458);
and U2661 (N_2661,N_2413,N_2324);
and U2662 (N_2662,N_2163,N_2409);
xor U2663 (N_2663,N_2002,N_2205);
nand U2664 (N_2664,N_2128,N_2306);
nand U2665 (N_2665,N_2219,N_2380);
and U2666 (N_2666,N_2494,N_2150);
and U2667 (N_2667,N_2130,N_2192);
or U2668 (N_2668,N_2207,N_2171);
and U2669 (N_2669,N_2096,N_2288);
nor U2670 (N_2670,N_2255,N_2327);
or U2671 (N_2671,N_2430,N_2408);
or U2672 (N_2672,N_2065,N_2054);
nand U2673 (N_2673,N_2470,N_2120);
nor U2674 (N_2674,N_2314,N_2340);
or U2675 (N_2675,N_2157,N_2191);
and U2676 (N_2676,N_2238,N_2139);
nand U2677 (N_2677,N_2445,N_2052);
or U2678 (N_2678,N_2243,N_2259);
and U2679 (N_2679,N_2039,N_2033);
or U2680 (N_2680,N_2465,N_2287);
nand U2681 (N_2681,N_2105,N_2283);
or U2682 (N_2682,N_2373,N_2267);
and U2683 (N_2683,N_2181,N_2437);
nor U2684 (N_2684,N_2250,N_2146);
nand U2685 (N_2685,N_2401,N_2143);
or U2686 (N_2686,N_2189,N_2279);
nand U2687 (N_2687,N_2386,N_2420);
nand U2688 (N_2688,N_2046,N_2358);
nor U2689 (N_2689,N_2407,N_2464);
and U2690 (N_2690,N_2325,N_2362);
or U2691 (N_2691,N_2228,N_2043);
nor U2692 (N_2692,N_2326,N_2416);
nor U2693 (N_2693,N_2335,N_2081);
nor U2694 (N_2694,N_2225,N_2155);
nor U2695 (N_2695,N_2073,N_2414);
or U2696 (N_2696,N_2104,N_2152);
nand U2697 (N_2697,N_2258,N_2264);
and U2698 (N_2698,N_2008,N_2294);
and U2699 (N_2699,N_2014,N_2066);
or U2700 (N_2700,N_2029,N_2299);
or U2701 (N_2701,N_2320,N_2359);
or U2702 (N_2702,N_2448,N_2298);
or U2703 (N_2703,N_2098,N_2419);
or U2704 (N_2704,N_2149,N_2193);
and U2705 (N_2705,N_2438,N_2194);
nand U2706 (N_2706,N_2153,N_2426);
or U2707 (N_2707,N_2140,N_2069);
and U2708 (N_2708,N_2136,N_2184);
or U2709 (N_2709,N_2094,N_2346);
nor U2710 (N_2710,N_2274,N_2431);
nand U2711 (N_2711,N_2021,N_2087);
or U2712 (N_2712,N_2348,N_2010);
nand U2713 (N_2713,N_2047,N_2176);
nand U2714 (N_2714,N_2227,N_2190);
nand U2715 (N_2715,N_2188,N_2042);
nand U2716 (N_2716,N_2490,N_2203);
or U2717 (N_2717,N_2099,N_2339);
nand U2718 (N_2718,N_2017,N_2249);
nand U2719 (N_2719,N_2000,N_2469);
nor U2720 (N_2720,N_2261,N_2310);
nand U2721 (N_2721,N_2159,N_2308);
or U2722 (N_2722,N_2158,N_2442);
and U2723 (N_2723,N_2354,N_2183);
nor U2724 (N_2724,N_2236,N_2347);
nor U2725 (N_2725,N_2398,N_2006);
nor U2726 (N_2726,N_2388,N_2474);
or U2727 (N_2727,N_2318,N_2091);
nand U2728 (N_2728,N_2113,N_2394);
nor U2729 (N_2729,N_2060,N_2328);
or U2730 (N_2730,N_2477,N_2271);
and U2731 (N_2731,N_2102,N_2165);
and U2732 (N_2732,N_2172,N_2275);
or U2733 (N_2733,N_2057,N_2070);
nand U2734 (N_2734,N_2239,N_2377);
and U2735 (N_2735,N_2262,N_2220);
and U2736 (N_2736,N_2100,N_2451);
nand U2737 (N_2737,N_2229,N_2221);
or U2738 (N_2738,N_2015,N_2480);
and U2739 (N_2739,N_2337,N_2185);
or U2740 (N_2740,N_2085,N_2381);
nand U2741 (N_2741,N_2122,N_2247);
or U2742 (N_2742,N_2496,N_2240);
or U2743 (N_2743,N_2341,N_2356);
nand U2744 (N_2744,N_2256,N_2463);
nor U2745 (N_2745,N_2443,N_2131);
and U2746 (N_2746,N_2281,N_2162);
or U2747 (N_2747,N_2282,N_2242);
and U2748 (N_2748,N_2051,N_2284);
and U2749 (N_2749,N_2109,N_2187);
or U2750 (N_2750,N_2007,N_2305);
nor U2751 (N_2751,N_2282,N_2109);
or U2752 (N_2752,N_2259,N_2367);
nor U2753 (N_2753,N_2230,N_2286);
nor U2754 (N_2754,N_2167,N_2238);
nor U2755 (N_2755,N_2052,N_2399);
nand U2756 (N_2756,N_2444,N_2252);
and U2757 (N_2757,N_2381,N_2145);
and U2758 (N_2758,N_2292,N_2400);
or U2759 (N_2759,N_2075,N_2056);
or U2760 (N_2760,N_2333,N_2218);
nor U2761 (N_2761,N_2188,N_2157);
nor U2762 (N_2762,N_2421,N_2191);
nor U2763 (N_2763,N_2465,N_2436);
nor U2764 (N_2764,N_2089,N_2362);
or U2765 (N_2765,N_2223,N_2398);
and U2766 (N_2766,N_2240,N_2447);
nand U2767 (N_2767,N_2247,N_2350);
nand U2768 (N_2768,N_2303,N_2274);
or U2769 (N_2769,N_2013,N_2368);
or U2770 (N_2770,N_2499,N_2356);
or U2771 (N_2771,N_2480,N_2166);
and U2772 (N_2772,N_2232,N_2492);
and U2773 (N_2773,N_2405,N_2460);
nor U2774 (N_2774,N_2306,N_2400);
and U2775 (N_2775,N_2419,N_2178);
or U2776 (N_2776,N_2150,N_2222);
and U2777 (N_2777,N_2464,N_2454);
nor U2778 (N_2778,N_2047,N_2239);
nor U2779 (N_2779,N_2420,N_2388);
or U2780 (N_2780,N_2121,N_2449);
or U2781 (N_2781,N_2374,N_2062);
nor U2782 (N_2782,N_2010,N_2340);
or U2783 (N_2783,N_2460,N_2421);
and U2784 (N_2784,N_2029,N_2039);
nand U2785 (N_2785,N_2273,N_2150);
nor U2786 (N_2786,N_2333,N_2154);
or U2787 (N_2787,N_2034,N_2160);
or U2788 (N_2788,N_2373,N_2353);
or U2789 (N_2789,N_2046,N_2148);
nand U2790 (N_2790,N_2360,N_2037);
nand U2791 (N_2791,N_2221,N_2120);
or U2792 (N_2792,N_2327,N_2221);
nand U2793 (N_2793,N_2335,N_2438);
or U2794 (N_2794,N_2044,N_2212);
nand U2795 (N_2795,N_2247,N_2129);
xor U2796 (N_2796,N_2017,N_2336);
nor U2797 (N_2797,N_2161,N_2234);
or U2798 (N_2798,N_2091,N_2031);
nor U2799 (N_2799,N_2158,N_2421);
nor U2800 (N_2800,N_2193,N_2136);
nor U2801 (N_2801,N_2276,N_2053);
nand U2802 (N_2802,N_2327,N_2257);
nand U2803 (N_2803,N_2282,N_2297);
and U2804 (N_2804,N_2291,N_2462);
and U2805 (N_2805,N_2164,N_2084);
nand U2806 (N_2806,N_2039,N_2167);
or U2807 (N_2807,N_2433,N_2015);
and U2808 (N_2808,N_2375,N_2000);
nor U2809 (N_2809,N_2087,N_2445);
or U2810 (N_2810,N_2030,N_2104);
nor U2811 (N_2811,N_2443,N_2496);
nand U2812 (N_2812,N_2485,N_2127);
nand U2813 (N_2813,N_2289,N_2414);
and U2814 (N_2814,N_2021,N_2389);
nor U2815 (N_2815,N_2350,N_2038);
nand U2816 (N_2816,N_2466,N_2233);
nor U2817 (N_2817,N_2051,N_2336);
nand U2818 (N_2818,N_2092,N_2371);
or U2819 (N_2819,N_2110,N_2405);
or U2820 (N_2820,N_2436,N_2178);
or U2821 (N_2821,N_2061,N_2426);
and U2822 (N_2822,N_2465,N_2498);
nand U2823 (N_2823,N_2113,N_2125);
or U2824 (N_2824,N_2035,N_2066);
and U2825 (N_2825,N_2332,N_2007);
nand U2826 (N_2826,N_2155,N_2404);
nor U2827 (N_2827,N_2370,N_2170);
nor U2828 (N_2828,N_2135,N_2247);
nand U2829 (N_2829,N_2143,N_2166);
or U2830 (N_2830,N_2167,N_2324);
nand U2831 (N_2831,N_2495,N_2444);
nor U2832 (N_2832,N_2150,N_2428);
nand U2833 (N_2833,N_2273,N_2023);
nand U2834 (N_2834,N_2089,N_2387);
nand U2835 (N_2835,N_2286,N_2260);
nor U2836 (N_2836,N_2035,N_2276);
or U2837 (N_2837,N_2071,N_2474);
or U2838 (N_2838,N_2196,N_2144);
nand U2839 (N_2839,N_2044,N_2320);
and U2840 (N_2840,N_2252,N_2340);
nor U2841 (N_2841,N_2462,N_2229);
or U2842 (N_2842,N_2134,N_2227);
nor U2843 (N_2843,N_2379,N_2030);
and U2844 (N_2844,N_2060,N_2435);
or U2845 (N_2845,N_2177,N_2073);
nand U2846 (N_2846,N_2013,N_2180);
nand U2847 (N_2847,N_2168,N_2157);
nor U2848 (N_2848,N_2069,N_2494);
nand U2849 (N_2849,N_2427,N_2271);
nand U2850 (N_2850,N_2369,N_2179);
or U2851 (N_2851,N_2076,N_2392);
nor U2852 (N_2852,N_2401,N_2200);
xor U2853 (N_2853,N_2247,N_2353);
and U2854 (N_2854,N_2124,N_2259);
or U2855 (N_2855,N_2014,N_2272);
or U2856 (N_2856,N_2473,N_2469);
nand U2857 (N_2857,N_2373,N_2366);
nor U2858 (N_2858,N_2245,N_2374);
nand U2859 (N_2859,N_2200,N_2313);
nor U2860 (N_2860,N_2054,N_2008);
nand U2861 (N_2861,N_2300,N_2083);
and U2862 (N_2862,N_2325,N_2205);
or U2863 (N_2863,N_2229,N_2364);
nand U2864 (N_2864,N_2254,N_2368);
and U2865 (N_2865,N_2393,N_2317);
nor U2866 (N_2866,N_2310,N_2431);
nand U2867 (N_2867,N_2394,N_2124);
nand U2868 (N_2868,N_2238,N_2043);
or U2869 (N_2869,N_2016,N_2488);
and U2870 (N_2870,N_2378,N_2018);
or U2871 (N_2871,N_2201,N_2211);
nor U2872 (N_2872,N_2221,N_2415);
and U2873 (N_2873,N_2330,N_2301);
and U2874 (N_2874,N_2129,N_2371);
or U2875 (N_2875,N_2425,N_2319);
and U2876 (N_2876,N_2113,N_2396);
and U2877 (N_2877,N_2274,N_2204);
nor U2878 (N_2878,N_2490,N_2307);
or U2879 (N_2879,N_2182,N_2351);
nor U2880 (N_2880,N_2224,N_2185);
or U2881 (N_2881,N_2330,N_2295);
nand U2882 (N_2882,N_2029,N_2347);
nor U2883 (N_2883,N_2408,N_2342);
and U2884 (N_2884,N_2032,N_2030);
and U2885 (N_2885,N_2108,N_2470);
and U2886 (N_2886,N_2045,N_2314);
nor U2887 (N_2887,N_2282,N_2201);
nand U2888 (N_2888,N_2209,N_2318);
or U2889 (N_2889,N_2114,N_2221);
nand U2890 (N_2890,N_2456,N_2194);
nand U2891 (N_2891,N_2282,N_2262);
nor U2892 (N_2892,N_2240,N_2330);
nand U2893 (N_2893,N_2482,N_2009);
and U2894 (N_2894,N_2363,N_2338);
nand U2895 (N_2895,N_2331,N_2088);
nand U2896 (N_2896,N_2053,N_2017);
nand U2897 (N_2897,N_2013,N_2340);
or U2898 (N_2898,N_2237,N_2257);
or U2899 (N_2899,N_2360,N_2191);
nor U2900 (N_2900,N_2208,N_2135);
or U2901 (N_2901,N_2221,N_2312);
nor U2902 (N_2902,N_2400,N_2457);
nand U2903 (N_2903,N_2359,N_2214);
nand U2904 (N_2904,N_2498,N_2022);
and U2905 (N_2905,N_2385,N_2005);
nand U2906 (N_2906,N_2255,N_2316);
xnor U2907 (N_2907,N_2349,N_2428);
nand U2908 (N_2908,N_2336,N_2386);
and U2909 (N_2909,N_2347,N_2329);
nor U2910 (N_2910,N_2407,N_2450);
nor U2911 (N_2911,N_2127,N_2495);
and U2912 (N_2912,N_2282,N_2026);
or U2913 (N_2913,N_2093,N_2474);
or U2914 (N_2914,N_2121,N_2242);
nand U2915 (N_2915,N_2153,N_2036);
or U2916 (N_2916,N_2341,N_2218);
or U2917 (N_2917,N_2329,N_2237);
and U2918 (N_2918,N_2462,N_2030);
nand U2919 (N_2919,N_2467,N_2258);
nand U2920 (N_2920,N_2238,N_2354);
and U2921 (N_2921,N_2012,N_2303);
nor U2922 (N_2922,N_2293,N_2352);
and U2923 (N_2923,N_2099,N_2361);
nor U2924 (N_2924,N_2361,N_2369);
nand U2925 (N_2925,N_2240,N_2181);
nor U2926 (N_2926,N_2406,N_2059);
nor U2927 (N_2927,N_2404,N_2147);
or U2928 (N_2928,N_2414,N_2227);
nand U2929 (N_2929,N_2104,N_2240);
or U2930 (N_2930,N_2085,N_2019);
nand U2931 (N_2931,N_2374,N_2070);
nor U2932 (N_2932,N_2098,N_2183);
nor U2933 (N_2933,N_2087,N_2487);
or U2934 (N_2934,N_2461,N_2002);
nand U2935 (N_2935,N_2486,N_2016);
nand U2936 (N_2936,N_2464,N_2479);
nand U2937 (N_2937,N_2040,N_2489);
or U2938 (N_2938,N_2029,N_2307);
nor U2939 (N_2939,N_2411,N_2478);
nand U2940 (N_2940,N_2044,N_2006);
nand U2941 (N_2941,N_2445,N_2150);
or U2942 (N_2942,N_2197,N_2161);
nand U2943 (N_2943,N_2492,N_2303);
and U2944 (N_2944,N_2317,N_2122);
or U2945 (N_2945,N_2123,N_2359);
nor U2946 (N_2946,N_2460,N_2499);
and U2947 (N_2947,N_2098,N_2107);
or U2948 (N_2948,N_2306,N_2152);
or U2949 (N_2949,N_2392,N_2320);
and U2950 (N_2950,N_2148,N_2196);
or U2951 (N_2951,N_2249,N_2294);
nand U2952 (N_2952,N_2317,N_2481);
and U2953 (N_2953,N_2318,N_2172);
nand U2954 (N_2954,N_2034,N_2280);
nor U2955 (N_2955,N_2146,N_2419);
and U2956 (N_2956,N_2463,N_2478);
or U2957 (N_2957,N_2495,N_2137);
nand U2958 (N_2958,N_2285,N_2302);
and U2959 (N_2959,N_2251,N_2087);
or U2960 (N_2960,N_2490,N_2466);
and U2961 (N_2961,N_2488,N_2242);
nor U2962 (N_2962,N_2424,N_2124);
nand U2963 (N_2963,N_2471,N_2410);
nor U2964 (N_2964,N_2216,N_2416);
nor U2965 (N_2965,N_2321,N_2403);
nor U2966 (N_2966,N_2012,N_2389);
and U2967 (N_2967,N_2075,N_2035);
or U2968 (N_2968,N_2344,N_2100);
xor U2969 (N_2969,N_2226,N_2105);
and U2970 (N_2970,N_2362,N_2030);
and U2971 (N_2971,N_2017,N_2418);
and U2972 (N_2972,N_2031,N_2408);
or U2973 (N_2973,N_2058,N_2157);
and U2974 (N_2974,N_2189,N_2164);
nor U2975 (N_2975,N_2408,N_2074);
nor U2976 (N_2976,N_2278,N_2318);
nand U2977 (N_2977,N_2081,N_2179);
nand U2978 (N_2978,N_2496,N_2040);
nand U2979 (N_2979,N_2144,N_2274);
or U2980 (N_2980,N_2487,N_2234);
or U2981 (N_2981,N_2062,N_2161);
and U2982 (N_2982,N_2423,N_2254);
or U2983 (N_2983,N_2482,N_2141);
nand U2984 (N_2984,N_2315,N_2468);
nand U2985 (N_2985,N_2329,N_2140);
nor U2986 (N_2986,N_2460,N_2258);
and U2987 (N_2987,N_2171,N_2365);
or U2988 (N_2988,N_2173,N_2409);
or U2989 (N_2989,N_2317,N_2025);
xnor U2990 (N_2990,N_2318,N_2166);
and U2991 (N_2991,N_2320,N_2434);
and U2992 (N_2992,N_2271,N_2058);
and U2993 (N_2993,N_2404,N_2074);
nor U2994 (N_2994,N_2001,N_2041);
nor U2995 (N_2995,N_2373,N_2073);
nor U2996 (N_2996,N_2463,N_2132);
nand U2997 (N_2997,N_2052,N_2349);
nor U2998 (N_2998,N_2147,N_2406);
nand U2999 (N_2999,N_2281,N_2031);
nor UO_0 (O_0,N_2881,N_2702);
nor UO_1 (O_1,N_2983,N_2990);
nand UO_2 (O_2,N_2855,N_2549);
nand UO_3 (O_3,N_2765,N_2595);
nor UO_4 (O_4,N_2759,N_2762);
and UO_5 (O_5,N_2524,N_2939);
or UO_6 (O_6,N_2701,N_2501);
nor UO_7 (O_7,N_2566,N_2737);
nand UO_8 (O_8,N_2796,N_2628);
nor UO_9 (O_9,N_2603,N_2999);
nor UO_10 (O_10,N_2948,N_2587);
nor UO_11 (O_11,N_2976,N_2538);
and UO_12 (O_12,N_2526,N_2950);
nand UO_13 (O_13,N_2898,N_2882);
or UO_14 (O_14,N_2854,N_2539);
nor UO_15 (O_15,N_2530,N_2716);
or UO_16 (O_16,N_2920,N_2704);
or UO_17 (O_17,N_2916,N_2993);
or UO_18 (O_18,N_2621,N_2975);
and UO_19 (O_19,N_2535,N_2864);
and UO_20 (O_20,N_2632,N_2819);
nor UO_21 (O_21,N_2921,N_2901);
or UO_22 (O_22,N_2778,N_2940);
nand UO_23 (O_23,N_2981,N_2690);
or UO_24 (O_24,N_2693,N_2679);
nand UO_25 (O_25,N_2803,N_2785);
or UO_26 (O_26,N_2805,N_2671);
nand UO_27 (O_27,N_2997,N_2531);
nor UO_28 (O_28,N_2746,N_2744);
and UO_29 (O_29,N_2893,N_2822);
or UO_30 (O_30,N_2637,N_2573);
or UO_31 (O_31,N_2706,N_2946);
or UO_32 (O_32,N_2646,N_2793);
or UO_33 (O_33,N_2982,N_2789);
nand UO_34 (O_34,N_2599,N_2675);
and UO_35 (O_35,N_2517,N_2825);
and UO_36 (O_36,N_2574,N_2771);
and UO_37 (O_37,N_2593,N_2724);
nor UO_38 (O_38,N_2634,N_2899);
nand UO_39 (O_39,N_2735,N_2721);
nand UO_40 (O_40,N_2842,N_2799);
or UO_41 (O_41,N_2583,N_2601);
and UO_42 (O_42,N_2745,N_2533);
nor UO_43 (O_43,N_2908,N_2510);
nor UO_44 (O_44,N_2889,N_2705);
or UO_45 (O_45,N_2584,N_2629);
or UO_46 (O_46,N_2725,N_2534);
and UO_47 (O_47,N_2890,N_2970);
and UO_48 (O_48,N_2585,N_2779);
nand UO_49 (O_49,N_2651,N_2772);
nor UO_50 (O_50,N_2888,N_2840);
nand UO_51 (O_51,N_2977,N_2521);
and UO_52 (O_52,N_2801,N_2857);
xor UO_53 (O_53,N_2775,N_2987);
nor UO_54 (O_54,N_2710,N_2995);
nand UO_55 (O_55,N_2512,N_2734);
or UO_56 (O_56,N_2672,N_2984);
and UO_57 (O_57,N_2794,N_2644);
nand UO_58 (O_58,N_2726,N_2811);
and UO_59 (O_59,N_2918,N_2786);
or UO_60 (O_60,N_2974,N_2572);
nor UO_61 (O_61,N_2795,N_2586);
and UO_62 (O_62,N_2518,N_2618);
or UO_63 (O_63,N_2782,N_2760);
or UO_64 (O_64,N_2508,N_2992);
and UO_65 (O_65,N_2807,N_2766);
and UO_66 (O_66,N_2617,N_2849);
and UO_67 (O_67,N_2653,N_2979);
nor UO_68 (O_68,N_2555,N_2522);
and UO_69 (O_69,N_2597,N_2816);
nand UO_70 (O_70,N_2592,N_2936);
nor UO_71 (O_71,N_2622,N_2541);
or UO_72 (O_72,N_2832,N_2620);
or UO_73 (O_73,N_2625,N_2758);
or UO_74 (O_74,N_2875,N_2770);
and UO_75 (O_75,N_2686,N_2868);
or UO_76 (O_76,N_2509,N_2960);
nor UO_77 (O_77,N_2713,N_2998);
and UO_78 (O_78,N_2626,N_2699);
nand UO_79 (O_79,N_2878,N_2945);
nand UO_80 (O_80,N_2678,N_2841);
nand UO_81 (O_81,N_2742,N_2567);
or UO_82 (O_82,N_2519,N_2876);
nor UO_83 (O_83,N_2767,N_2696);
or UO_84 (O_84,N_2565,N_2663);
or UO_85 (O_85,N_2902,N_2931);
nor UO_86 (O_86,N_2907,N_2588);
or UO_87 (O_87,N_2787,N_2930);
or UO_88 (O_88,N_2718,N_2935);
and UO_89 (O_89,N_2543,N_2667);
nor UO_90 (O_90,N_2577,N_2873);
nor UO_91 (O_91,N_2809,N_2514);
nand UO_92 (O_92,N_2925,N_2648);
nor UO_93 (O_93,N_2738,N_2863);
nand UO_94 (O_94,N_2967,N_2978);
or UO_95 (O_95,N_2523,N_2835);
or UO_96 (O_96,N_2641,N_2631);
or UO_97 (O_97,N_2537,N_2790);
nor UO_98 (O_98,N_2818,N_2972);
or UO_99 (O_99,N_2717,N_2958);
nand UO_100 (O_100,N_2502,N_2886);
and UO_101 (O_101,N_2607,N_2853);
and UO_102 (O_102,N_2828,N_2548);
and UO_103 (O_103,N_2910,N_2783);
and UO_104 (O_104,N_2985,N_2844);
nor UO_105 (O_105,N_2866,N_2688);
nand UO_106 (O_106,N_2837,N_2906);
nand UO_107 (O_107,N_2529,N_2571);
and UO_108 (O_108,N_2552,N_2851);
nor UO_109 (O_109,N_2860,N_2943);
and UO_110 (O_110,N_2895,N_2870);
nand UO_111 (O_111,N_2773,N_2934);
nor UO_112 (O_112,N_2557,N_2569);
or UO_113 (O_113,N_2937,N_2560);
or UO_114 (O_114,N_2674,N_2885);
and UO_115 (O_115,N_2676,N_2989);
and UO_116 (O_116,N_2662,N_2823);
and UO_117 (O_117,N_2961,N_2944);
or UO_118 (O_118,N_2610,N_2558);
nor UO_119 (O_119,N_2732,N_2660);
nand UO_120 (O_120,N_2956,N_2719);
nor UO_121 (O_121,N_2747,N_2954);
and UO_122 (O_122,N_2743,N_2691);
nor UO_123 (O_123,N_2589,N_2904);
nor UO_124 (O_124,N_2761,N_2709);
nor UO_125 (O_125,N_2513,N_2687);
nand UO_126 (O_126,N_2838,N_2915);
or UO_127 (O_127,N_2968,N_2645);
nor UO_128 (O_128,N_2768,N_2612);
nor UO_129 (O_129,N_2623,N_2722);
and UO_130 (O_130,N_2579,N_2568);
nor UO_131 (O_131,N_2856,N_2581);
or UO_132 (O_132,N_2681,N_2695);
nor UO_133 (O_133,N_2707,N_2896);
or UO_134 (O_134,N_2833,N_2959);
or UO_135 (O_135,N_2666,N_2836);
and UO_136 (O_136,N_2536,N_2843);
nand UO_137 (O_137,N_2503,N_2802);
nand UO_138 (O_138,N_2845,N_2880);
and UO_139 (O_139,N_2784,N_2812);
and UO_140 (O_140,N_2909,N_2764);
nor UO_141 (O_141,N_2846,N_2605);
nand UO_142 (O_142,N_2624,N_2955);
nor UO_143 (O_143,N_2847,N_2730);
or UO_144 (O_144,N_2797,N_2578);
and UO_145 (O_145,N_2994,N_2776);
nand UO_146 (O_146,N_2542,N_2963);
and UO_147 (O_147,N_2545,N_2698);
or UO_148 (O_148,N_2570,N_2774);
or UO_149 (O_149,N_2657,N_2996);
nand UO_150 (O_150,N_2810,N_2669);
or UO_151 (O_151,N_2755,N_2532);
nor UO_152 (O_152,N_2665,N_2932);
or UO_153 (O_153,N_2897,N_2913);
or UO_154 (O_154,N_2938,N_2600);
or UO_155 (O_155,N_2576,N_2694);
or UO_156 (O_156,N_2551,N_2563);
nand UO_157 (O_157,N_2727,N_2941);
xnor UO_158 (O_158,N_2928,N_2650);
or UO_159 (O_159,N_2692,N_2652);
nor UO_160 (O_160,N_2731,N_2824);
or UO_161 (O_161,N_2630,N_2988);
or UO_162 (O_162,N_2594,N_2712);
nand UO_163 (O_163,N_2554,N_2754);
nand UO_164 (O_164,N_2639,N_2613);
nand UO_165 (O_165,N_2608,N_2606);
or UO_166 (O_166,N_2750,N_2830);
or UO_167 (O_167,N_2872,N_2962);
or UO_168 (O_168,N_2813,N_2611);
nand UO_169 (O_169,N_2942,N_2867);
nor UO_170 (O_170,N_2923,N_2527);
and UO_171 (O_171,N_2991,N_2804);
nand UO_172 (O_172,N_2839,N_2850);
or UO_173 (O_173,N_2800,N_2520);
and UO_174 (O_174,N_2553,N_2861);
nand UO_175 (O_175,N_2929,N_2602);
or UO_176 (O_176,N_2505,N_2753);
or UO_177 (O_177,N_2966,N_2643);
or UO_178 (O_178,N_2964,N_2635);
and UO_179 (O_179,N_2757,N_2673);
or UO_180 (O_180,N_2798,N_2740);
and UO_181 (O_181,N_2777,N_2654);
and UO_182 (O_182,N_2806,N_2682);
nor UO_183 (O_183,N_2865,N_2728);
nand UO_184 (O_184,N_2905,N_2769);
and UO_185 (O_185,N_2927,N_2661);
nor UO_186 (O_186,N_2763,N_2922);
and UO_187 (O_187,N_2969,N_2792);
nor UO_188 (O_188,N_2658,N_2751);
nand UO_189 (O_189,N_2525,N_2820);
or UO_190 (O_190,N_2596,N_2914);
nand UO_191 (O_191,N_2604,N_2649);
or UO_192 (O_192,N_2700,N_2703);
nor UO_193 (O_193,N_2924,N_2590);
nor UO_194 (O_194,N_2831,N_2808);
and UO_195 (O_195,N_2874,N_2827);
and UO_196 (O_196,N_2511,N_2619);
and UO_197 (O_197,N_2507,N_2957);
xnor UO_198 (O_198,N_2684,N_2729);
nand UO_199 (O_199,N_2642,N_2965);
nor UO_200 (O_200,N_2500,N_2791);
xnor UO_201 (O_201,N_2756,N_2616);
nand UO_202 (O_202,N_2677,N_2561);
or UO_203 (O_203,N_2980,N_2598);
and UO_204 (O_204,N_2638,N_2656);
nand UO_205 (O_205,N_2550,N_2711);
nand UO_206 (O_206,N_2826,N_2556);
nor UO_207 (O_207,N_2564,N_2953);
nor UO_208 (O_208,N_2670,N_2871);
and UO_209 (O_209,N_2540,N_2951);
and UO_210 (O_210,N_2926,N_2919);
and UO_211 (O_211,N_2852,N_2894);
or UO_212 (O_212,N_2971,N_2834);
and UO_213 (O_213,N_2933,N_2917);
or UO_214 (O_214,N_2614,N_2715);
or UO_215 (O_215,N_2515,N_2859);
nand UO_216 (O_216,N_2633,N_2697);
or UO_217 (O_217,N_2862,N_2733);
and UO_218 (O_218,N_2903,N_2683);
nand UO_219 (O_219,N_2748,N_2640);
or UO_220 (O_220,N_2952,N_2575);
nor UO_221 (O_221,N_2720,N_2506);
and UO_222 (O_222,N_2814,N_2562);
and UO_223 (O_223,N_2591,N_2869);
or UO_224 (O_224,N_2883,N_2528);
nor UO_225 (O_225,N_2636,N_2516);
nand UO_226 (O_226,N_2664,N_2609);
and UO_227 (O_227,N_2736,N_2547);
nand UO_228 (O_228,N_2815,N_2973);
nor UO_229 (O_229,N_2685,N_2689);
nor UO_230 (O_230,N_2559,N_2668);
and UO_231 (O_231,N_2627,N_2504);
or UO_232 (O_232,N_2680,N_2817);
or UO_233 (O_233,N_2912,N_2821);
or UO_234 (O_234,N_2848,N_2781);
and UO_235 (O_235,N_2887,N_2580);
nand UO_236 (O_236,N_2947,N_2723);
nor UO_237 (O_237,N_2655,N_2752);
and UO_238 (O_238,N_2892,N_2780);
and UO_239 (O_239,N_2708,N_2911);
or UO_240 (O_240,N_2647,N_2829);
nor UO_241 (O_241,N_2546,N_2891);
or UO_242 (O_242,N_2949,N_2739);
and UO_243 (O_243,N_2544,N_2858);
nor UO_244 (O_244,N_2749,N_2884);
nand UO_245 (O_245,N_2877,N_2879);
nand UO_246 (O_246,N_2900,N_2615);
nand UO_247 (O_247,N_2986,N_2714);
nand UO_248 (O_248,N_2659,N_2582);
or UO_249 (O_249,N_2741,N_2788);
and UO_250 (O_250,N_2614,N_2967);
and UO_251 (O_251,N_2961,N_2922);
nor UO_252 (O_252,N_2764,N_2802);
nand UO_253 (O_253,N_2610,N_2847);
or UO_254 (O_254,N_2505,N_2664);
nand UO_255 (O_255,N_2509,N_2562);
or UO_256 (O_256,N_2627,N_2626);
nand UO_257 (O_257,N_2697,N_2833);
nor UO_258 (O_258,N_2652,N_2860);
nor UO_259 (O_259,N_2718,N_2511);
and UO_260 (O_260,N_2605,N_2956);
and UO_261 (O_261,N_2634,N_2901);
nand UO_262 (O_262,N_2940,N_2586);
and UO_263 (O_263,N_2613,N_2523);
nand UO_264 (O_264,N_2971,N_2535);
or UO_265 (O_265,N_2674,N_2799);
or UO_266 (O_266,N_2526,N_2535);
nand UO_267 (O_267,N_2533,N_2992);
or UO_268 (O_268,N_2799,N_2902);
or UO_269 (O_269,N_2855,N_2744);
or UO_270 (O_270,N_2954,N_2990);
and UO_271 (O_271,N_2757,N_2827);
nor UO_272 (O_272,N_2836,N_2533);
or UO_273 (O_273,N_2778,N_2751);
or UO_274 (O_274,N_2995,N_2969);
nand UO_275 (O_275,N_2651,N_2559);
or UO_276 (O_276,N_2651,N_2702);
nand UO_277 (O_277,N_2689,N_2927);
or UO_278 (O_278,N_2611,N_2844);
nand UO_279 (O_279,N_2957,N_2877);
or UO_280 (O_280,N_2973,N_2616);
nor UO_281 (O_281,N_2684,N_2835);
nor UO_282 (O_282,N_2769,N_2953);
or UO_283 (O_283,N_2513,N_2551);
nand UO_284 (O_284,N_2784,N_2877);
nand UO_285 (O_285,N_2676,N_2720);
nand UO_286 (O_286,N_2703,N_2778);
or UO_287 (O_287,N_2629,N_2915);
or UO_288 (O_288,N_2699,N_2753);
or UO_289 (O_289,N_2800,N_2570);
or UO_290 (O_290,N_2629,N_2932);
nor UO_291 (O_291,N_2775,N_2900);
nand UO_292 (O_292,N_2630,N_2724);
and UO_293 (O_293,N_2640,N_2912);
and UO_294 (O_294,N_2847,N_2574);
and UO_295 (O_295,N_2822,N_2734);
nand UO_296 (O_296,N_2782,N_2776);
and UO_297 (O_297,N_2990,N_2669);
nand UO_298 (O_298,N_2694,N_2711);
or UO_299 (O_299,N_2575,N_2671);
nand UO_300 (O_300,N_2608,N_2779);
or UO_301 (O_301,N_2727,N_2691);
nor UO_302 (O_302,N_2818,N_2635);
nor UO_303 (O_303,N_2781,N_2906);
and UO_304 (O_304,N_2763,N_2748);
nor UO_305 (O_305,N_2798,N_2632);
nand UO_306 (O_306,N_2519,N_2996);
nand UO_307 (O_307,N_2671,N_2500);
or UO_308 (O_308,N_2665,N_2887);
or UO_309 (O_309,N_2559,N_2689);
nor UO_310 (O_310,N_2627,N_2940);
or UO_311 (O_311,N_2904,N_2881);
or UO_312 (O_312,N_2753,N_2599);
and UO_313 (O_313,N_2714,N_2779);
and UO_314 (O_314,N_2518,N_2886);
nand UO_315 (O_315,N_2701,N_2816);
or UO_316 (O_316,N_2651,N_2913);
nand UO_317 (O_317,N_2581,N_2693);
nand UO_318 (O_318,N_2937,N_2763);
and UO_319 (O_319,N_2797,N_2717);
and UO_320 (O_320,N_2870,N_2657);
or UO_321 (O_321,N_2959,N_2633);
nand UO_322 (O_322,N_2993,N_2755);
or UO_323 (O_323,N_2884,N_2736);
and UO_324 (O_324,N_2779,N_2962);
nand UO_325 (O_325,N_2647,N_2859);
nor UO_326 (O_326,N_2601,N_2520);
or UO_327 (O_327,N_2605,N_2571);
nand UO_328 (O_328,N_2762,N_2689);
nand UO_329 (O_329,N_2976,N_2796);
and UO_330 (O_330,N_2893,N_2973);
nand UO_331 (O_331,N_2706,N_2745);
xor UO_332 (O_332,N_2705,N_2596);
nand UO_333 (O_333,N_2904,N_2832);
nor UO_334 (O_334,N_2537,N_2905);
nand UO_335 (O_335,N_2781,N_2888);
nand UO_336 (O_336,N_2700,N_2603);
or UO_337 (O_337,N_2636,N_2845);
or UO_338 (O_338,N_2958,N_2951);
or UO_339 (O_339,N_2906,N_2796);
xnor UO_340 (O_340,N_2555,N_2707);
or UO_341 (O_341,N_2853,N_2504);
xor UO_342 (O_342,N_2617,N_2520);
or UO_343 (O_343,N_2591,N_2501);
or UO_344 (O_344,N_2850,N_2970);
and UO_345 (O_345,N_2869,N_2719);
nand UO_346 (O_346,N_2937,N_2967);
or UO_347 (O_347,N_2835,N_2677);
nand UO_348 (O_348,N_2911,N_2523);
or UO_349 (O_349,N_2921,N_2523);
and UO_350 (O_350,N_2733,N_2855);
or UO_351 (O_351,N_2737,N_2676);
or UO_352 (O_352,N_2864,N_2625);
nor UO_353 (O_353,N_2989,N_2589);
nor UO_354 (O_354,N_2593,N_2776);
or UO_355 (O_355,N_2996,N_2686);
nor UO_356 (O_356,N_2891,N_2904);
and UO_357 (O_357,N_2858,N_2961);
nor UO_358 (O_358,N_2742,N_2730);
nand UO_359 (O_359,N_2836,N_2638);
nor UO_360 (O_360,N_2719,N_2739);
nor UO_361 (O_361,N_2904,N_2500);
and UO_362 (O_362,N_2801,N_2559);
and UO_363 (O_363,N_2732,N_2601);
nor UO_364 (O_364,N_2639,N_2813);
or UO_365 (O_365,N_2711,N_2825);
nand UO_366 (O_366,N_2763,N_2838);
nor UO_367 (O_367,N_2778,N_2732);
or UO_368 (O_368,N_2714,N_2902);
or UO_369 (O_369,N_2789,N_2934);
or UO_370 (O_370,N_2713,N_2749);
and UO_371 (O_371,N_2504,N_2655);
nor UO_372 (O_372,N_2886,N_2737);
nor UO_373 (O_373,N_2678,N_2607);
nor UO_374 (O_374,N_2574,N_2742);
nor UO_375 (O_375,N_2540,N_2530);
nand UO_376 (O_376,N_2741,N_2841);
or UO_377 (O_377,N_2630,N_2606);
nand UO_378 (O_378,N_2954,N_2559);
nand UO_379 (O_379,N_2541,N_2878);
and UO_380 (O_380,N_2739,N_2827);
nand UO_381 (O_381,N_2833,N_2971);
or UO_382 (O_382,N_2814,N_2594);
or UO_383 (O_383,N_2704,N_2669);
or UO_384 (O_384,N_2714,N_2649);
nand UO_385 (O_385,N_2560,N_2960);
nor UO_386 (O_386,N_2953,N_2963);
and UO_387 (O_387,N_2679,N_2956);
nor UO_388 (O_388,N_2513,N_2658);
nand UO_389 (O_389,N_2943,N_2883);
or UO_390 (O_390,N_2588,N_2500);
and UO_391 (O_391,N_2565,N_2725);
nand UO_392 (O_392,N_2751,N_2669);
or UO_393 (O_393,N_2780,N_2658);
and UO_394 (O_394,N_2721,N_2945);
nor UO_395 (O_395,N_2629,N_2959);
and UO_396 (O_396,N_2905,N_2666);
or UO_397 (O_397,N_2573,N_2628);
nand UO_398 (O_398,N_2644,N_2695);
nor UO_399 (O_399,N_2792,N_2695);
nand UO_400 (O_400,N_2972,N_2668);
nand UO_401 (O_401,N_2848,N_2994);
nand UO_402 (O_402,N_2827,N_2882);
nor UO_403 (O_403,N_2599,N_2987);
nor UO_404 (O_404,N_2542,N_2808);
nor UO_405 (O_405,N_2824,N_2727);
nor UO_406 (O_406,N_2637,N_2812);
or UO_407 (O_407,N_2858,N_2621);
nand UO_408 (O_408,N_2721,N_2715);
and UO_409 (O_409,N_2831,N_2693);
nand UO_410 (O_410,N_2752,N_2595);
nand UO_411 (O_411,N_2780,N_2987);
or UO_412 (O_412,N_2580,N_2504);
nor UO_413 (O_413,N_2594,N_2976);
nor UO_414 (O_414,N_2573,N_2769);
nand UO_415 (O_415,N_2693,N_2612);
nor UO_416 (O_416,N_2573,N_2874);
or UO_417 (O_417,N_2777,N_2585);
nor UO_418 (O_418,N_2642,N_2684);
and UO_419 (O_419,N_2604,N_2693);
nand UO_420 (O_420,N_2877,N_2641);
nand UO_421 (O_421,N_2688,N_2872);
nor UO_422 (O_422,N_2717,N_2738);
nor UO_423 (O_423,N_2633,N_2917);
nand UO_424 (O_424,N_2712,N_2932);
or UO_425 (O_425,N_2968,N_2558);
nand UO_426 (O_426,N_2731,N_2701);
nor UO_427 (O_427,N_2727,N_2515);
nand UO_428 (O_428,N_2779,N_2507);
or UO_429 (O_429,N_2511,N_2539);
and UO_430 (O_430,N_2908,N_2780);
and UO_431 (O_431,N_2551,N_2853);
and UO_432 (O_432,N_2953,N_2531);
nor UO_433 (O_433,N_2869,N_2938);
nand UO_434 (O_434,N_2659,N_2559);
or UO_435 (O_435,N_2527,N_2820);
nor UO_436 (O_436,N_2941,N_2731);
or UO_437 (O_437,N_2833,N_2916);
and UO_438 (O_438,N_2850,N_2964);
or UO_439 (O_439,N_2637,N_2932);
nand UO_440 (O_440,N_2794,N_2934);
and UO_441 (O_441,N_2984,N_2658);
nor UO_442 (O_442,N_2863,N_2909);
nor UO_443 (O_443,N_2846,N_2740);
or UO_444 (O_444,N_2968,N_2651);
and UO_445 (O_445,N_2627,N_2909);
nor UO_446 (O_446,N_2729,N_2981);
nand UO_447 (O_447,N_2786,N_2602);
nand UO_448 (O_448,N_2504,N_2503);
nor UO_449 (O_449,N_2841,N_2773);
nor UO_450 (O_450,N_2605,N_2584);
and UO_451 (O_451,N_2581,N_2977);
and UO_452 (O_452,N_2779,N_2737);
or UO_453 (O_453,N_2611,N_2826);
and UO_454 (O_454,N_2852,N_2733);
or UO_455 (O_455,N_2581,N_2880);
or UO_456 (O_456,N_2759,N_2855);
or UO_457 (O_457,N_2569,N_2769);
nor UO_458 (O_458,N_2594,N_2836);
nand UO_459 (O_459,N_2935,N_2864);
or UO_460 (O_460,N_2827,N_2919);
or UO_461 (O_461,N_2646,N_2989);
or UO_462 (O_462,N_2608,N_2884);
nor UO_463 (O_463,N_2755,N_2527);
nand UO_464 (O_464,N_2691,N_2828);
nor UO_465 (O_465,N_2633,N_2549);
and UO_466 (O_466,N_2808,N_2590);
nor UO_467 (O_467,N_2840,N_2639);
nand UO_468 (O_468,N_2557,N_2799);
or UO_469 (O_469,N_2838,N_2916);
nor UO_470 (O_470,N_2681,N_2835);
nand UO_471 (O_471,N_2796,N_2570);
or UO_472 (O_472,N_2975,N_2817);
nor UO_473 (O_473,N_2885,N_2590);
nor UO_474 (O_474,N_2956,N_2798);
nand UO_475 (O_475,N_2845,N_2673);
and UO_476 (O_476,N_2866,N_2620);
or UO_477 (O_477,N_2771,N_2693);
nand UO_478 (O_478,N_2621,N_2532);
or UO_479 (O_479,N_2725,N_2531);
nand UO_480 (O_480,N_2665,N_2626);
and UO_481 (O_481,N_2607,N_2791);
nor UO_482 (O_482,N_2841,N_2932);
and UO_483 (O_483,N_2515,N_2894);
and UO_484 (O_484,N_2813,N_2670);
nand UO_485 (O_485,N_2768,N_2933);
nand UO_486 (O_486,N_2751,N_2580);
and UO_487 (O_487,N_2966,N_2844);
nand UO_488 (O_488,N_2744,N_2726);
nand UO_489 (O_489,N_2710,N_2821);
nor UO_490 (O_490,N_2858,N_2586);
nand UO_491 (O_491,N_2993,N_2801);
or UO_492 (O_492,N_2544,N_2869);
xnor UO_493 (O_493,N_2500,N_2621);
nor UO_494 (O_494,N_2878,N_2509);
or UO_495 (O_495,N_2658,N_2849);
nand UO_496 (O_496,N_2857,N_2779);
nand UO_497 (O_497,N_2907,N_2626);
and UO_498 (O_498,N_2767,N_2563);
or UO_499 (O_499,N_2520,N_2885);
endmodule