module basic_500_3000_500_15_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_475,In_459);
or U1 (N_1,In_126,In_381);
xor U2 (N_2,In_227,In_272);
xor U3 (N_3,In_34,In_450);
nor U4 (N_4,In_442,In_104);
xnor U5 (N_5,In_81,In_330);
xnor U6 (N_6,In_476,In_41);
or U7 (N_7,In_491,In_148);
nand U8 (N_8,In_301,In_370);
xnor U9 (N_9,In_343,In_128);
xnor U10 (N_10,In_277,In_36);
nor U11 (N_11,In_218,In_294);
or U12 (N_12,In_235,In_7);
or U13 (N_13,In_44,In_72);
and U14 (N_14,In_27,In_319);
nand U15 (N_15,In_152,In_295);
nor U16 (N_16,In_496,In_140);
xor U17 (N_17,In_264,In_14);
or U18 (N_18,In_422,In_324);
nand U19 (N_19,In_130,In_401);
nor U20 (N_20,In_125,In_311);
or U21 (N_21,In_177,In_349);
and U22 (N_22,In_68,In_179);
nand U23 (N_23,In_413,In_67);
and U24 (N_24,In_409,In_304);
or U25 (N_25,In_172,In_8);
or U26 (N_26,In_99,In_223);
xor U27 (N_27,In_63,In_320);
or U28 (N_28,In_468,In_121);
nand U29 (N_29,In_166,In_392);
or U30 (N_30,In_372,In_191);
nor U31 (N_31,In_342,In_169);
xnor U32 (N_32,In_79,In_228);
or U33 (N_33,In_13,In_131);
xor U34 (N_34,In_215,In_415);
xor U35 (N_35,In_245,In_209);
nor U36 (N_36,In_205,In_335);
nand U37 (N_37,In_302,In_113);
nor U38 (N_38,In_388,In_90);
and U39 (N_39,In_73,In_426);
or U40 (N_40,In_135,In_280);
xor U41 (N_41,In_256,In_32);
nand U42 (N_42,In_486,In_250);
nor U43 (N_43,In_16,In_400);
nor U44 (N_44,In_282,In_395);
xor U45 (N_45,In_274,In_3);
xnor U46 (N_46,In_178,In_208);
or U47 (N_47,In_407,In_481);
nor U48 (N_48,In_203,In_193);
nand U49 (N_49,In_144,In_421);
or U50 (N_50,In_216,In_50);
nor U51 (N_51,In_168,In_346);
nand U52 (N_52,In_240,In_487);
and U53 (N_53,In_490,In_150);
nor U54 (N_54,In_316,In_229);
nand U55 (N_55,In_305,In_397);
nand U56 (N_56,In_202,In_437);
xnor U57 (N_57,In_290,In_380);
xnor U58 (N_58,In_431,In_165);
nor U59 (N_59,In_410,In_232);
nor U60 (N_60,In_428,In_321);
or U61 (N_61,In_173,In_97);
nand U62 (N_62,In_315,In_260);
and U63 (N_63,In_281,In_136);
and U64 (N_64,In_341,In_45);
nor U65 (N_65,In_248,In_257);
nand U66 (N_66,In_84,In_484);
nor U67 (N_67,In_350,In_347);
and U68 (N_68,In_270,In_275);
or U69 (N_69,In_210,In_78);
nor U70 (N_70,In_58,In_112);
nand U71 (N_71,In_391,In_389);
or U72 (N_72,In_93,In_366);
and U73 (N_73,In_473,In_263);
xnor U74 (N_74,In_306,In_207);
nand U75 (N_75,In_153,In_106);
nand U76 (N_76,In_190,In_92);
and U77 (N_77,In_226,In_19);
nor U78 (N_78,In_379,In_2);
and U79 (N_79,In_384,In_181);
or U80 (N_80,In_162,In_157);
or U81 (N_81,In_31,In_292);
nor U82 (N_82,In_364,In_35);
xnor U83 (N_83,In_20,In_189);
xor U84 (N_84,In_246,In_103);
nor U85 (N_85,In_489,In_60);
or U86 (N_86,In_465,In_488);
nor U87 (N_87,In_377,In_262);
nand U88 (N_88,In_253,In_495);
or U89 (N_89,In_61,In_77);
nor U90 (N_90,In_435,In_17);
and U91 (N_91,In_474,In_98);
or U92 (N_92,In_333,In_182);
or U93 (N_93,In_382,In_398);
and U94 (N_94,In_278,In_239);
and U95 (N_95,In_116,In_322);
xnor U96 (N_96,In_361,In_463);
or U97 (N_97,In_441,In_149);
nand U98 (N_98,In_18,In_214);
or U99 (N_99,In_477,In_86);
nand U100 (N_100,In_309,In_143);
nand U101 (N_101,In_11,In_254);
xnor U102 (N_102,In_9,In_453);
nor U103 (N_103,In_313,In_6);
nand U104 (N_104,In_243,In_376);
or U105 (N_105,In_458,In_120);
nand U106 (N_106,In_53,In_328);
nor U107 (N_107,In_28,In_286);
xor U108 (N_108,In_323,In_483);
nand U109 (N_109,In_429,In_115);
nand U110 (N_110,In_404,In_114);
or U111 (N_111,In_466,In_362);
xnor U112 (N_112,In_498,In_141);
xnor U113 (N_113,In_417,In_187);
and U114 (N_114,In_49,In_145);
and U115 (N_115,In_357,In_183);
nor U116 (N_116,In_457,In_273);
and U117 (N_117,In_101,In_374);
xor U118 (N_118,In_180,In_470);
xor U119 (N_119,In_219,In_76);
nor U120 (N_120,In_186,In_80);
nor U121 (N_121,In_224,In_440);
xor U122 (N_122,In_199,In_146);
nor U123 (N_123,In_110,In_62);
nand U124 (N_124,In_124,In_430);
and U125 (N_125,In_46,In_326);
nor U126 (N_126,In_332,In_279);
and U127 (N_127,In_26,In_452);
nor U128 (N_128,In_151,In_345);
nor U129 (N_129,In_43,In_95);
nand U130 (N_130,In_327,In_414);
or U131 (N_131,In_237,In_138);
nand U132 (N_132,In_184,In_455);
nand U133 (N_133,In_51,In_105);
or U134 (N_134,In_348,In_242);
nor U135 (N_135,In_298,In_204);
xnor U136 (N_136,In_267,In_185);
and U137 (N_137,In_408,In_192);
nand U138 (N_138,In_155,In_351);
nand U139 (N_139,In_159,In_307);
nor U140 (N_140,In_170,In_297);
nand U141 (N_141,In_353,In_499);
nand U142 (N_142,In_161,In_25);
nor U143 (N_143,In_329,In_434);
nor U144 (N_144,In_85,In_369);
xor U145 (N_145,In_30,In_354);
or U146 (N_146,In_375,In_259);
xnor U147 (N_147,In_94,In_39);
and U148 (N_148,In_37,In_399);
nand U149 (N_149,In_478,In_424);
nand U150 (N_150,In_334,In_439);
or U151 (N_151,In_331,In_176);
xor U152 (N_152,In_265,In_132);
xnor U153 (N_153,In_129,In_188);
or U154 (N_154,In_83,In_56);
or U155 (N_155,In_427,In_196);
or U156 (N_156,In_127,In_195);
nor U157 (N_157,In_238,In_462);
or U158 (N_158,In_212,In_137);
xor U159 (N_159,In_108,In_367);
or U160 (N_160,In_446,In_418);
or U161 (N_161,In_269,In_449);
or U162 (N_162,In_247,In_285);
and U163 (N_163,In_387,In_40);
or U164 (N_164,In_249,In_461);
or U165 (N_165,In_472,In_206);
nor U166 (N_166,In_493,In_59);
or U167 (N_167,In_23,In_33);
or U168 (N_168,In_296,In_52);
nand U169 (N_169,In_123,In_406);
nand U170 (N_170,In_222,In_471);
nor U171 (N_171,In_117,In_303);
and U172 (N_172,In_139,In_433);
xnor U173 (N_173,In_289,In_102);
and U174 (N_174,In_174,In_485);
nor U175 (N_175,In_251,In_255);
or U176 (N_176,In_69,In_160);
nand U177 (N_177,In_454,In_48);
and U178 (N_178,In_213,In_65);
nor U179 (N_179,In_344,In_432);
nor U180 (N_180,In_100,In_314);
nor U181 (N_181,In_312,In_87);
nand U182 (N_182,In_365,In_57);
or U183 (N_183,In_198,In_142);
and U184 (N_184,In_480,In_119);
and U185 (N_185,In_197,In_420);
xor U186 (N_186,In_283,In_419);
and U187 (N_187,In_211,In_308);
nand U188 (N_188,In_469,In_360);
nor U189 (N_189,In_38,In_71);
xnor U190 (N_190,In_1,In_147);
nor U191 (N_191,In_10,In_443);
nand U192 (N_192,In_436,In_118);
nand U193 (N_193,In_405,In_167);
and U194 (N_194,In_82,In_24);
nand U195 (N_195,In_194,In_133);
xor U196 (N_196,In_393,In_15);
and U197 (N_197,In_336,In_284);
nor U198 (N_198,In_288,In_359);
nand U199 (N_199,In_412,In_261);
xor U200 (N_200,In_355,N_88);
nor U201 (N_201,In_107,N_130);
xnor U202 (N_202,In_371,N_37);
nand U203 (N_203,In_231,In_386);
nand U204 (N_204,In_337,In_134);
xor U205 (N_205,In_299,In_394);
and U206 (N_206,N_173,N_170);
nand U207 (N_207,N_57,In_66);
or U208 (N_208,N_9,In_220);
or U209 (N_209,N_7,N_83);
nand U210 (N_210,N_140,N_159);
and U211 (N_211,N_119,In_74);
nand U212 (N_212,N_70,N_120);
nand U213 (N_213,N_112,N_158);
nor U214 (N_214,N_67,N_38);
xor U215 (N_215,N_90,N_124);
nor U216 (N_216,In_122,N_107);
and U217 (N_217,N_2,In_29);
or U218 (N_218,N_103,N_139);
nor U219 (N_219,In_383,In_423);
or U220 (N_220,N_80,N_151);
or U221 (N_221,N_41,In_200);
and U222 (N_222,N_165,N_46);
and U223 (N_223,N_128,In_158);
nand U224 (N_224,In_236,N_102);
nand U225 (N_225,In_171,N_133);
or U226 (N_226,In_266,In_287);
nand U227 (N_227,N_18,N_42);
or U228 (N_228,In_54,N_21);
and U229 (N_229,N_28,N_121);
or U230 (N_230,In_268,In_467);
xnor U231 (N_231,In_293,In_0);
nand U232 (N_232,N_180,N_181);
nor U233 (N_233,In_221,N_95);
and U234 (N_234,In_416,N_68);
xor U235 (N_235,In_492,N_199);
nand U236 (N_236,In_276,N_50);
xnor U237 (N_237,N_51,N_27);
nand U238 (N_238,In_64,N_153);
and U239 (N_239,In_358,N_94);
and U240 (N_240,N_135,N_187);
and U241 (N_241,N_148,N_1);
and U242 (N_242,In_425,In_352);
or U243 (N_243,N_150,N_194);
xor U244 (N_244,N_185,N_3);
nand U245 (N_245,In_448,In_4);
or U246 (N_246,N_11,N_144);
nand U247 (N_247,N_190,N_177);
nor U248 (N_248,N_101,N_23);
nor U249 (N_249,N_193,N_164);
or U250 (N_250,N_10,In_22);
or U251 (N_251,N_113,In_300);
xor U252 (N_252,In_91,N_74);
and U253 (N_253,In_363,N_24);
and U254 (N_254,In_325,In_373);
nand U255 (N_255,N_108,N_157);
xnor U256 (N_256,N_54,N_35);
nor U257 (N_257,N_189,In_368);
nor U258 (N_258,In_390,In_385);
xnor U259 (N_259,N_43,N_123);
nor U260 (N_260,N_63,In_403);
xor U261 (N_261,N_71,In_156);
and U262 (N_262,N_22,In_21);
nand U263 (N_263,N_195,N_106);
xnor U264 (N_264,In_233,N_100);
nor U265 (N_265,N_86,N_197);
and U266 (N_266,N_84,N_64);
or U267 (N_267,N_176,N_55);
or U268 (N_268,N_174,N_141);
and U269 (N_269,N_122,In_494);
and U270 (N_270,N_97,N_40);
nand U271 (N_271,In_89,In_75);
xor U272 (N_272,N_138,N_126);
nor U273 (N_273,In_258,N_52);
xor U274 (N_274,In_47,In_411);
xor U275 (N_275,N_60,N_166);
nor U276 (N_276,N_171,N_12);
xor U277 (N_277,N_169,In_164);
and U278 (N_278,In_497,N_184);
and U279 (N_279,N_26,N_129);
nand U280 (N_280,N_0,In_456);
and U281 (N_281,N_92,N_79);
and U282 (N_282,In_163,In_12);
or U283 (N_283,N_98,N_178);
xnor U284 (N_284,N_183,N_182);
nand U285 (N_285,In_291,N_168);
nor U286 (N_286,In_201,In_460);
and U287 (N_287,N_155,N_82);
nor U288 (N_288,N_186,N_152);
and U289 (N_289,N_156,N_58);
or U290 (N_290,N_32,In_317);
nor U291 (N_291,N_89,N_134);
nor U292 (N_292,In_175,N_62);
and U293 (N_293,N_142,N_34);
or U294 (N_294,N_5,In_482);
or U295 (N_295,In_378,In_444);
nand U296 (N_296,N_78,In_447);
or U297 (N_297,In_70,In_396);
nand U298 (N_298,N_45,N_149);
xor U299 (N_299,N_4,In_340);
or U300 (N_300,N_19,N_115);
or U301 (N_301,N_48,In_109);
nor U302 (N_302,N_47,N_146);
and U303 (N_303,In_230,In_111);
nor U304 (N_304,N_59,N_117);
or U305 (N_305,N_125,N_17);
or U306 (N_306,N_147,N_105);
nor U307 (N_307,N_53,N_111);
nand U308 (N_308,In_271,N_66);
nand U309 (N_309,N_172,In_464);
nor U310 (N_310,In_241,N_49);
nor U311 (N_311,N_29,N_61);
and U312 (N_312,In_402,N_30);
nor U313 (N_313,N_13,N_44);
and U314 (N_314,N_25,In_310);
xnor U315 (N_315,N_72,N_85);
nand U316 (N_316,In_339,N_76);
or U317 (N_317,N_162,N_104);
or U318 (N_318,In_88,N_73);
and U319 (N_319,N_145,N_167);
nand U320 (N_320,N_163,In_217);
nand U321 (N_321,In_451,N_20);
xnor U322 (N_322,N_16,N_96);
and U323 (N_323,N_137,N_39);
xnor U324 (N_324,In_96,In_244);
nand U325 (N_325,N_143,In_445);
nand U326 (N_326,N_99,N_109);
or U327 (N_327,N_179,N_36);
nand U328 (N_328,N_6,N_56);
nor U329 (N_329,N_118,N_175);
nand U330 (N_330,In_42,In_252);
nand U331 (N_331,N_15,N_198);
xor U332 (N_332,In_154,In_356);
nor U333 (N_333,N_33,In_55);
and U334 (N_334,N_196,N_75);
and U335 (N_335,N_191,N_160);
nand U336 (N_336,N_77,N_116);
nand U337 (N_337,In_479,N_188);
and U338 (N_338,N_69,N_161);
and U339 (N_339,N_154,In_438);
or U340 (N_340,N_81,N_131);
xor U341 (N_341,N_87,N_91);
xnor U342 (N_342,N_192,N_31);
xnor U343 (N_343,N_65,N_14);
nor U344 (N_344,N_93,N_132);
nand U345 (N_345,N_110,In_225);
or U346 (N_346,N_114,N_136);
or U347 (N_347,N_8,In_5);
and U348 (N_348,In_338,In_234);
nor U349 (N_349,In_318,N_127);
nand U350 (N_350,In_416,N_81);
xor U351 (N_351,N_70,N_139);
nand U352 (N_352,In_230,N_122);
nor U353 (N_353,N_35,In_220);
nand U354 (N_354,In_363,N_138);
nand U355 (N_355,N_197,N_192);
nand U356 (N_356,In_21,In_74);
or U357 (N_357,N_1,In_175);
xor U358 (N_358,N_185,In_234);
nand U359 (N_359,In_74,N_108);
nand U360 (N_360,N_147,N_46);
and U361 (N_361,N_86,N_20);
or U362 (N_362,N_59,N_64);
and U363 (N_363,N_90,N_175);
nor U364 (N_364,N_131,N_156);
nor U365 (N_365,N_126,N_84);
and U366 (N_366,N_129,N_138);
nand U367 (N_367,N_50,N_161);
or U368 (N_368,In_467,N_91);
nand U369 (N_369,N_38,In_70);
xnor U370 (N_370,In_55,In_154);
nor U371 (N_371,N_55,N_28);
nor U372 (N_372,N_64,In_482);
nand U373 (N_373,N_171,N_149);
or U374 (N_374,In_55,N_175);
nor U375 (N_375,N_153,In_494);
and U376 (N_376,N_0,N_156);
or U377 (N_377,N_104,N_148);
or U378 (N_378,In_200,N_124);
xor U379 (N_379,N_54,In_371);
nand U380 (N_380,N_54,N_179);
and U381 (N_381,N_52,In_339);
xor U382 (N_382,In_447,N_70);
xnor U383 (N_383,N_120,N_197);
xor U384 (N_384,In_225,N_126);
and U385 (N_385,N_44,In_109);
or U386 (N_386,N_182,N_121);
and U387 (N_387,N_69,N_129);
xor U388 (N_388,In_217,N_138);
or U389 (N_389,N_172,N_33);
or U390 (N_390,N_135,In_266);
or U391 (N_391,In_325,N_63);
xnor U392 (N_392,In_134,N_181);
nand U393 (N_393,N_174,N_36);
nand U394 (N_394,N_108,In_200);
or U395 (N_395,N_79,N_149);
nor U396 (N_396,N_169,N_144);
nand U397 (N_397,In_54,In_122);
and U398 (N_398,N_175,N_120);
or U399 (N_399,N_68,In_171);
or U400 (N_400,N_222,N_204);
or U401 (N_401,N_240,N_274);
xnor U402 (N_402,N_369,N_216);
and U403 (N_403,N_244,N_374);
and U404 (N_404,N_285,N_366);
xor U405 (N_405,N_316,N_261);
or U406 (N_406,N_383,N_237);
and U407 (N_407,N_349,N_289);
nand U408 (N_408,N_245,N_296);
or U409 (N_409,N_334,N_267);
and U410 (N_410,N_276,N_231);
and U411 (N_411,N_229,N_365);
nand U412 (N_412,N_256,N_243);
nor U413 (N_413,N_338,N_246);
and U414 (N_414,N_208,N_309);
xor U415 (N_415,N_386,N_201);
xor U416 (N_416,N_337,N_311);
nor U417 (N_417,N_302,N_393);
and U418 (N_418,N_265,N_292);
and U419 (N_419,N_320,N_220);
nor U420 (N_420,N_226,N_249);
and U421 (N_421,N_368,N_340);
nand U422 (N_422,N_397,N_378);
nor U423 (N_423,N_271,N_205);
xnor U424 (N_424,N_317,N_336);
nor U425 (N_425,N_203,N_219);
xnor U426 (N_426,N_392,N_348);
and U427 (N_427,N_206,N_312);
and U428 (N_428,N_324,N_293);
nand U429 (N_429,N_364,N_234);
and U430 (N_430,N_253,N_225);
xor U431 (N_431,N_335,N_269);
nand U432 (N_432,N_298,N_211);
xnor U433 (N_433,N_343,N_279);
and U434 (N_434,N_347,N_357);
or U435 (N_435,N_248,N_236);
and U436 (N_436,N_318,N_356);
or U437 (N_437,N_282,N_218);
and U438 (N_438,N_328,N_341);
nor U439 (N_439,N_251,N_344);
or U440 (N_440,N_322,N_326);
xor U441 (N_441,N_270,N_315);
and U442 (N_442,N_278,N_329);
or U443 (N_443,N_352,N_370);
xnor U444 (N_444,N_387,N_323);
and U445 (N_445,N_373,N_227);
or U446 (N_446,N_358,N_254);
and U447 (N_447,N_228,N_307);
nand U448 (N_448,N_263,N_286);
nor U449 (N_449,N_310,N_262);
xnor U450 (N_450,N_332,N_390);
and U451 (N_451,N_259,N_272);
xnor U452 (N_452,N_295,N_207);
nand U453 (N_453,N_372,N_200);
xnor U454 (N_454,N_345,N_301);
nand U455 (N_455,N_255,N_210);
nand U456 (N_456,N_327,N_233);
or U457 (N_457,N_388,N_221);
xnor U458 (N_458,N_297,N_223);
xnor U459 (N_459,N_213,N_304);
and U460 (N_460,N_353,N_252);
and U461 (N_461,N_367,N_280);
xnor U462 (N_462,N_242,N_232);
or U463 (N_463,N_291,N_362);
nand U464 (N_464,N_238,N_371);
nand U465 (N_465,N_377,N_394);
xor U466 (N_466,N_308,N_381);
or U467 (N_467,N_287,N_257);
or U468 (N_468,N_235,N_268);
or U469 (N_469,N_283,N_342);
nor U470 (N_470,N_399,N_314);
and U471 (N_471,N_277,N_351);
xor U472 (N_472,N_380,N_375);
and U473 (N_473,N_350,N_379);
nor U474 (N_474,N_260,N_212);
nand U475 (N_475,N_319,N_209);
xor U476 (N_476,N_273,N_266);
and U477 (N_477,N_214,N_331);
nor U478 (N_478,N_346,N_275);
nand U479 (N_479,N_306,N_224);
or U480 (N_480,N_288,N_215);
nor U481 (N_481,N_264,N_284);
nor U482 (N_482,N_391,N_360);
nand U483 (N_483,N_300,N_395);
xnor U484 (N_484,N_230,N_250);
nand U485 (N_485,N_217,N_361);
and U486 (N_486,N_363,N_355);
and U487 (N_487,N_247,N_299);
nand U488 (N_488,N_359,N_202);
nor U489 (N_489,N_376,N_339);
or U490 (N_490,N_385,N_382);
xnor U491 (N_491,N_294,N_239);
nor U492 (N_492,N_330,N_389);
xnor U493 (N_493,N_333,N_396);
and U494 (N_494,N_281,N_305);
nand U495 (N_495,N_398,N_354);
nand U496 (N_496,N_384,N_241);
xor U497 (N_497,N_325,N_303);
xnor U498 (N_498,N_313,N_258);
xor U499 (N_499,N_290,N_321);
and U500 (N_500,N_229,N_392);
nand U501 (N_501,N_395,N_218);
or U502 (N_502,N_278,N_220);
nand U503 (N_503,N_319,N_292);
and U504 (N_504,N_351,N_242);
or U505 (N_505,N_340,N_280);
nor U506 (N_506,N_309,N_347);
nor U507 (N_507,N_383,N_251);
xnor U508 (N_508,N_394,N_334);
nor U509 (N_509,N_274,N_291);
nor U510 (N_510,N_301,N_351);
or U511 (N_511,N_206,N_351);
nor U512 (N_512,N_345,N_389);
or U513 (N_513,N_333,N_314);
nor U514 (N_514,N_357,N_313);
and U515 (N_515,N_330,N_392);
and U516 (N_516,N_322,N_385);
or U517 (N_517,N_276,N_359);
and U518 (N_518,N_255,N_208);
nor U519 (N_519,N_281,N_205);
xor U520 (N_520,N_234,N_250);
nand U521 (N_521,N_212,N_379);
nand U522 (N_522,N_381,N_355);
or U523 (N_523,N_363,N_273);
or U524 (N_524,N_332,N_353);
or U525 (N_525,N_318,N_244);
or U526 (N_526,N_335,N_376);
or U527 (N_527,N_365,N_393);
or U528 (N_528,N_324,N_238);
and U529 (N_529,N_261,N_356);
and U530 (N_530,N_255,N_266);
nand U531 (N_531,N_272,N_391);
nor U532 (N_532,N_320,N_380);
and U533 (N_533,N_323,N_223);
xnor U534 (N_534,N_277,N_233);
nand U535 (N_535,N_277,N_257);
xor U536 (N_536,N_366,N_271);
or U537 (N_537,N_359,N_265);
nor U538 (N_538,N_314,N_329);
xnor U539 (N_539,N_225,N_223);
nor U540 (N_540,N_238,N_281);
and U541 (N_541,N_207,N_322);
nor U542 (N_542,N_261,N_353);
nor U543 (N_543,N_266,N_295);
nor U544 (N_544,N_221,N_276);
xor U545 (N_545,N_353,N_395);
nor U546 (N_546,N_298,N_291);
and U547 (N_547,N_316,N_253);
and U548 (N_548,N_319,N_237);
or U549 (N_549,N_242,N_317);
xnor U550 (N_550,N_387,N_362);
xnor U551 (N_551,N_214,N_347);
nand U552 (N_552,N_239,N_344);
nor U553 (N_553,N_270,N_272);
nor U554 (N_554,N_242,N_274);
nor U555 (N_555,N_290,N_388);
nand U556 (N_556,N_246,N_278);
and U557 (N_557,N_283,N_367);
or U558 (N_558,N_289,N_370);
nand U559 (N_559,N_266,N_292);
nand U560 (N_560,N_280,N_388);
and U561 (N_561,N_381,N_340);
nor U562 (N_562,N_280,N_372);
nor U563 (N_563,N_348,N_241);
or U564 (N_564,N_367,N_355);
xnor U565 (N_565,N_265,N_204);
or U566 (N_566,N_270,N_335);
or U567 (N_567,N_355,N_347);
xor U568 (N_568,N_273,N_378);
xnor U569 (N_569,N_265,N_338);
or U570 (N_570,N_207,N_345);
xor U571 (N_571,N_386,N_271);
xnor U572 (N_572,N_300,N_367);
nand U573 (N_573,N_286,N_298);
and U574 (N_574,N_298,N_225);
or U575 (N_575,N_374,N_384);
nand U576 (N_576,N_354,N_366);
nand U577 (N_577,N_219,N_261);
or U578 (N_578,N_292,N_371);
and U579 (N_579,N_270,N_256);
nor U580 (N_580,N_295,N_322);
nor U581 (N_581,N_390,N_342);
or U582 (N_582,N_323,N_247);
and U583 (N_583,N_208,N_263);
and U584 (N_584,N_259,N_203);
nand U585 (N_585,N_280,N_278);
nand U586 (N_586,N_207,N_286);
nand U587 (N_587,N_236,N_216);
xnor U588 (N_588,N_279,N_350);
xnor U589 (N_589,N_210,N_254);
nand U590 (N_590,N_369,N_291);
nor U591 (N_591,N_316,N_220);
and U592 (N_592,N_221,N_271);
nand U593 (N_593,N_312,N_330);
or U594 (N_594,N_383,N_238);
xor U595 (N_595,N_272,N_343);
nor U596 (N_596,N_351,N_245);
and U597 (N_597,N_283,N_268);
or U598 (N_598,N_246,N_256);
or U599 (N_599,N_258,N_204);
nand U600 (N_600,N_579,N_447);
nor U601 (N_601,N_450,N_592);
or U602 (N_602,N_488,N_509);
and U603 (N_603,N_591,N_465);
nand U604 (N_604,N_444,N_584);
nor U605 (N_605,N_451,N_479);
nand U606 (N_606,N_484,N_470);
or U607 (N_607,N_569,N_422);
and U608 (N_608,N_515,N_421);
or U609 (N_609,N_504,N_405);
nand U610 (N_610,N_524,N_463);
nand U611 (N_611,N_525,N_483);
nor U612 (N_612,N_431,N_429);
nor U613 (N_613,N_566,N_523);
nand U614 (N_614,N_555,N_564);
or U615 (N_615,N_439,N_597);
nor U616 (N_616,N_559,N_599);
nor U617 (N_617,N_590,N_578);
and U618 (N_618,N_454,N_589);
or U619 (N_619,N_430,N_588);
or U620 (N_620,N_542,N_593);
nand U621 (N_621,N_471,N_527);
or U622 (N_622,N_496,N_434);
and U623 (N_623,N_554,N_416);
xor U624 (N_624,N_413,N_459);
nor U625 (N_625,N_464,N_548);
nor U626 (N_626,N_576,N_533);
and U627 (N_627,N_546,N_433);
or U628 (N_628,N_445,N_475);
or U629 (N_629,N_580,N_577);
xor U630 (N_630,N_507,N_538);
and U631 (N_631,N_521,N_478);
or U632 (N_632,N_587,N_449);
nand U633 (N_633,N_474,N_508);
nor U634 (N_634,N_410,N_428);
xor U635 (N_635,N_531,N_598);
and U636 (N_636,N_506,N_565);
and U637 (N_637,N_520,N_477);
and U638 (N_638,N_424,N_539);
and U639 (N_639,N_582,N_518);
nand U640 (N_640,N_408,N_452);
xor U641 (N_641,N_446,N_594);
nor U642 (N_642,N_519,N_522);
nand U643 (N_643,N_406,N_400);
xor U644 (N_644,N_402,N_420);
or U645 (N_645,N_499,N_516);
xnor U646 (N_646,N_498,N_487);
xor U647 (N_647,N_404,N_571);
and U648 (N_648,N_411,N_540);
xnor U649 (N_649,N_415,N_455);
nor U650 (N_650,N_562,N_423);
nor U651 (N_651,N_510,N_417);
nor U652 (N_652,N_403,N_543);
nand U653 (N_653,N_526,N_448);
and U654 (N_654,N_556,N_502);
nor U655 (N_655,N_456,N_468);
xor U656 (N_656,N_586,N_409);
nor U657 (N_657,N_442,N_419);
nand U658 (N_658,N_440,N_435);
xnor U659 (N_659,N_407,N_414);
nor U660 (N_660,N_494,N_561);
nand U661 (N_661,N_437,N_476);
and U662 (N_662,N_472,N_441);
xnor U663 (N_663,N_466,N_558);
xor U664 (N_664,N_505,N_560);
or U665 (N_665,N_575,N_547);
and U666 (N_666,N_492,N_427);
xor U667 (N_667,N_552,N_534);
xnor U668 (N_668,N_567,N_493);
nor U669 (N_669,N_432,N_473);
and U670 (N_670,N_425,N_536);
nand U671 (N_671,N_570,N_528);
and U672 (N_672,N_568,N_500);
or U673 (N_673,N_460,N_596);
or U674 (N_674,N_486,N_563);
or U675 (N_675,N_557,N_501);
nand U676 (N_676,N_482,N_495);
or U677 (N_677,N_458,N_490);
xnor U678 (N_678,N_443,N_489);
or U679 (N_679,N_595,N_457);
or U680 (N_680,N_401,N_545);
xor U681 (N_681,N_573,N_436);
and U682 (N_682,N_480,N_514);
xnor U683 (N_683,N_549,N_530);
and U684 (N_684,N_544,N_550);
nand U685 (N_685,N_551,N_412);
and U686 (N_686,N_535,N_512);
nand U687 (N_687,N_585,N_438);
or U688 (N_688,N_529,N_461);
nand U689 (N_689,N_453,N_426);
or U690 (N_690,N_467,N_497);
nand U691 (N_691,N_462,N_572);
and U692 (N_692,N_503,N_517);
and U693 (N_693,N_485,N_541);
or U694 (N_694,N_491,N_574);
nor U695 (N_695,N_553,N_418);
xor U696 (N_696,N_537,N_581);
and U697 (N_697,N_513,N_532);
or U698 (N_698,N_583,N_481);
xor U699 (N_699,N_511,N_469);
nor U700 (N_700,N_457,N_429);
xor U701 (N_701,N_578,N_459);
nor U702 (N_702,N_482,N_531);
nand U703 (N_703,N_550,N_579);
or U704 (N_704,N_443,N_439);
nor U705 (N_705,N_503,N_407);
and U706 (N_706,N_507,N_422);
nor U707 (N_707,N_447,N_418);
nand U708 (N_708,N_569,N_587);
nand U709 (N_709,N_483,N_558);
and U710 (N_710,N_596,N_502);
and U711 (N_711,N_525,N_512);
and U712 (N_712,N_543,N_546);
nand U713 (N_713,N_412,N_414);
or U714 (N_714,N_477,N_584);
xnor U715 (N_715,N_506,N_558);
or U716 (N_716,N_524,N_589);
nor U717 (N_717,N_400,N_504);
nand U718 (N_718,N_538,N_447);
or U719 (N_719,N_416,N_579);
nor U720 (N_720,N_432,N_426);
and U721 (N_721,N_579,N_563);
xor U722 (N_722,N_436,N_524);
or U723 (N_723,N_505,N_470);
and U724 (N_724,N_415,N_584);
xnor U725 (N_725,N_548,N_536);
or U726 (N_726,N_591,N_544);
xnor U727 (N_727,N_426,N_435);
nand U728 (N_728,N_587,N_562);
and U729 (N_729,N_551,N_405);
or U730 (N_730,N_455,N_557);
nand U731 (N_731,N_568,N_531);
or U732 (N_732,N_557,N_477);
xnor U733 (N_733,N_523,N_506);
nand U734 (N_734,N_583,N_448);
or U735 (N_735,N_407,N_496);
nor U736 (N_736,N_567,N_416);
nand U737 (N_737,N_461,N_403);
and U738 (N_738,N_428,N_422);
nand U739 (N_739,N_588,N_419);
nand U740 (N_740,N_475,N_488);
nand U741 (N_741,N_579,N_420);
or U742 (N_742,N_590,N_441);
nand U743 (N_743,N_581,N_506);
xor U744 (N_744,N_544,N_503);
nor U745 (N_745,N_565,N_456);
and U746 (N_746,N_587,N_413);
xor U747 (N_747,N_424,N_400);
nor U748 (N_748,N_481,N_469);
nand U749 (N_749,N_412,N_555);
nand U750 (N_750,N_477,N_560);
or U751 (N_751,N_442,N_464);
and U752 (N_752,N_557,N_561);
and U753 (N_753,N_506,N_415);
and U754 (N_754,N_492,N_499);
nand U755 (N_755,N_488,N_409);
and U756 (N_756,N_516,N_439);
or U757 (N_757,N_490,N_460);
nand U758 (N_758,N_473,N_507);
xnor U759 (N_759,N_596,N_576);
and U760 (N_760,N_503,N_401);
xor U761 (N_761,N_418,N_483);
or U762 (N_762,N_410,N_497);
and U763 (N_763,N_516,N_501);
or U764 (N_764,N_443,N_563);
and U765 (N_765,N_595,N_556);
and U766 (N_766,N_590,N_462);
or U767 (N_767,N_548,N_456);
or U768 (N_768,N_484,N_429);
nand U769 (N_769,N_544,N_439);
or U770 (N_770,N_532,N_444);
and U771 (N_771,N_516,N_454);
nor U772 (N_772,N_403,N_508);
nor U773 (N_773,N_469,N_405);
or U774 (N_774,N_510,N_551);
xor U775 (N_775,N_479,N_557);
nor U776 (N_776,N_491,N_401);
nor U777 (N_777,N_494,N_402);
xor U778 (N_778,N_539,N_500);
or U779 (N_779,N_497,N_443);
nor U780 (N_780,N_568,N_593);
and U781 (N_781,N_476,N_471);
nor U782 (N_782,N_577,N_500);
or U783 (N_783,N_520,N_415);
nor U784 (N_784,N_573,N_500);
nor U785 (N_785,N_533,N_535);
xnor U786 (N_786,N_550,N_455);
and U787 (N_787,N_522,N_405);
or U788 (N_788,N_419,N_581);
and U789 (N_789,N_593,N_582);
nor U790 (N_790,N_509,N_483);
nand U791 (N_791,N_528,N_416);
and U792 (N_792,N_478,N_414);
nand U793 (N_793,N_434,N_424);
nand U794 (N_794,N_446,N_501);
and U795 (N_795,N_446,N_566);
nor U796 (N_796,N_488,N_442);
or U797 (N_797,N_566,N_555);
and U798 (N_798,N_423,N_586);
nand U799 (N_799,N_463,N_413);
and U800 (N_800,N_647,N_610);
nand U801 (N_801,N_778,N_615);
nand U802 (N_802,N_606,N_718);
xor U803 (N_803,N_795,N_691);
and U804 (N_804,N_627,N_739);
and U805 (N_805,N_765,N_721);
xnor U806 (N_806,N_640,N_629);
xnor U807 (N_807,N_658,N_614);
and U808 (N_808,N_790,N_632);
or U809 (N_809,N_793,N_748);
and U810 (N_810,N_684,N_603);
and U811 (N_811,N_730,N_744);
and U812 (N_812,N_751,N_667);
or U813 (N_813,N_693,N_673);
and U814 (N_814,N_668,N_738);
and U815 (N_815,N_787,N_723);
nand U816 (N_816,N_724,N_659);
nor U817 (N_817,N_764,N_621);
nor U818 (N_818,N_653,N_690);
or U819 (N_819,N_754,N_758);
nor U820 (N_820,N_752,N_734);
xnor U821 (N_821,N_685,N_678);
or U822 (N_822,N_650,N_605);
and U823 (N_823,N_789,N_637);
xnor U824 (N_824,N_742,N_745);
nor U825 (N_825,N_657,N_737);
nor U826 (N_826,N_676,N_722);
nand U827 (N_827,N_607,N_686);
nor U828 (N_828,N_689,N_631);
or U829 (N_829,N_639,N_717);
xor U830 (N_830,N_783,N_604);
and U831 (N_831,N_648,N_706);
and U832 (N_832,N_756,N_772);
or U833 (N_833,N_620,N_645);
nor U834 (N_834,N_712,N_600);
xnor U835 (N_835,N_763,N_628);
xor U836 (N_836,N_710,N_630);
nand U837 (N_837,N_771,N_731);
and U838 (N_838,N_687,N_609);
xnor U839 (N_839,N_677,N_635);
nor U840 (N_840,N_773,N_683);
or U841 (N_841,N_746,N_695);
nor U842 (N_842,N_702,N_799);
nor U843 (N_843,N_762,N_633);
and U844 (N_844,N_665,N_675);
nor U845 (N_845,N_708,N_726);
xnor U846 (N_846,N_661,N_617);
xor U847 (N_847,N_651,N_688);
nand U848 (N_848,N_619,N_774);
nor U849 (N_849,N_612,N_743);
xnor U850 (N_850,N_796,N_707);
xnor U851 (N_851,N_732,N_670);
xnor U852 (N_852,N_644,N_750);
nor U853 (N_853,N_643,N_666);
and U854 (N_854,N_757,N_641);
nor U855 (N_855,N_692,N_798);
xnor U856 (N_856,N_785,N_608);
nand U857 (N_857,N_791,N_733);
xor U858 (N_858,N_664,N_662);
xnor U859 (N_859,N_770,N_618);
nor U860 (N_860,N_611,N_699);
xor U861 (N_861,N_696,N_705);
or U862 (N_862,N_613,N_735);
or U863 (N_863,N_719,N_680);
nand U864 (N_864,N_786,N_652);
nand U865 (N_865,N_716,N_741);
and U866 (N_866,N_601,N_674);
or U867 (N_867,N_655,N_715);
and U868 (N_868,N_700,N_749);
nand U869 (N_869,N_642,N_624);
or U870 (N_870,N_703,N_681);
or U871 (N_871,N_760,N_672);
or U872 (N_872,N_679,N_711);
or U873 (N_873,N_602,N_697);
nor U874 (N_874,N_797,N_669);
or U875 (N_875,N_780,N_788);
or U876 (N_876,N_779,N_755);
nor U877 (N_877,N_759,N_616);
and U878 (N_878,N_794,N_713);
nor U879 (N_879,N_792,N_775);
and U880 (N_880,N_761,N_725);
or U881 (N_881,N_777,N_634);
and U882 (N_882,N_660,N_626);
nand U883 (N_883,N_714,N_656);
xor U884 (N_884,N_727,N_646);
or U885 (N_885,N_698,N_701);
or U886 (N_886,N_736,N_654);
nor U887 (N_887,N_766,N_782);
and U888 (N_888,N_622,N_747);
nor U889 (N_889,N_623,N_753);
nor U890 (N_890,N_636,N_625);
or U891 (N_891,N_694,N_649);
nand U892 (N_892,N_728,N_781);
nor U893 (N_893,N_663,N_784);
xnor U894 (N_894,N_740,N_638);
nand U895 (N_895,N_768,N_767);
and U896 (N_896,N_682,N_720);
and U897 (N_897,N_671,N_729);
xor U898 (N_898,N_769,N_709);
nand U899 (N_899,N_704,N_776);
and U900 (N_900,N_731,N_673);
nor U901 (N_901,N_769,N_761);
nor U902 (N_902,N_694,N_770);
nand U903 (N_903,N_750,N_753);
xnor U904 (N_904,N_777,N_682);
and U905 (N_905,N_741,N_734);
xor U906 (N_906,N_653,N_673);
or U907 (N_907,N_695,N_630);
nor U908 (N_908,N_707,N_743);
nand U909 (N_909,N_650,N_668);
nor U910 (N_910,N_794,N_635);
nand U911 (N_911,N_745,N_748);
nor U912 (N_912,N_649,N_667);
xor U913 (N_913,N_676,N_692);
and U914 (N_914,N_627,N_619);
xor U915 (N_915,N_610,N_770);
or U916 (N_916,N_768,N_652);
xor U917 (N_917,N_690,N_769);
or U918 (N_918,N_736,N_651);
nand U919 (N_919,N_719,N_689);
or U920 (N_920,N_676,N_666);
or U921 (N_921,N_660,N_728);
nor U922 (N_922,N_646,N_752);
nand U923 (N_923,N_636,N_628);
xnor U924 (N_924,N_605,N_789);
nand U925 (N_925,N_776,N_720);
nand U926 (N_926,N_785,N_679);
nor U927 (N_927,N_633,N_780);
or U928 (N_928,N_713,N_661);
xor U929 (N_929,N_786,N_623);
nand U930 (N_930,N_634,N_606);
xnor U931 (N_931,N_636,N_688);
or U932 (N_932,N_655,N_625);
and U933 (N_933,N_646,N_613);
xnor U934 (N_934,N_685,N_644);
nor U935 (N_935,N_706,N_655);
xor U936 (N_936,N_639,N_689);
nor U937 (N_937,N_667,N_700);
nor U938 (N_938,N_644,N_665);
or U939 (N_939,N_778,N_696);
xor U940 (N_940,N_724,N_729);
and U941 (N_941,N_660,N_710);
xor U942 (N_942,N_730,N_759);
or U943 (N_943,N_619,N_604);
and U944 (N_944,N_730,N_619);
nand U945 (N_945,N_673,N_697);
and U946 (N_946,N_758,N_680);
nor U947 (N_947,N_602,N_751);
and U948 (N_948,N_649,N_751);
nor U949 (N_949,N_685,N_765);
nor U950 (N_950,N_749,N_792);
xor U951 (N_951,N_664,N_657);
nand U952 (N_952,N_766,N_771);
xnor U953 (N_953,N_766,N_745);
xnor U954 (N_954,N_709,N_705);
nor U955 (N_955,N_795,N_667);
or U956 (N_956,N_728,N_717);
or U957 (N_957,N_637,N_774);
nand U958 (N_958,N_757,N_600);
xor U959 (N_959,N_606,N_686);
or U960 (N_960,N_611,N_609);
xor U961 (N_961,N_635,N_727);
nand U962 (N_962,N_726,N_751);
nor U963 (N_963,N_680,N_777);
and U964 (N_964,N_725,N_700);
and U965 (N_965,N_672,N_727);
or U966 (N_966,N_674,N_739);
and U967 (N_967,N_714,N_718);
nor U968 (N_968,N_609,N_728);
or U969 (N_969,N_655,N_747);
xor U970 (N_970,N_776,N_746);
nor U971 (N_971,N_636,N_610);
xor U972 (N_972,N_647,N_619);
nor U973 (N_973,N_718,N_693);
and U974 (N_974,N_655,N_667);
or U975 (N_975,N_739,N_631);
xor U976 (N_976,N_710,N_619);
xor U977 (N_977,N_773,N_731);
xor U978 (N_978,N_658,N_700);
and U979 (N_979,N_796,N_645);
xor U980 (N_980,N_720,N_670);
or U981 (N_981,N_638,N_726);
nand U982 (N_982,N_621,N_687);
or U983 (N_983,N_732,N_664);
or U984 (N_984,N_640,N_799);
nand U985 (N_985,N_680,N_753);
or U986 (N_986,N_663,N_779);
xor U987 (N_987,N_799,N_782);
nand U988 (N_988,N_685,N_742);
and U989 (N_989,N_665,N_715);
nand U990 (N_990,N_694,N_740);
nand U991 (N_991,N_790,N_700);
nand U992 (N_992,N_604,N_659);
and U993 (N_993,N_621,N_679);
nand U994 (N_994,N_688,N_674);
nor U995 (N_995,N_684,N_755);
xnor U996 (N_996,N_609,N_706);
xor U997 (N_997,N_739,N_647);
or U998 (N_998,N_621,N_635);
or U999 (N_999,N_666,N_707);
or U1000 (N_1000,N_874,N_849);
and U1001 (N_1001,N_956,N_975);
nand U1002 (N_1002,N_830,N_808);
and U1003 (N_1003,N_887,N_816);
and U1004 (N_1004,N_854,N_916);
xor U1005 (N_1005,N_805,N_933);
nor U1006 (N_1006,N_983,N_813);
or U1007 (N_1007,N_811,N_831);
and U1008 (N_1008,N_869,N_803);
nand U1009 (N_1009,N_826,N_952);
nand U1010 (N_1010,N_878,N_827);
xnor U1011 (N_1011,N_876,N_832);
nor U1012 (N_1012,N_911,N_865);
or U1013 (N_1013,N_927,N_839);
or U1014 (N_1014,N_947,N_877);
nand U1015 (N_1015,N_898,N_972);
xnor U1016 (N_1016,N_879,N_840);
and U1017 (N_1017,N_939,N_906);
nand U1018 (N_1018,N_809,N_868);
and U1019 (N_1019,N_838,N_930);
xnor U1020 (N_1020,N_988,N_902);
and U1021 (N_1021,N_821,N_872);
xor U1022 (N_1022,N_938,N_885);
or U1023 (N_1023,N_934,N_950);
xor U1024 (N_1024,N_932,N_920);
or U1025 (N_1025,N_817,N_800);
xnor U1026 (N_1026,N_856,N_814);
or U1027 (N_1027,N_941,N_867);
nand U1028 (N_1028,N_833,N_993);
xnor U1029 (N_1029,N_863,N_844);
and U1030 (N_1030,N_900,N_894);
xor U1031 (N_1031,N_922,N_995);
xnor U1032 (N_1032,N_946,N_967);
or U1033 (N_1033,N_974,N_982);
xor U1034 (N_1034,N_979,N_893);
xor U1035 (N_1035,N_918,N_819);
nand U1036 (N_1036,N_908,N_858);
nand U1037 (N_1037,N_822,N_945);
nor U1038 (N_1038,N_812,N_815);
nor U1039 (N_1039,N_870,N_954);
xor U1040 (N_1040,N_961,N_855);
xnor U1041 (N_1041,N_823,N_861);
xor U1042 (N_1042,N_901,N_969);
nor U1043 (N_1043,N_853,N_896);
xor U1044 (N_1044,N_966,N_905);
nand U1045 (N_1045,N_936,N_940);
xnor U1046 (N_1046,N_977,N_909);
or U1047 (N_1047,N_804,N_985);
nand U1048 (N_1048,N_978,N_976);
or U1049 (N_1049,N_992,N_802);
or U1050 (N_1050,N_889,N_997);
nand U1051 (N_1051,N_944,N_964);
and U1052 (N_1052,N_824,N_828);
and U1053 (N_1053,N_955,N_834);
or U1054 (N_1054,N_829,N_953);
nand U1055 (N_1055,N_951,N_903);
and U1056 (N_1056,N_990,N_937);
or U1057 (N_1057,N_980,N_994);
nand U1058 (N_1058,N_960,N_852);
or U1059 (N_1059,N_860,N_913);
or U1060 (N_1060,N_904,N_931);
or U1061 (N_1061,N_881,N_917);
xnor U1062 (N_1062,N_957,N_910);
and U1063 (N_1063,N_847,N_971);
nor U1064 (N_1064,N_801,N_970);
nor U1065 (N_1065,N_818,N_890);
and U1066 (N_1066,N_897,N_871);
or U1067 (N_1067,N_880,N_959);
nand U1068 (N_1068,N_943,N_851);
or U1069 (N_1069,N_843,N_912);
nor U1070 (N_1070,N_987,N_899);
nor U1071 (N_1071,N_806,N_973);
or U1072 (N_1072,N_883,N_984);
and U1073 (N_1073,N_928,N_935);
xor U1074 (N_1074,N_857,N_859);
nand U1075 (N_1075,N_942,N_810);
and U1076 (N_1076,N_996,N_875);
nand U1077 (N_1077,N_929,N_891);
or U1078 (N_1078,N_921,N_835);
and U1079 (N_1079,N_884,N_825);
and U1080 (N_1080,N_965,N_914);
and U1081 (N_1081,N_949,N_998);
xnor U1082 (N_1082,N_925,N_850);
nor U1083 (N_1083,N_907,N_968);
xor U1084 (N_1084,N_836,N_963);
nor U1085 (N_1085,N_986,N_807);
xnor U1086 (N_1086,N_841,N_962);
and U1087 (N_1087,N_915,N_888);
and U1088 (N_1088,N_895,N_873);
and U1089 (N_1089,N_892,N_919);
nand U1090 (N_1090,N_864,N_923);
nor U1091 (N_1091,N_846,N_989);
or U1092 (N_1092,N_991,N_958);
and U1093 (N_1093,N_886,N_882);
and U1094 (N_1094,N_820,N_837);
or U1095 (N_1095,N_999,N_848);
or U1096 (N_1096,N_866,N_862);
nand U1097 (N_1097,N_981,N_924);
or U1098 (N_1098,N_926,N_842);
nor U1099 (N_1099,N_948,N_845);
and U1100 (N_1100,N_936,N_842);
nand U1101 (N_1101,N_930,N_938);
and U1102 (N_1102,N_857,N_978);
nor U1103 (N_1103,N_823,N_841);
xnor U1104 (N_1104,N_970,N_924);
xnor U1105 (N_1105,N_862,N_951);
or U1106 (N_1106,N_805,N_839);
nand U1107 (N_1107,N_956,N_808);
nor U1108 (N_1108,N_970,N_820);
xor U1109 (N_1109,N_916,N_903);
or U1110 (N_1110,N_988,N_972);
nor U1111 (N_1111,N_843,N_927);
or U1112 (N_1112,N_810,N_801);
nand U1113 (N_1113,N_931,N_971);
or U1114 (N_1114,N_830,N_944);
or U1115 (N_1115,N_928,N_961);
and U1116 (N_1116,N_823,N_876);
and U1117 (N_1117,N_883,N_817);
nor U1118 (N_1118,N_819,N_892);
or U1119 (N_1119,N_877,N_893);
xor U1120 (N_1120,N_833,N_848);
nand U1121 (N_1121,N_921,N_994);
nand U1122 (N_1122,N_981,N_937);
nand U1123 (N_1123,N_925,N_806);
nand U1124 (N_1124,N_869,N_937);
and U1125 (N_1125,N_809,N_918);
xor U1126 (N_1126,N_824,N_906);
xnor U1127 (N_1127,N_907,N_873);
xor U1128 (N_1128,N_832,N_972);
nor U1129 (N_1129,N_957,N_968);
and U1130 (N_1130,N_995,N_824);
and U1131 (N_1131,N_967,N_972);
and U1132 (N_1132,N_855,N_925);
or U1133 (N_1133,N_931,N_890);
and U1134 (N_1134,N_883,N_818);
xnor U1135 (N_1135,N_835,N_830);
and U1136 (N_1136,N_890,N_917);
nor U1137 (N_1137,N_853,N_974);
nor U1138 (N_1138,N_863,N_919);
nor U1139 (N_1139,N_857,N_823);
nand U1140 (N_1140,N_818,N_913);
and U1141 (N_1141,N_963,N_933);
nor U1142 (N_1142,N_941,N_801);
nor U1143 (N_1143,N_919,N_960);
and U1144 (N_1144,N_860,N_821);
and U1145 (N_1145,N_908,N_953);
or U1146 (N_1146,N_914,N_866);
and U1147 (N_1147,N_849,N_837);
nand U1148 (N_1148,N_993,N_951);
or U1149 (N_1149,N_969,N_970);
xnor U1150 (N_1150,N_882,N_988);
or U1151 (N_1151,N_865,N_980);
nor U1152 (N_1152,N_825,N_892);
xor U1153 (N_1153,N_816,N_807);
and U1154 (N_1154,N_964,N_945);
and U1155 (N_1155,N_837,N_975);
and U1156 (N_1156,N_958,N_933);
nand U1157 (N_1157,N_886,N_910);
xnor U1158 (N_1158,N_968,N_825);
nor U1159 (N_1159,N_809,N_925);
xnor U1160 (N_1160,N_828,N_823);
and U1161 (N_1161,N_928,N_824);
xnor U1162 (N_1162,N_924,N_882);
or U1163 (N_1163,N_983,N_944);
or U1164 (N_1164,N_954,N_853);
nand U1165 (N_1165,N_836,N_837);
nand U1166 (N_1166,N_827,N_910);
nand U1167 (N_1167,N_817,N_854);
and U1168 (N_1168,N_801,N_825);
or U1169 (N_1169,N_865,N_985);
or U1170 (N_1170,N_982,N_869);
xor U1171 (N_1171,N_878,N_874);
nand U1172 (N_1172,N_942,N_829);
or U1173 (N_1173,N_936,N_946);
and U1174 (N_1174,N_957,N_822);
xnor U1175 (N_1175,N_847,N_882);
nor U1176 (N_1176,N_834,N_947);
and U1177 (N_1177,N_824,N_834);
and U1178 (N_1178,N_953,N_803);
xor U1179 (N_1179,N_819,N_925);
and U1180 (N_1180,N_989,N_821);
xor U1181 (N_1181,N_865,N_886);
nor U1182 (N_1182,N_869,N_887);
nand U1183 (N_1183,N_937,N_866);
and U1184 (N_1184,N_914,N_864);
or U1185 (N_1185,N_948,N_804);
and U1186 (N_1186,N_997,N_944);
nand U1187 (N_1187,N_909,N_847);
nand U1188 (N_1188,N_970,N_916);
xor U1189 (N_1189,N_830,N_880);
nor U1190 (N_1190,N_931,N_818);
nand U1191 (N_1191,N_859,N_802);
xor U1192 (N_1192,N_860,N_950);
and U1193 (N_1193,N_817,N_963);
nor U1194 (N_1194,N_923,N_861);
xor U1195 (N_1195,N_827,N_830);
or U1196 (N_1196,N_818,N_858);
and U1197 (N_1197,N_969,N_896);
nand U1198 (N_1198,N_962,N_912);
xor U1199 (N_1199,N_867,N_912);
nand U1200 (N_1200,N_1147,N_1091);
or U1201 (N_1201,N_1018,N_1079);
nor U1202 (N_1202,N_1136,N_1043);
nand U1203 (N_1203,N_1123,N_1001);
and U1204 (N_1204,N_1060,N_1089);
or U1205 (N_1205,N_1139,N_1116);
and U1206 (N_1206,N_1087,N_1110);
xnor U1207 (N_1207,N_1048,N_1085);
and U1208 (N_1208,N_1167,N_1101);
and U1209 (N_1209,N_1005,N_1163);
nand U1210 (N_1210,N_1190,N_1099);
nand U1211 (N_1211,N_1040,N_1002);
nand U1212 (N_1212,N_1143,N_1119);
or U1213 (N_1213,N_1198,N_1105);
xnor U1214 (N_1214,N_1028,N_1093);
xnor U1215 (N_1215,N_1017,N_1042);
and U1216 (N_1216,N_1192,N_1193);
or U1217 (N_1217,N_1035,N_1014);
and U1218 (N_1218,N_1088,N_1084);
nor U1219 (N_1219,N_1162,N_1082);
and U1220 (N_1220,N_1007,N_1160);
xnor U1221 (N_1221,N_1174,N_1130);
xnor U1222 (N_1222,N_1065,N_1076);
nand U1223 (N_1223,N_1061,N_1164);
xor U1224 (N_1224,N_1086,N_1183);
and U1225 (N_1225,N_1075,N_1027);
nand U1226 (N_1226,N_1132,N_1000);
nor U1227 (N_1227,N_1071,N_1172);
nand U1228 (N_1228,N_1097,N_1050);
nand U1229 (N_1229,N_1072,N_1054);
xnor U1230 (N_1230,N_1073,N_1003);
nor U1231 (N_1231,N_1041,N_1008);
xnor U1232 (N_1232,N_1055,N_1185);
and U1233 (N_1233,N_1153,N_1184);
or U1234 (N_1234,N_1051,N_1175);
nand U1235 (N_1235,N_1166,N_1009);
or U1236 (N_1236,N_1078,N_1062);
and U1237 (N_1237,N_1010,N_1169);
xor U1238 (N_1238,N_1100,N_1070);
and U1239 (N_1239,N_1052,N_1187);
nor U1240 (N_1240,N_1094,N_1049);
and U1241 (N_1241,N_1151,N_1083);
xor U1242 (N_1242,N_1016,N_1170);
nand U1243 (N_1243,N_1135,N_1121);
or U1244 (N_1244,N_1020,N_1063);
or U1245 (N_1245,N_1114,N_1181);
nor U1246 (N_1246,N_1140,N_1154);
or U1247 (N_1247,N_1109,N_1178);
nor U1248 (N_1248,N_1068,N_1157);
or U1249 (N_1249,N_1102,N_1039);
or U1250 (N_1250,N_1098,N_1186);
nor U1251 (N_1251,N_1038,N_1194);
or U1252 (N_1252,N_1066,N_1176);
xor U1253 (N_1253,N_1196,N_1004);
xor U1254 (N_1254,N_1156,N_1113);
xnor U1255 (N_1255,N_1161,N_1031);
or U1256 (N_1256,N_1059,N_1129);
xnor U1257 (N_1257,N_1015,N_1125);
and U1258 (N_1258,N_1037,N_1112);
nand U1259 (N_1259,N_1025,N_1159);
xnor U1260 (N_1260,N_1165,N_1021);
xnor U1261 (N_1261,N_1131,N_1173);
nor U1262 (N_1262,N_1029,N_1189);
or U1263 (N_1263,N_1106,N_1120);
nand U1264 (N_1264,N_1179,N_1056);
xnor U1265 (N_1265,N_1108,N_1057);
nand U1266 (N_1266,N_1133,N_1158);
xnor U1267 (N_1267,N_1006,N_1117);
or U1268 (N_1268,N_1107,N_1069);
xnor U1269 (N_1269,N_1180,N_1011);
or U1270 (N_1270,N_1146,N_1191);
nor U1271 (N_1271,N_1032,N_1023);
and U1272 (N_1272,N_1044,N_1118);
and U1273 (N_1273,N_1019,N_1155);
or U1274 (N_1274,N_1026,N_1012);
or U1275 (N_1275,N_1024,N_1013);
nand U1276 (N_1276,N_1092,N_1077);
and U1277 (N_1277,N_1064,N_1182);
and U1278 (N_1278,N_1144,N_1149);
nor U1279 (N_1279,N_1150,N_1067);
nor U1280 (N_1280,N_1053,N_1022);
xor U1281 (N_1281,N_1148,N_1127);
and U1282 (N_1282,N_1134,N_1081);
and U1283 (N_1283,N_1104,N_1188);
nand U1284 (N_1284,N_1096,N_1033);
nor U1285 (N_1285,N_1030,N_1036);
xnor U1286 (N_1286,N_1045,N_1168);
or U1287 (N_1287,N_1047,N_1103);
nand U1288 (N_1288,N_1177,N_1195);
xnor U1289 (N_1289,N_1122,N_1126);
nor U1290 (N_1290,N_1034,N_1080);
or U1291 (N_1291,N_1141,N_1142);
nor U1292 (N_1292,N_1145,N_1090);
and U1293 (N_1293,N_1074,N_1197);
xnor U1294 (N_1294,N_1115,N_1058);
nand U1295 (N_1295,N_1128,N_1138);
or U1296 (N_1296,N_1095,N_1111);
or U1297 (N_1297,N_1199,N_1171);
or U1298 (N_1298,N_1124,N_1137);
and U1299 (N_1299,N_1152,N_1046);
nor U1300 (N_1300,N_1140,N_1112);
nor U1301 (N_1301,N_1099,N_1067);
xor U1302 (N_1302,N_1182,N_1184);
or U1303 (N_1303,N_1083,N_1149);
or U1304 (N_1304,N_1042,N_1124);
or U1305 (N_1305,N_1079,N_1029);
and U1306 (N_1306,N_1099,N_1038);
and U1307 (N_1307,N_1062,N_1166);
xor U1308 (N_1308,N_1143,N_1196);
and U1309 (N_1309,N_1194,N_1110);
or U1310 (N_1310,N_1093,N_1120);
and U1311 (N_1311,N_1043,N_1013);
xnor U1312 (N_1312,N_1152,N_1072);
or U1313 (N_1313,N_1129,N_1136);
xor U1314 (N_1314,N_1187,N_1119);
or U1315 (N_1315,N_1162,N_1104);
xnor U1316 (N_1316,N_1081,N_1163);
xnor U1317 (N_1317,N_1153,N_1023);
nor U1318 (N_1318,N_1016,N_1002);
nand U1319 (N_1319,N_1163,N_1112);
xnor U1320 (N_1320,N_1094,N_1156);
or U1321 (N_1321,N_1049,N_1160);
nor U1322 (N_1322,N_1085,N_1195);
nor U1323 (N_1323,N_1026,N_1147);
nor U1324 (N_1324,N_1137,N_1182);
xor U1325 (N_1325,N_1013,N_1169);
xnor U1326 (N_1326,N_1125,N_1000);
xor U1327 (N_1327,N_1119,N_1152);
or U1328 (N_1328,N_1175,N_1048);
or U1329 (N_1329,N_1194,N_1075);
nand U1330 (N_1330,N_1126,N_1182);
and U1331 (N_1331,N_1156,N_1074);
or U1332 (N_1332,N_1197,N_1069);
or U1333 (N_1333,N_1130,N_1081);
xnor U1334 (N_1334,N_1159,N_1007);
or U1335 (N_1335,N_1058,N_1094);
and U1336 (N_1336,N_1157,N_1193);
nand U1337 (N_1337,N_1112,N_1040);
nand U1338 (N_1338,N_1190,N_1155);
and U1339 (N_1339,N_1042,N_1046);
or U1340 (N_1340,N_1031,N_1149);
or U1341 (N_1341,N_1076,N_1108);
or U1342 (N_1342,N_1102,N_1060);
and U1343 (N_1343,N_1042,N_1098);
xnor U1344 (N_1344,N_1185,N_1125);
and U1345 (N_1345,N_1130,N_1117);
xnor U1346 (N_1346,N_1035,N_1118);
nor U1347 (N_1347,N_1074,N_1103);
and U1348 (N_1348,N_1087,N_1002);
nand U1349 (N_1349,N_1169,N_1167);
nand U1350 (N_1350,N_1077,N_1082);
nand U1351 (N_1351,N_1176,N_1177);
or U1352 (N_1352,N_1194,N_1018);
nand U1353 (N_1353,N_1137,N_1120);
nor U1354 (N_1354,N_1070,N_1137);
and U1355 (N_1355,N_1156,N_1038);
nor U1356 (N_1356,N_1074,N_1110);
nor U1357 (N_1357,N_1174,N_1147);
and U1358 (N_1358,N_1026,N_1146);
and U1359 (N_1359,N_1041,N_1164);
or U1360 (N_1360,N_1054,N_1067);
or U1361 (N_1361,N_1069,N_1103);
nand U1362 (N_1362,N_1011,N_1063);
nor U1363 (N_1363,N_1166,N_1049);
and U1364 (N_1364,N_1087,N_1161);
nand U1365 (N_1365,N_1108,N_1000);
and U1366 (N_1366,N_1090,N_1112);
xnor U1367 (N_1367,N_1138,N_1083);
and U1368 (N_1368,N_1130,N_1074);
xnor U1369 (N_1369,N_1170,N_1061);
and U1370 (N_1370,N_1150,N_1192);
or U1371 (N_1371,N_1194,N_1189);
xor U1372 (N_1372,N_1027,N_1095);
and U1373 (N_1373,N_1014,N_1076);
and U1374 (N_1374,N_1167,N_1109);
nor U1375 (N_1375,N_1148,N_1170);
nor U1376 (N_1376,N_1000,N_1057);
xor U1377 (N_1377,N_1148,N_1178);
xor U1378 (N_1378,N_1138,N_1170);
or U1379 (N_1379,N_1103,N_1143);
nor U1380 (N_1380,N_1014,N_1166);
nand U1381 (N_1381,N_1178,N_1108);
or U1382 (N_1382,N_1160,N_1191);
nor U1383 (N_1383,N_1012,N_1155);
nand U1384 (N_1384,N_1043,N_1045);
nand U1385 (N_1385,N_1164,N_1193);
xnor U1386 (N_1386,N_1174,N_1153);
or U1387 (N_1387,N_1099,N_1191);
nand U1388 (N_1388,N_1146,N_1172);
nor U1389 (N_1389,N_1128,N_1012);
nand U1390 (N_1390,N_1166,N_1108);
or U1391 (N_1391,N_1186,N_1026);
nor U1392 (N_1392,N_1076,N_1169);
xor U1393 (N_1393,N_1004,N_1185);
nand U1394 (N_1394,N_1060,N_1154);
nand U1395 (N_1395,N_1020,N_1034);
xor U1396 (N_1396,N_1125,N_1191);
nand U1397 (N_1397,N_1029,N_1129);
or U1398 (N_1398,N_1125,N_1082);
or U1399 (N_1399,N_1102,N_1162);
or U1400 (N_1400,N_1328,N_1300);
nor U1401 (N_1401,N_1327,N_1324);
xor U1402 (N_1402,N_1267,N_1313);
nor U1403 (N_1403,N_1240,N_1205);
nand U1404 (N_1404,N_1270,N_1356);
and U1405 (N_1405,N_1298,N_1312);
nand U1406 (N_1406,N_1353,N_1350);
nor U1407 (N_1407,N_1372,N_1385);
nand U1408 (N_1408,N_1293,N_1305);
xnor U1409 (N_1409,N_1303,N_1316);
nand U1410 (N_1410,N_1254,N_1322);
xor U1411 (N_1411,N_1245,N_1359);
or U1412 (N_1412,N_1277,N_1249);
and U1413 (N_1413,N_1225,N_1292);
and U1414 (N_1414,N_1229,N_1250);
nor U1415 (N_1415,N_1258,N_1263);
nor U1416 (N_1416,N_1237,N_1318);
xnor U1417 (N_1417,N_1280,N_1389);
and U1418 (N_1418,N_1275,N_1202);
nand U1419 (N_1419,N_1309,N_1382);
or U1420 (N_1420,N_1379,N_1321);
and U1421 (N_1421,N_1325,N_1252);
or U1422 (N_1422,N_1266,N_1354);
and U1423 (N_1423,N_1374,N_1251);
nand U1424 (N_1424,N_1387,N_1391);
nor U1425 (N_1425,N_1357,N_1208);
nand U1426 (N_1426,N_1299,N_1212);
and U1427 (N_1427,N_1232,N_1295);
nor U1428 (N_1428,N_1209,N_1235);
nand U1429 (N_1429,N_1338,N_1222);
xor U1430 (N_1430,N_1366,N_1219);
nor U1431 (N_1431,N_1296,N_1283);
and U1432 (N_1432,N_1394,N_1220);
xor U1433 (N_1433,N_1213,N_1215);
and U1434 (N_1434,N_1261,N_1247);
or U1435 (N_1435,N_1290,N_1302);
xor U1436 (N_1436,N_1336,N_1314);
or U1437 (N_1437,N_1272,N_1398);
and U1438 (N_1438,N_1268,N_1370);
nor U1439 (N_1439,N_1315,N_1367);
xor U1440 (N_1440,N_1282,N_1386);
xnor U1441 (N_1441,N_1392,N_1349);
nand U1442 (N_1442,N_1226,N_1230);
or U1443 (N_1443,N_1363,N_1294);
or U1444 (N_1444,N_1239,N_1358);
xnor U1445 (N_1445,N_1348,N_1375);
nor U1446 (N_1446,N_1378,N_1393);
xor U1447 (N_1447,N_1264,N_1371);
or U1448 (N_1448,N_1259,N_1326);
nor U1449 (N_1449,N_1238,N_1278);
or U1450 (N_1450,N_1204,N_1364);
nand U1451 (N_1451,N_1216,N_1285);
xor U1452 (N_1452,N_1241,N_1288);
nor U1453 (N_1453,N_1311,N_1373);
or U1454 (N_1454,N_1233,N_1257);
or U1455 (N_1455,N_1210,N_1224);
or U1456 (N_1456,N_1339,N_1360);
xnor U1457 (N_1457,N_1337,N_1397);
and U1458 (N_1458,N_1301,N_1279);
xor U1459 (N_1459,N_1200,N_1203);
xnor U1460 (N_1460,N_1323,N_1376);
or U1461 (N_1461,N_1351,N_1236);
or U1462 (N_1462,N_1377,N_1355);
nor U1463 (N_1463,N_1248,N_1221);
or U1464 (N_1464,N_1380,N_1369);
and U1465 (N_1465,N_1310,N_1262);
or U1466 (N_1466,N_1329,N_1227);
and U1467 (N_1467,N_1214,N_1289);
or U1468 (N_1468,N_1286,N_1399);
and U1469 (N_1469,N_1287,N_1284);
and U1470 (N_1470,N_1304,N_1368);
or U1471 (N_1471,N_1384,N_1343);
nand U1472 (N_1472,N_1217,N_1365);
xnor U1473 (N_1473,N_1345,N_1332);
or U1474 (N_1474,N_1396,N_1390);
nand U1475 (N_1475,N_1260,N_1320);
xnor U1476 (N_1476,N_1234,N_1223);
nand U1477 (N_1477,N_1206,N_1346);
nor U1478 (N_1478,N_1231,N_1342);
nand U1479 (N_1479,N_1273,N_1242);
or U1480 (N_1480,N_1333,N_1347);
nand U1481 (N_1481,N_1253,N_1308);
or U1482 (N_1482,N_1317,N_1362);
xor U1483 (N_1483,N_1243,N_1271);
and U1484 (N_1484,N_1265,N_1341);
or U1485 (N_1485,N_1381,N_1281);
nor U1486 (N_1486,N_1297,N_1361);
xor U1487 (N_1487,N_1269,N_1330);
nor U1488 (N_1488,N_1335,N_1383);
and U1489 (N_1489,N_1307,N_1319);
or U1490 (N_1490,N_1246,N_1276);
and U1491 (N_1491,N_1207,N_1218);
and U1492 (N_1492,N_1395,N_1331);
or U1493 (N_1493,N_1388,N_1274);
or U1494 (N_1494,N_1201,N_1211);
nand U1495 (N_1495,N_1340,N_1344);
nand U1496 (N_1496,N_1256,N_1228);
and U1497 (N_1497,N_1306,N_1255);
nand U1498 (N_1498,N_1352,N_1334);
or U1499 (N_1499,N_1244,N_1291);
nand U1500 (N_1500,N_1328,N_1251);
and U1501 (N_1501,N_1326,N_1323);
or U1502 (N_1502,N_1308,N_1273);
and U1503 (N_1503,N_1308,N_1299);
xnor U1504 (N_1504,N_1396,N_1372);
xnor U1505 (N_1505,N_1275,N_1305);
and U1506 (N_1506,N_1331,N_1317);
nor U1507 (N_1507,N_1271,N_1228);
nand U1508 (N_1508,N_1282,N_1361);
or U1509 (N_1509,N_1203,N_1268);
nor U1510 (N_1510,N_1290,N_1226);
xor U1511 (N_1511,N_1296,N_1232);
xnor U1512 (N_1512,N_1361,N_1296);
nand U1513 (N_1513,N_1378,N_1270);
nor U1514 (N_1514,N_1202,N_1370);
xor U1515 (N_1515,N_1275,N_1303);
and U1516 (N_1516,N_1359,N_1227);
xor U1517 (N_1517,N_1323,N_1329);
nand U1518 (N_1518,N_1313,N_1251);
or U1519 (N_1519,N_1327,N_1387);
or U1520 (N_1520,N_1282,N_1297);
or U1521 (N_1521,N_1377,N_1276);
and U1522 (N_1522,N_1282,N_1360);
or U1523 (N_1523,N_1389,N_1275);
or U1524 (N_1524,N_1292,N_1254);
or U1525 (N_1525,N_1232,N_1231);
nand U1526 (N_1526,N_1296,N_1281);
nor U1527 (N_1527,N_1265,N_1241);
nor U1528 (N_1528,N_1280,N_1349);
or U1529 (N_1529,N_1366,N_1292);
xnor U1530 (N_1530,N_1358,N_1304);
and U1531 (N_1531,N_1396,N_1395);
nand U1532 (N_1532,N_1361,N_1250);
nand U1533 (N_1533,N_1391,N_1212);
nor U1534 (N_1534,N_1284,N_1320);
nand U1535 (N_1535,N_1248,N_1238);
or U1536 (N_1536,N_1254,N_1290);
or U1537 (N_1537,N_1284,N_1347);
nand U1538 (N_1538,N_1276,N_1217);
and U1539 (N_1539,N_1345,N_1202);
nor U1540 (N_1540,N_1285,N_1333);
nor U1541 (N_1541,N_1210,N_1207);
and U1542 (N_1542,N_1357,N_1365);
and U1543 (N_1543,N_1376,N_1205);
xnor U1544 (N_1544,N_1239,N_1374);
and U1545 (N_1545,N_1331,N_1240);
nand U1546 (N_1546,N_1323,N_1391);
nand U1547 (N_1547,N_1385,N_1362);
xor U1548 (N_1548,N_1302,N_1377);
xor U1549 (N_1549,N_1313,N_1341);
nand U1550 (N_1550,N_1258,N_1304);
or U1551 (N_1551,N_1323,N_1324);
xnor U1552 (N_1552,N_1204,N_1330);
nand U1553 (N_1553,N_1328,N_1255);
xnor U1554 (N_1554,N_1201,N_1397);
nor U1555 (N_1555,N_1329,N_1336);
or U1556 (N_1556,N_1322,N_1354);
and U1557 (N_1557,N_1286,N_1252);
nand U1558 (N_1558,N_1360,N_1384);
xor U1559 (N_1559,N_1202,N_1395);
xor U1560 (N_1560,N_1384,N_1216);
nor U1561 (N_1561,N_1233,N_1313);
or U1562 (N_1562,N_1383,N_1205);
and U1563 (N_1563,N_1220,N_1296);
nor U1564 (N_1564,N_1260,N_1365);
and U1565 (N_1565,N_1377,N_1201);
or U1566 (N_1566,N_1356,N_1391);
nand U1567 (N_1567,N_1229,N_1321);
xor U1568 (N_1568,N_1272,N_1379);
nor U1569 (N_1569,N_1359,N_1200);
xnor U1570 (N_1570,N_1213,N_1318);
nand U1571 (N_1571,N_1388,N_1233);
nor U1572 (N_1572,N_1393,N_1283);
nand U1573 (N_1573,N_1207,N_1242);
nor U1574 (N_1574,N_1229,N_1249);
nand U1575 (N_1575,N_1332,N_1324);
nand U1576 (N_1576,N_1393,N_1305);
and U1577 (N_1577,N_1294,N_1345);
nor U1578 (N_1578,N_1219,N_1305);
xor U1579 (N_1579,N_1305,N_1243);
xor U1580 (N_1580,N_1395,N_1267);
nor U1581 (N_1581,N_1302,N_1370);
nor U1582 (N_1582,N_1379,N_1206);
xor U1583 (N_1583,N_1305,N_1354);
nor U1584 (N_1584,N_1316,N_1362);
nand U1585 (N_1585,N_1323,N_1312);
or U1586 (N_1586,N_1243,N_1367);
nand U1587 (N_1587,N_1393,N_1333);
or U1588 (N_1588,N_1388,N_1296);
nand U1589 (N_1589,N_1282,N_1317);
or U1590 (N_1590,N_1347,N_1386);
xor U1591 (N_1591,N_1314,N_1253);
and U1592 (N_1592,N_1317,N_1302);
xor U1593 (N_1593,N_1251,N_1201);
xnor U1594 (N_1594,N_1205,N_1299);
nor U1595 (N_1595,N_1247,N_1204);
or U1596 (N_1596,N_1233,N_1269);
nor U1597 (N_1597,N_1285,N_1231);
and U1598 (N_1598,N_1263,N_1218);
nand U1599 (N_1599,N_1359,N_1235);
xor U1600 (N_1600,N_1415,N_1534);
nor U1601 (N_1601,N_1460,N_1456);
xnor U1602 (N_1602,N_1492,N_1569);
and U1603 (N_1603,N_1462,N_1487);
xor U1604 (N_1604,N_1543,N_1524);
or U1605 (N_1605,N_1437,N_1590);
or U1606 (N_1606,N_1436,N_1575);
nor U1607 (N_1607,N_1435,N_1446);
xnor U1608 (N_1608,N_1461,N_1542);
xor U1609 (N_1609,N_1591,N_1544);
and U1610 (N_1610,N_1523,N_1598);
nand U1611 (N_1611,N_1422,N_1599);
nand U1612 (N_1612,N_1440,N_1494);
or U1613 (N_1613,N_1561,N_1439);
nor U1614 (N_1614,N_1552,N_1597);
and U1615 (N_1615,N_1533,N_1499);
nand U1616 (N_1616,N_1537,N_1486);
xnor U1617 (N_1617,N_1476,N_1589);
nand U1618 (N_1618,N_1596,N_1491);
nor U1619 (N_1619,N_1516,N_1570);
or U1620 (N_1620,N_1459,N_1470);
and U1621 (N_1621,N_1582,N_1554);
nand U1622 (N_1622,N_1424,N_1421);
xnor U1623 (N_1623,N_1485,N_1566);
xor U1624 (N_1624,N_1426,N_1443);
nand U1625 (N_1625,N_1507,N_1584);
nand U1626 (N_1626,N_1528,N_1432);
xor U1627 (N_1627,N_1464,N_1560);
xnor U1628 (N_1628,N_1553,N_1581);
nor U1629 (N_1629,N_1483,N_1402);
and U1630 (N_1630,N_1411,N_1577);
and U1631 (N_1631,N_1510,N_1425);
or U1632 (N_1632,N_1587,N_1466);
nor U1633 (N_1633,N_1509,N_1413);
nand U1634 (N_1634,N_1428,N_1481);
nor U1635 (N_1635,N_1420,N_1520);
nand U1636 (N_1636,N_1595,N_1448);
nor U1637 (N_1637,N_1457,N_1519);
nor U1638 (N_1638,N_1592,N_1530);
and U1639 (N_1639,N_1532,N_1450);
or U1640 (N_1640,N_1430,N_1555);
nor U1641 (N_1641,N_1500,N_1517);
and U1642 (N_1642,N_1564,N_1540);
nand U1643 (N_1643,N_1538,N_1414);
nor U1644 (N_1644,N_1479,N_1452);
and U1645 (N_1645,N_1445,N_1558);
xor U1646 (N_1646,N_1586,N_1493);
and U1647 (N_1647,N_1508,N_1515);
nor U1648 (N_1648,N_1451,N_1573);
xor U1649 (N_1649,N_1511,N_1548);
nor U1650 (N_1650,N_1468,N_1471);
nor U1651 (N_1651,N_1469,N_1531);
and U1652 (N_1652,N_1467,N_1495);
or U1653 (N_1653,N_1423,N_1473);
nor U1654 (N_1654,N_1417,N_1409);
and U1655 (N_1655,N_1477,N_1463);
and U1656 (N_1656,N_1490,N_1489);
nand U1657 (N_1657,N_1505,N_1458);
and U1658 (N_1658,N_1583,N_1449);
and U1659 (N_1659,N_1416,N_1410);
nand U1660 (N_1660,N_1400,N_1518);
or U1661 (N_1661,N_1447,N_1427);
nor U1662 (N_1662,N_1498,N_1551);
xnor U1663 (N_1663,N_1547,N_1567);
nor U1664 (N_1664,N_1585,N_1512);
xnor U1665 (N_1665,N_1568,N_1401);
nand U1666 (N_1666,N_1588,N_1444);
or U1667 (N_1667,N_1442,N_1478);
nand U1668 (N_1668,N_1407,N_1502);
and U1669 (N_1669,N_1521,N_1541);
xnor U1670 (N_1670,N_1431,N_1441);
and U1671 (N_1671,N_1565,N_1539);
nor U1672 (N_1672,N_1506,N_1406);
nand U1673 (N_1673,N_1455,N_1454);
nor U1674 (N_1674,N_1503,N_1412);
nor U1675 (N_1675,N_1572,N_1571);
or U1676 (N_1676,N_1549,N_1497);
or U1677 (N_1677,N_1434,N_1557);
xor U1678 (N_1678,N_1522,N_1580);
and U1679 (N_1679,N_1562,N_1403);
xnor U1680 (N_1680,N_1559,N_1474);
nand U1681 (N_1681,N_1545,N_1438);
nor U1682 (N_1682,N_1496,N_1419);
nand U1683 (N_1683,N_1556,N_1594);
and U1684 (N_1684,N_1484,N_1529);
xnor U1685 (N_1685,N_1404,N_1405);
xnor U1686 (N_1686,N_1504,N_1550);
nor U1687 (N_1687,N_1525,N_1433);
nand U1688 (N_1688,N_1536,N_1408);
xnor U1689 (N_1689,N_1526,N_1527);
and U1690 (N_1690,N_1482,N_1535);
and U1691 (N_1691,N_1453,N_1514);
and U1692 (N_1692,N_1480,N_1501);
and U1693 (N_1693,N_1563,N_1513);
or U1694 (N_1694,N_1465,N_1593);
nand U1695 (N_1695,N_1574,N_1475);
nor U1696 (N_1696,N_1579,N_1488);
and U1697 (N_1697,N_1418,N_1546);
or U1698 (N_1698,N_1578,N_1576);
or U1699 (N_1699,N_1472,N_1429);
nor U1700 (N_1700,N_1544,N_1560);
nand U1701 (N_1701,N_1419,N_1560);
nor U1702 (N_1702,N_1404,N_1482);
and U1703 (N_1703,N_1454,N_1473);
nor U1704 (N_1704,N_1405,N_1461);
or U1705 (N_1705,N_1489,N_1473);
and U1706 (N_1706,N_1549,N_1561);
xor U1707 (N_1707,N_1420,N_1523);
nor U1708 (N_1708,N_1447,N_1444);
nand U1709 (N_1709,N_1489,N_1508);
xnor U1710 (N_1710,N_1527,N_1471);
nor U1711 (N_1711,N_1501,N_1464);
or U1712 (N_1712,N_1454,N_1503);
or U1713 (N_1713,N_1451,N_1540);
and U1714 (N_1714,N_1503,N_1494);
or U1715 (N_1715,N_1420,N_1426);
or U1716 (N_1716,N_1504,N_1406);
xor U1717 (N_1717,N_1576,N_1426);
nor U1718 (N_1718,N_1492,N_1517);
nand U1719 (N_1719,N_1488,N_1457);
or U1720 (N_1720,N_1538,N_1487);
nor U1721 (N_1721,N_1588,N_1426);
nand U1722 (N_1722,N_1518,N_1434);
nand U1723 (N_1723,N_1472,N_1459);
xor U1724 (N_1724,N_1580,N_1573);
and U1725 (N_1725,N_1513,N_1468);
nand U1726 (N_1726,N_1549,N_1542);
and U1727 (N_1727,N_1506,N_1544);
nand U1728 (N_1728,N_1576,N_1477);
or U1729 (N_1729,N_1406,N_1521);
and U1730 (N_1730,N_1405,N_1532);
nand U1731 (N_1731,N_1589,N_1583);
nand U1732 (N_1732,N_1592,N_1414);
or U1733 (N_1733,N_1526,N_1554);
and U1734 (N_1734,N_1450,N_1579);
nor U1735 (N_1735,N_1425,N_1464);
nor U1736 (N_1736,N_1497,N_1524);
xor U1737 (N_1737,N_1409,N_1489);
xor U1738 (N_1738,N_1439,N_1545);
xor U1739 (N_1739,N_1549,N_1530);
xnor U1740 (N_1740,N_1500,N_1526);
xnor U1741 (N_1741,N_1571,N_1452);
nor U1742 (N_1742,N_1466,N_1478);
nand U1743 (N_1743,N_1508,N_1514);
nand U1744 (N_1744,N_1528,N_1521);
nand U1745 (N_1745,N_1599,N_1589);
xor U1746 (N_1746,N_1580,N_1542);
nand U1747 (N_1747,N_1596,N_1451);
xnor U1748 (N_1748,N_1457,N_1455);
xnor U1749 (N_1749,N_1453,N_1406);
nand U1750 (N_1750,N_1411,N_1528);
nor U1751 (N_1751,N_1402,N_1459);
and U1752 (N_1752,N_1477,N_1570);
nand U1753 (N_1753,N_1488,N_1480);
nor U1754 (N_1754,N_1482,N_1425);
or U1755 (N_1755,N_1592,N_1521);
xor U1756 (N_1756,N_1508,N_1422);
nor U1757 (N_1757,N_1544,N_1551);
or U1758 (N_1758,N_1492,N_1541);
nor U1759 (N_1759,N_1410,N_1419);
or U1760 (N_1760,N_1573,N_1417);
nand U1761 (N_1761,N_1430,N_1569);
nor U1762 (N_1762,N_1458,N_1519);
nor U1763 (N_1763,N_1474,N_1593);
nand U1764 (N_1764,N_1521,N_1571);
xor U1765 (N_1765,N_1409,N_1443);
or U1766 (N_1766,N_1461,N_1565);
and U1767 (N_1767,N_1588,N_1437);
or U1768 (N_1768,N_1475,N_1581);
and U1769 (N_1769,N_1434,N_1448);
nor U1770 (N_1770,N_1554,N_1504);
and U1771 (N_1771,N_1480,N_1574);
or U1772 (N_1772,N_1442,N_1569);
nor U1773 (N_1773,N_1462,N_1542);
or U1774 (N_1774,N_1571,N_1547);
or U1775 (N_1775,N_1498,N_1401);
and U1776 (N_1776,N_1533,N_1477);
xnor U1777 (N_1777,N_1453,N_1537);
or U1778 (N_1778,N_1469,N_1433);
nor U1779 (N_1779,N_1545,N_1504);
xnor U1780 (N_1780,N_1530,N_1587);
or U1781 (N_1781,N_1541,N_1557);
nor U1782 (N_1782,N_1483,N_1435);
nand U1783 (N_1783,N_1565,N_1403);
or U1784 (N_1784,N_1503,N_1469);
nand U1785 (N_1785,N_1493,N_1557);
nor U1786 (N_1786,N_1512,N_1539);
and U1787 (N_1787,N_1512,N_1409);
or U1788 (N_1788,N_1497,N_1491);
or U1789 (N_1789,N_1469,N_1499);
nand U1790 (N_1790,N_1591,N_1494);
xor U1791 (N_1791,N_1407,N_1415);
and U1792 (N_1792,N_1462,N_1428);
nor U1793 (N_1793,N_1543,N_1464);
xnor U1794 (N_1794,N_1527,N_1594);
or U1795 (N_1795,N_1530,N_1569);
and U1796 (N_1796,N_1404,N_1558);
and U1797 (N_1797,N_1589,N_1585);
nor U1798 (N_1798,N_1417,N_1450);
and U1799 (N_1799,N_1524,N_1515);
or U1800 (N_1800,N_1778,N_1699);
and U1801 (N_1801,N_1673,N_1654);
nor U1802 (N_1802,N_1723,N_1793);
nor U1803 (N_1803,N_1650,N_1610);
nor U1804 (N_1804,N_1792,N_1718);
nand U1805 (N_1805,N_1720,N_1712);
or U1806 (N_1806,N_1794,N_1668);
or U1807 (N_1807,N_1693,N_1675);
and U1808 (N_1808,N_1714,N_1696);
or U1809 (N_1809,N_1782,N_1708);
xnor U1810 (N_1810,N_1760,N_1613);
or U1811 (N_1811,N_1796,N_1616);
nor U1812 (N_1812,N_1608,N_1715);
or U1813 (N_1813,N_1759,N_1647);
or U1814 (N_1814,N_1659,N_1648);
or U1815 (N_1815,N_1605,N_1651);
nor U1816 (N_1816,N_1698,N_1713);
or U1817 (N_1817,N_1634,N_1627);
and U1818 (N_1818,N_1612,N_1685);
xor U1819 (N_1819,N_1756,N_1764);
or U1820 (N_1820,N_1641,N_1609);
xnor U1821 (N_1821,N_1640,N_1744);
nor U1822 (N_1822,N_1623,N_1680);
nand U1823 (N_1823,N_1674,N_1746);
and U1824 (N_1824,N_1692,N_1797);
nor U1825 (N_1825,N_1777,N_1730);
nor U1826 (N_1826,N_1615,N_1652);
or U1827 (N_1827,N_1733,N_1672);
and U1828 (N_1828,N_1681,N_1774);
nor U1829 (N_1829,N_1656,N_1717);
nand U1830 (N_1830,N_1614,N_1761);
nand U1831 (N_1831,N_1742,N_1706);
xnor U1832 (N_1832,N_1791,N_1687);
xnor U1833 (N_1833,N_1664,N_1737);
xnor U1834 (N_1834,N_1728,N_1618);
nor U1835 (N_1835,N_1683,N_1787);
and U1836 (N_1836,N_1768,N_1762);
or U1837 (N_1837,N_1653,N_1619);
or U1838 (N_1838,N_1789,N_1725);
xnor U1839 (N_1839,N_1646,N_1741);
nor U1840 (N_1840,N_1748,N_1738);
and U1841 (N_1841,N_1790,N_1663);
xor U1842 (N_1842,N_1766,N_1783);
nand U1843 (N_1843,N_1604,N_1719);
nand U1844 (N_1844,N_1637,N_1765);
nand U1845 (N_1845,N_1669,N_1658);
or U1846 (N_1846,N_1779,N_1731);
nor U1847 (N_1847,N_1703,N_1670);
and U1848 (N_1848,N_1657,N_1622);
or U1849 (N_1849,N_1769,N_1620);
nand U1850 (N_1850,N_1773,N_1788);
xor U1851 (N_1851,N_1727,N_1607);
or U1852 (N_1852,N_1666,N_1721);
xnor U1853 (N_1853,N_1753,N_1763);
nand U1854 (N_1854,N_1690,N_1635);
nand U1855 (N_1855,N_1661,N_1624);
nor U1856 (N_1856,N_1688,N_1636);
and U1857 (N_1857,N_1707,N_1691);
xnor U1858 (N_1858,N_1735,N_1722);
and U1859 (N_1859,N_1677,N_1705);
nor U1860 (N_1860,N_1785,N_1770);
nor U1861 (N_1861,N_1625,N_1655);
nor U1862 (N_1862,N_1602,N_1600);
nor U1863 (N_1863,N_1642,N_1665);
nor U1864 (N_1864,N_1694,N_1617);
xor U1865 (N_1865,N_1724,N_1786);
and U1866 (N_1866,N_1601,N_1775);
and U1867 (N_1867,N_1784,N_1678);
or U1868 (N_1868,N_1795,N_1684);
and U1869 (N_1869,N_1649,N_1732);
nor U1870 (N_1870,N_1743,N_1754);
nor U1871 (N_1871,N_1697,N_1639);
and U1872 (N_1872,N_1729,N_1716);
or U1873 (N_1873,N_1630,N_1799);
nand U1874 (N_1874,N_1633,N_1701);
nor U1875 (N_1875,N_1662,N_1780);
nand U1876 (N_1876,N_1676,N_1745);
xor U1877 (N_1877,N_1734,N_1645);
nor U1878 (N_1878,N_1772,N_1758);
nor U1879 (N_1879,N_1626,N_1689);
or U1880 (N_1880,N_1781,N_1767);
nor U1881 (N_1881,N_1747,N_1644);
xor U1882 (N_1882,N_1638,N_1632);
nor U1883 (N_1883,N_1771,N_1629);
or U1884 (N_1884,N_1776,N_1757);
and U1885 (N_1885,N_1749,N_1710);
and U1886 (N_1886,N_1679,N_1686);
nor U1887 (N_1887,N_1739,N_1740);
and U1888 (N_1888,N_1711,N_1660);
or U1889 (N_1889,N_1682,N_1798);
nor U1890 (N_1890,N_1755,N_1671);
nor U1891 (N_1891,N_1709,N_1667);
nand U1892 (N_1892,N_1752,N_1695);
and U1893 (N_1893,N_1611,N_1606);
and U1894 (N_1894,N_1628,N_1702);
xnor U1895 (N_1895,N_1726,N_1603);
and U1896 (N_1896,N_1621,N_1631);
xnor U1897 (N_1897,N_1751,N_1700);
or U1898 (N_1898,N_1736,N_1643);
and U1899 (N_1899,N_1750,N_1704);
and U1900 (N_1900,N_1750,N_1724);
xor U1901 (N_1901,N_1675,N_1697);
or U1902 (N_1902,N_1679,N_1799);
xor U1903 (N_1903,N_1687,N_1752);
nor U1904 (N_1904,N_1601,N_1627);
and U1905 (N_1905,N_1755,N_1645);
xor U1906 (N_1906,N_1785,N_1679);
nor U1907 (N_1907,N_1746,N_1658);
nor U1908 (N_1908,N_1703,N_1743);
nor U1909 (N_1909,N_1625,N_1740);
nor U1910 (N_1910,N_1698,N_1783);
nand U1911 (N_1911,N_1664,N_1721);
and U1912 (N_1912,N_1694,N_1786);
or U1913 (N_1913,N_1734,N_1751);
or U1914 (N_1914,N_1632,N_1727);
xnor U1915 (N_1915,N_1616,N_1703);
or U1916 (N_1916,N_1602,N_1782);
or U1917 (N_1917,N_1610,N_1626);
xnor U1918 (N_1918,N_1639,N_1728);
nand U1919 (N_1919,N_1713,N_1636);
nand U1920 (N_1920,N_1796,N_1658);
and U1921 (N_1921,N_1673,N_1645);
or U1922 (N_1922,N_1791,N_1788);
nand U1923 (N_1923,N_1612,N_1762);
xnor U1924 (N_1924,N_1786,N_1616);
nor U1925 (N_1925,N_1791,N_1724);
or U1926 (N_1926,N_1602,N_1648);
and U1927 (N_1927,N_1688,N_1722);
and U1928 (N_1928,N_1730,N_1736);
nor U1929 (N_1929,N_1766,N_1773);
or U1930 (N_1930,N_1686,N_1730);
and U1931 (N_1931,N_1774,N_1640);
nand U1932 (N_1932,N_1781,N_1778);
nor U1933 (N_1933,N_1634,N_1684);
nor U1934 (N_1934,N_1741,N_1706);
and U1935 (N_1935,N_1740,N_1646);
or U1936 (N_1936,N_1765,N_1749);
or U1937 (N_1937,N_1612,N_1711);
nor U1938 (N_1938,N_1715,N_1799);
and U1939 (N_1939,N_1628,N_1782);
xor U1940 (N_1940,N_1769,N_1797);
or U1941 (N_1941,N_1618,N_1664);
nor U1942 (N_1942,N_1726,N_1666);
nand U1943 (N_1943,N_1724,N_1709);
or U1944 (N_1944,N_1625,N_1676);
xnor U1945 (N_1945,N_1778,N_1608);
and U1946 (N_1946,N_1688,N_1604);
nor U1947 (N_1947,N_1601,N_1698);
and U1948 (N_1948,N_1679,N_1655);
xnor U1949 (N_1949,N_1665,N_1779);
xor U1950 (N_1950,N_1630,N_1693);
and U1951 (N_1951,N_1659,N_1785);
nor U1952 (N_1952,N_1760,N_1604);
nor U1953 (N_1953,N_1607,N_1725);
and U1954 (N_1954,N_1641,N_1784);
nor U1955 (N_1955,N_1752,N_1648);
nand U1956 (N_1956,N_1773,N_1607);
or U1957 (N_1957,N_1786,N_1635);
and U1958 (N_1958,N_1796,N_1604);
or U1959 (N_1959,N_1708,N_1648);
nor U1960 (N_1960,N_1759,N_1673);
nor U1961 (N_1961,N_1703,N_1729);
nor U1962 (N_1962,N_1798,N_1694);
nand U1963 (N_1963,N_1601,N_1690);
or U1964 (N_1964,N_1755,N_1641);
nand U1965 (N_1965,N_1631,N_1770);
and U1966 (N_1966,N_1744,N_1757);
or U1967 (N_1967,N_1727,N_1634);
nor U1968 (N_1968,N_1679,N_1755);
and U1969 (N_1969,N_1630,N_1764);
nand U1970 (N_1970,N_1623,N_1780);
nor U1971 (N_1971,N_1686,N_1692);
and U1972 (N_1972,N_1678,N_1679);
nand U1973 (N_1973,N_1720,N_1792);
nand U1974 (N_1974,N_1672,N_1617);
or U1975 (N_1975,N_1755,N_1789);
xnor U1976 (N_1976,N_1601,N_1663);
or U1977 (N_1977,N_1736,N_1756);
xor U1978 (N_1978,N_1734,N_1799);
nor U1979 (N_1979,N_1667,N_1760);
or U1980 (N_1980,N_1742,N_1674);
or U1981 (N_1981,N_1656,N_1704);
xnor U1982 (N_1982,N_1754,N_1667);
or U1983 (N_1983,N_1614,N_1685);
xnor U1984 (N_1984,N_1745,N_1719);
nand U1985 (N_1985,N_1637,N_1763);
or U1986 (N_1986,N_1676,N_1752);
nand U1987 (N_1987,N_1703,N_1750);
nor U1988 (N_1988,N_1751,N_1752);
xor U1989 (N_1989,N_1717,N_1693);
nor U1990 (N_1990,N_1653,N_1623);
nand U1991 (N_1991,N_1740,N_1743);
nand U1992 (N_1992,N_1774,N_1747);
nand U1993 (N_1993,N_1795,N_1762);
xor U1994 (N_1994,N_1671,N_1712);
xnor U1995 (N_1995,N_1788,N_1678);
nor U1996 (N_1996,N_1788,N_1701);
nand U1997 (N_1997,N_1754,N_1671);
or U1998 (N_1998,N_1650,N_1798);
nor U1999 (N_1999,N_1701,N_1659);
nand U2000 (N_2000,N_1913,N_1932);
and U2001 (N_2001,N_1842,N_1960);
and U2002 (N_2002,N_1945,N_1867);
or U2003 (N_2003,N_1880,N_1897);
nand U2004 (N_2004,N_1895,N_1820);
nor U2005 (N_2005,N_1924,N_1969);
and U2006 (N_2006,N_1978,N_1966);
or U2007 (N_2007,N_1826,N_1912);
or U2008 (N_2008,N_1935,N_1955);
and U2009 (N_2009,N_1837,N_1828);
nor U2010 (N_2010,N_1954,N_1900);
or U2011 (N_2011,N_1878,N_1958);
and U2012 (N_2012,N_1870,N_1965);
nor U2013 (N_2013,N_1940,N_1967);
and U2014 (N_2014,N_1996,N_1810);
or U2015 (N_2015,N_1861,N_1865);
xor U2016 (N_2016,N_1929,N_1835);
or U2017 (N_2017,N_1852,N_1931);
or U2018 (N_2018,N_1845,N_1890);
nand U2019 (N_2019,N_1823,N_1882);
and U2020 (N_2020,N_1893,N_1812);
nor U2021 (N_2021,N_1829,N_1903);
or U2022 (N_2022,N_1862,N_1858);
and U2023 (N_2023,N_1983,N_1970);
or U2024 (N_2024,N_1991,N_1839);
or U2025 (N_2025,N_1821,N_1989);
or U2026 (N_2026,N_1941,N_1951);
or U2027 (N_2027,N_1961,N_1864);
and U2028 (N_2028,N_1918,N_1926);
and U2029 (N_2029,N_1928,N_1899);
and U2030 (N_2030,N_1849,N_1855);
or U2031 (N_2031,N_1942,N_1898);
nand U2032 (N_2032,N_1840,N_1847);
or U2033 (N_2033,N_1885,N_1988);
nand U2034 (N_2034,N_1914,N_1871);
nand U2035 (N_2035,N_1892,N_1806);
nor U2036 (N_2036,N_1923,N_1987);
nor U2037 (N_2037,N_1868,N_1805);
xor U2038 (N_2038,N_1943,N_1836);
or U2039 (N_2039,N_1887,N_1971);
and U2040 (N_2040,N_1911,N_1869);
xnor U2041 (N_2041,N_1877,N_1891);
or U2042 (N_2042,N_1848,N_1956);
nor U2043 (N_2043,N_1815,N_1997);
or U2044 (N_2044,N_1982,N_1909);
xor U2045 (N_2045,N_1896,N_1916);
nand U2046 (N_2046,N_1857,N_1832);
nand U2047 (N_2047,N_1936,N_1894);
xnor U2048 (N_2048,N_1811,N_1949);
nand U2049 (N_2049,N_1854,N_1994);
and U2050 (N_2050,N_1904,N_1992);
or U2051 (N_2051,N_1937,N_1803);
nand U2052 (N_2052,N_1883,N_1860);
xnor U2053 (N_2053,N_1843,N_1950);
and U2054 (N_2054,N_1827,N_1998);
nand U2055 (N_2055,N_1984,N_1925);
xnor U2056 (N_2056,N_1999,N_1963);
nor U2057 (N_2057,N_1920,N_1800);
xor U2058 (N_2058,N_1946,N_1830);
xor U2059 (N_2059,N_1927,N_1974);
and U2060 (N_2060,N_1939,N_1986);
nand U2061 (N_2061,N_1853,N_1816);
and U2062 (N_2062,N_1844,N_1850);
nand U2063 (N_2063,N_1980,N_1952);
nor U2064 (N_2064,N_1834,N_1804);
nand U2065 (N_2065,N_1873,N_1995);
xnor U2066 (N_2066,N_1964,N_1917);
or U2067 (N_2067,N_1808,N_1851);
nand U2068 (N_2068,N_1863,N_1957);
or U2069 (N_2069,N_1976,N_1933);
nand U2070 (N_2070,N_1874,N_1807);
nor U2071 (N_2071,N_1977,N_1975);
xnor U2072 (N_2072,N_1901,N_1902);
or U2073 (N_2073,N_1915,N_1825);
nor U2074 (N_2074,N_1802,N_1872);
and U2075 (N_2075,N_1824,N_1884);
and U2076 (N_2076,N_1968,N_1906);
xor U2077 (N_2077,N_1889,N_1841);
nor U2078 (N_2078,N_1934,N_1938);
nand U2079 (N_2079,N_1993,N_1990);
nand U2080 (N_2080,N_1822,N_1985);
nand U2081 (N_2081,N_1818,N_1981);
nand U2082 (N_2082,N_1886,N_1846);
nor U2083 (N_2083,N_1876,N_1908);
xnor U2084 (N_2084,N_1859,N_1881);
nor U2085 (N_2085,N_1831,N_1819);
or U2086 (N_2086,N_1919,N_1962);
nand U2087 (N_2087,N_1801,N_1907);
nor U2088 (N_2088,N_1922,N_1905);
nor U2089 (N_2089,N_1814,N_1959);
xor U2090 (N_2090,N_1944,N_1973);
or U2091 (N_2091,N_1888,N_1947);
xor U2092 (N_2092,N_1972,N_1948);
and U2093 (N_2093,N_1809,N_1813);
or U2094 (N_2094,N_1921,N_1875);
xnor U2095 (N_2095,N_1953,N_1833);
nand U2096 (N_2096,N_1838,N_1866);
nand U2097 (N_2097,N_1930,N_1879);
and U2098 (N_2098,N_1910,N_1817);
nor U2099 (N_2099,N_1979,N_1856);
xor U2100 (N_2100,N_1801,N_1863);
xnor U2101 (N_2101,N_1945,N_1936);
nand U2102 (N_2102,N_1868,N_1806);
nor U2103 (N_2103,N_1913,N_1859);
xnor U2104 (N_2104,N_1856,N_1847);
or U2105 (N_2105,N_1940,N_1959);
or U2106 (N_2106,N_1826,N_1846);
xnor U2107 (N_2107,N_1875,N_1971);
or U2108 (N_2108,N_1854,N_1990);
nor U2109 (N_2109,N_1980,N_1873);
nand U2110 (N_2110,N_1976,N_1816);
nor U2111 (N_2111,N_1923,N_1848);
or U2112 (N_2112,N_1930,N_1857);
and U2113 (N_2113,N_1885,N_1827);
or U2114 (N_2114,N_1913,N_1836);
nor U2115 (N_2115,N_1802,N_1828);
xnor U2116 (N_2116,N_1860,N_1870);
or U2117 (N_2117,N_1812,N_1894);
or U2118 (N_2118,N_1913,N_1891);
and U2119 (N_2119,N_1978,N_1934);
nor U2120 (N_2120,N_1805,N_1817);
xor U2121 (N_2121,N_1878,N_1969);
or U2122 (N_2122,N_1940,N_1890);
nor U2123 (N_2123,N_1985,N_1823);
or U2124 (N_2124,N_1840,N_1819);
nand U2125 (N_2125,N_1835,N_1844);
nor U2126 (N_2126,N_1904,N_1909);
xor U2127 (N_2127,N_1876,N_1922);
or U2128 (N_2128,N_1832,N_1840);
xor U2129 (N_2129,N_1955,N_1834);
nor U2130 (N_2130,N_1839,N_1985);
nand U2131 (N_2131,N_1970,N_1806);
and U2132 (N_2132,N_1943,N_1942);
nor U2133 (N_2133,N_1800,N_1832);
xnor U2134 (N_2134,N_1944,N_1837);
nand U2135 (N_2135,N_1942,N_1968);
or U2136 (N_2136,N_1892,N_1945);
nor U2137 (N_2137,N_1928,N_1835);
nor U2138 (N_2138,N_1843,N_1813);
xor U2139 (N_2139,N_1901,N_1868);
xor U2140 (N_2140,N_1923,N_1847);
and U2141 (N_2141,N_1895,N_1975);
nor U2142 (N_2142,N_1999,N_1980);
or U2143 (N_2143,N_1986,N_1888);
nand U2144 (N_2144,N_1800,N_1884);
xnor U2145 (N_2145,N_1952,N_1937);
xnor U2146 (N_2146,N_1900,N_1862);
and U2147 (N_2147,N_1804,N_1951);
nor U2148 (N_2148,N_1979,N_1950);
and U2149 (N_2149,N_1836,N_1984);
nor U2150 (N_2150,N_1928,N_1960);
nand U2151 (N_2151,N_1938,N_1992);
or U2152 (N_2152,N_1850,N_1837);
or U2153 (N_2153,N_1941,N_1958);
xor U2154 (N_2154,N_1839,N_1934);
nand U2155 (N_2155,N_1898,N_1944);
xor U2156 (N_2156,N_1871,N_1874);
or U2157 (N_2157,N_1813,N_1869);
and U2158 (N_2158,N_1929,N_1926);
xnor U2159 (N_2159,N_1816,N_1842);
nand U2160 (N_2160,N_1857,N_1879);
and U2161 (N_2161,N_1966,N_1813);
and U2162 (N_2162,N_1854,N_1967);
and U2163 (N_2163,N_1985,N_1820);
or U2164 (N_2164,N_1878,N_1803);
xnor U2165 (N_2165,N_1939,N_1971);
and U2166 (N_2166,N_1963,N_1941);
nand U2167 (N_2167,N_1867,N_1892);
or U2168 (N_2168,N_1820,N_1938);
and U2169 (N_2169,N_1850,N_1956);
nand U2170 (N_2170,N_1929,N_1902);
or U2171 (N_2171,N_1839,N_1996);
and U2172 (N_2172,N_1936,N_1988);
and U2173 (N_2173,N_1868,N_1918);
nor U2174 (N_2174,N_1808,N_1886);
xnor U2175 (N_2175,N_1975,N_1832);
nor U2176 (N_2176,N_1932,N_1802);
nor U2177 (N_2177,N_1829,N_1957);
xnor U2178 (N_2178,N_1930,N_1849);
and U2179 (N_2179,N_1892,N_1854);
nor U2180 (N_2180,N_1863,N_1839);
and U2181 (N_2181,N_1920,N_1861);
or U2182 (N_2182,N_1989,N_1995);
and U2183 (N_2183,N_1822,N_1885);
nand U2184 (N_2184,N_1807,N_1875);
nor U2185 (N_2185,N_1940,N_1996);
or U2186 (N_2186,N_1897,N_1816);
nor U2187 (N_2187,N_1920,N_1895);
or U2188 (N_2188,N_1936,N_1975);
nor U2189 (N_2189,N_1895,N_1952);
nand U2190 (N_2190,N_1854,N_1909);
and U2191 (N_2191,N_1837,N_1978);
or U2192 (N_2192,N_1816,N_1867);
nand U2193 (N_2193,N_1805,N_1815);
nor U2194 (N_2194,N_1822,N_1873);
nor U2195 (N_2195,N_1879,N_1945);
xnor U2196 (N_2196,N_1834,N_1845);
xnor U2197 (N_2197,N_1983,N_1956);
xnor U2198 (N_2198,N_1806,N_1836);
nand U2199 (N_2199,N_1902,N_1875);
nand U2200 (N_2200,N_2083,N_2031);
nand U2201 (N_2201,N_2171,N_2142);
or U2202 (N_2202,N_2094,N_2101);
nor U2203 (N_2203,N_2067,N_2127);
nor U2204 (N_2204,N_2059,N_2087);
xnor U2205 (N_2205,N_2074,N_2140);
xnor U2206 (N_2206,N_2118,N_2153);
xnor U2207 (N_2207,N_2050,N_2058);
nor U2208 (N_2208,N_2183,N_2145);
or U2209 (N_2209,N_2052,N_2103);
and U2210 (N_2210,N_2150,N_2049);
nand U2211 (N_2211,N_2048,N_2016);
or U2212 (N_2212,N_2198,N_2028);
or U2213 (N_2213,N_2141,N_2129);
and U2214 (N_2214,N_2014,N_2023);
xnor U2215 (N_2215,N_2071,N_2089);
and U2216 (N_2216,N_2199,N_2196);
and U2217 (N_2217,N_2166,N_2197);
nor U2218 (N_2218,N_2072,N_2119);
nor U2219 (N_2219,N_2175,N_2109);
nor U2220 (N_2220,N_2027,N_2161);
nor U2221 (N_2221,N_2130,N_2047);
or U2222 (N_2222,N_2054,N_2181);
xor U2223 (N_2223,N_2068,N_2173);
or U2224 (N_2224,N_2154,N_2172);
or U2225 (N_2225,N_2004,N_2105);
nand U2226 (N_2226,N_2156,N_2164);
nand U2227 (N_2227,N_2106,N_2104);
nand U2228 (N_2228,N_2082,N_2099);
or U2229 (N_2229,N_2045,N_2177);
and U2230 (N_2230,N_2081,N_2152);
nor U2231 (N_2231,N_2147,N_2114);
and U2232 (N_2232,N_2026,N_2003);
and U2233 (N_2233,N_2034,N_2182);
and U2234 (N_2234,N_2139,N_2123);
xnor U2235 (N_2235,N_2008,N_2036);
nand U2236 (N_2236,N_2030,N_2192);
nor U2237 (N_2237,N_2079,N_2057);
xor U2238 (N_2238,N_2029,N_2005);
xor U2239 (N_2239,N_2124,N_2013);
and U2240 (N_2240,N_2085,N_2137);
xnor U2241 (N_2241,N_2033,N_2159);
nor U2242 (N_2242,N_2095,N_2151);
xor U2243 (N_2243,N_2162,N_2160);
and U2244 (N_2244,N_2138,N_2111);
nor U2245 (N_2245,N_2126,N_2170);
nand U2246 (N_2246,N_2148,N_2186);
and U2247 (N_2247,N_2179,N_2097);
or U2248 (N_2248,N_2012,N_2178);
nor U2249 (N_2249,N_2102,N_2060);
xnor U2250 (N_2250,N_2121,N_2132);
nor U2251 (N_2251,N_2163,N_2017);
and U2252 (N_2252,N_2006,N_2146);
nor U2253 (N_2253,N_2195,N_2010);
and U2254 (N_2254,N_2168,N_2035);
and U2255 (N_2255,N_2053,N_2041);
nor U2256 (N_2256,N_2077,N_2158);
and U2257 (N_2257,N_2064,N_2125);
nor U2258 (N_2258,N_2143,N_2063);
nand U2259 (N_2259,N_2002,N_2176);
xnor U2260 (N_2260,N_2075,N_2021);
xor U2261 (N_2261,N_2009,N_2133);
xnor U2262 (N_2262,N_2084,N_2062);
nand U2263 (N_2263,N_2135,N_2011);
or U2264 (N_2264,N_2190,N_2113);
nor U2265 (N_2265,N_2073,N_2065);
or U2266 (N_2266,N_2107,N_2024);
nor U2267 (N_2267,N_2020,N_2191);
nor U2268 (N_2268,N_2018,N_2076);
nand U2269 (N_2269,N_2001,N_2185);
or U2270 (N_2270,N_2116,N_2066);
nor U2271 (N_2271,N_2043,N_2007);
or U2272 (N_2272,N_2110,N_2044);
or U2273 (N_2273,N_2037,N_2056);
nor U2274 (N_2274,N_2108,N_2167);
nand U2275 (N_2275,N_2080,N_2100);
xnor U2276 (N_2276,N_2165,N_2122);
nand U2277 (N_2277,N_2098,N_2038);
and U2278 (N_2278,N_2019,N_2180);
nor U2279 (N_2279,N_2040,N_2078);
and U2280 (N_2280,N_2144,N_2069);
nand U2281 (N_2281,N_2025,N_2032);
xor U2282 (N_2282,N_2136,N_2188);
xnor U2283 (N_2283,N_2015,N_2134);
xor U2284 (N_2284,N_2194,N_2187);
or U2285 (N_2285,N_2051,N_2022);
nand U2286 (N_2286,N_2184,N_2091);
xor U2287 (N_2287,N_2117,N_2169);
and U2288 (N_2288,N_2046,N_2174);
xnor U2289 (N_2289,N_2131,N_2092);
nand U2290 (N_2290,N_2193,N_2086);
xor U2291 (N_2291,N_2149,N_2090);
or U2292 (N_2292,N_2042,N_2157);
and U2293 (N_2293,N_2128,N_2115);
and U2294 (N_2294,N_2070,N_2112);
xor U2295 (N_2295,N_2088,N_2093);
nand U2296 (N_2296,N_2096,N_2000);
nor U2297 (N_2297,N_2055,N_2120);
or U2298 (N_2298,N_2039,N_2155);
nor U2299 (N_2299,N_2189,N_2061);
nand U2300 (N_2300,N_2166,N_2108);
xor U2301 (N_2301,N_2174,N_2017);
xor U2302 (N_2302,N_2097,N_2108);
nand U2303 (N_2303,N_2177,N_2035);
nor U2304 (N_2304,N_2057,N_2108);
or U2305 (N_2305,N_2010,N_2087);
or U2306 (N_2306,N_2032,N_2117);
xnor U2307 (N_2307,N_2040,N_2198);
and U2308 (N_2308,N_2186,N_2022);
nor U2309 (N_2309,N_2039,N_2095);
and U2310 (N_2310,N_2076,N_2106);
nor U2311 (N_2311,N_2074,N_2179);
nand U2312 (N_2312,N_2141,N_2099);
xnor U2313 (N_2313,N_2144,N_2148);
nor U2314 (N_2314,N_2196,N_2109);
or U2315 (N_2315,N_2068,N_2191);
or U2316 (N_2316,N_2121,N_2147);
nor U2317 (N_2317,N_2165,N_2151);
xor U2318 (N_2318,N_2012,N_2161);
or U2319 (N_2319,N_2037,N_2116);
or U2320 (N_2320,N_2178,N_2096);
or U2321 (N_2321,N_2132,N_2176);
nor U2322 (N_2322,N_2069,N_2055);
or U2323 (N_2323,N_2049,N_2076);
nand U2324 (N_2324,N_2070,N_2188);
nor U2325 (N_2325,N_2003,N_2162);
xnor U2326 (N_2326,N_2194,N_2048);
nand U2327 (N_2327,N_2094,N_2078);
nand U2328 (N_2328,N_2150,N_2183);
xor U2329 (N_2329,N_2175,N_2162);
xnor U2330 (N_2330,N_2063,N_2040);
or U2331 (N_2331,N_2131,N_2027);
and U2332 (N_2332,N_2148,N_2074);
and U2333 (N_2333,N_2020,N_2098);
and U2334 (N_2334,N_2146,N_2043);
and U2335 (N_2335,N_2050,N_2166);
nand U2336 (N_2336,N_2168,N_2132);
nor U2337 (N_2337,N_2062,N_2173);
and U2338 (N_2338,N_2166,N_2161);
xnor U2339 (N_2339,N_2105,N_2064);
xor U2340 (N_2340,N_2028,N_2164);
nor U2341 (N_2341,N_2178,N_2153);
or U2342 (N_2342,N_2145,N_2008);
xnor U2343 (N_2343,N_2037,N_2101);
or U2344 (N_2344,N_2121,N_2128);
nand U2345 (N_2345,N_2174,N_2161);
xnor U2346 (N_2346,N_2039,N_2189);
or U2347 (N_2347,N_2063,N_2002);
or U2348 (N_2348,N_2124,N_2151);
or U2349 (N_2349,N_2011,N_2104);
or U2350 (N_2350,N_2002,N_2160);
or U2351 (N_2351,N_2060,N_2069);
nand U2352 (N_2352,N_2032,N_2152);
nor U2353 (N_2353,N_2178,N_2145);
nor U2354 (N_2354,N_2172,N_2096);
xor U2355 (N_2355,N_2103,N_2185);
nor U2356 (N_2356,N_2198,N_2107);
nor U2357 (N_2357,N_2011,N_2009);
nor U2358 (N_2358,N_2141,N_2059);
or U2359 (N_2359,N_2006,N_2101);
or U2360 (N_2360,N_2041,N_2097);
and U2361 (N_2361,N_2011,N_2117);
nand U2362 (N_2362,N_2185,N_2015);
nand U2363 (N_2363,N_2055,N_2068);
nand U2364 (N_2364,N_2042,N_2030);
or U2365 (N_2365,N_2041,N_2082);
nand U2366 (N_2366,N_2104,N_2043);
and U2367 (N_2367,N_2098,N_2109);
or U2368 (N_2368,N_2177,N_2049);
nand U2369 (N_2369,N_2022,N_2188);
nor U2370 (N_2370,N_2189,N_2154);
nor U2371 (N_2371,N_2068,N_2131);
xnor U2372 (N_2372,N_2006,N_2032);
xnor U2373 (N_2373,N_2164,N_2035);
xor U2374 (N_2374,N_2102,N_2094);
or U2375 (N_2375,N_2065,N_2068);
nand U2376 (N_2376,N_2064,N_2075);
or U2377 (N_2377,N_2040,N_2085);
or U2378 (N_2378,N_2151,N_2047);
nand U2379 (N_2379,N_2030,N_2059);
nor U2380 (N_2380,N_2134,N_2099);
and U2381 (N_2381,N_2166,N_2115);
or U2382 (N_2382,N_2145,N_2034);
and U2383 (N_2383,N_2050,N_2077);
nor U2384 (N_2384,N_2107,N_2018);
xor U2385 (N_2385,N_2105,N_2089);
or U2386 (N_2386,N_2088,N_2000);
xnor U2387 (N_2387,N_2145,N_2096);
nor U2388 (N_2388,N_2176,N_2116);
nor U2389 (N_2389,N_2029,N_2135);
nor U2390 (N_2390,N_2194,N_2088);
nand U2391 (N_2391,N_2049,N_2016);
and U2392 (N_2392,N_2094,N_2124);
nand U2393 (N_2393,N_2185,N_2161);
and U2394 (N_2394,N_2111,N_2070);
nor U2395 (N_2395,N_2015,N_2068);
nor U2396 (N_2396,N_2199,N_2075);
and U2397 (N_2397,N_2097,N_2075);
or U2398 (N_2398,N_2171,N_2025);
or U2399 (N_2399,N_2091,N_2097);
nand U2400 (N_2400,N_2285,N_2210);
and U2401 (N_2401,N_2383,N_2351);
and U2402 (N_2402,N_2221,N_2263);
nand U2403 (N_2403,N_2363,N_2374);
nor U2404 (N_2404,N_2229,N_2271);
xor U2405 (N_2405,N_2218,N_2333);
and U2406 (N_2406,N_2284,N_2370);
xnor U2407 (N_2407,N_2272,N_2328);
xor U2408 (N_2408,N_2340,N_2323);
nor U2409 (N_2409,N_2364,N_2329);
and U2410 (N_2410,N_2317,N_2341);
nor U2411 (N_2411,N_2399,N_2280);
and U2412 (N_2412,N_2278,N_2264);
xnor U2413 (N_2413,N_2287,N_2299);
or U2414 (N_2414,N_2262,N_2313);
nand U2415 (N_2415,N_2297,N_2352);
nand U2416 (N_2416,N_2378,N_2225);
and U2417 (N_2417,N_2224,N_2350);
or U2418 (N_2418,N_2296,N_2345);
and U2419 (N_2419,N_2355,N_2222);
or U2420 (N_2420,N_2200,N_2311);
nor U2421 (N_2421,N_2377,N_2281);
and U2422 (N_2422,N_2246,N_2301);
and U2423 (N_2423,N_2213,N_2368);
or U2424 (N_2424,N_2273,N_2236);
and U2425 (N_2425,N_2392,N_2255);
nand U2426 (N_2426,N_2387,N_2336);
nor U2427 (N_2427,N_2361,N_2390);
xor U2428 (N_2428,N_2310,N_2293);
nand U2429 (N_2429,N_2233,N_2360);
or U2430 (N_2430,N_2204,N_2248);
or U2431 (N_2431,N_2217,N_2291);
xor U2432 (N_2432,N_2395,N_2302);
nand U2433 (N_2433,N_2373,N_2325);
nand U2434 (N_2434,N_2295,N_2207);
or U2435 (N_2435,N_2226,N_2257);
xnor U2436 (N_2436,N_2259,N_2211);
nor U2437 (N_2437,N_2309,N_2234);
nor U2438 (N_2438,N_2335,N_2300);
nand U2439 (N_2439,N_2240,N_2356);
nand U2440 (N_2440,N_2321,N_2375);
nand U2441 (N_2441,N_2282,N_2275);
and U2442 (N_2442,N_2288,N_2290);
or U2443 (N_2443,N_2319,N_2388);
or U2444 (N_2444,N_2214,N_2372);
xnor U2445 (N_2445,N_2279,N_2371);
xnor U2446 (N_2446,N_2343,N_2230);
nand U2447 (N_2447,N_2249,N_2324);
or U2448 (N_2448,N_2330,N_2289);
nand U2449 (N_2449,N_2338,N_2252);
xnor U2450 (N_2450,N_2267,N_2380);
nand U2451 (N_2451,N_2251,N_2339);
nor U2452 (N_2452,N_2250,N_2232);
or U2453 (N_2453,N_2349,N_2382);
nand U2454 (N_2454,N_2358,N_2359);
and U2455 (N_2455,N_2318,N_2294);
nand U2456 (N_2456,N_2235,N_2208);
nand U2457 (N_2457,N_2209,N_2277);
and U2458 (N_2458,N_2316,N_2376);
and U2459 (N_2459,N_2315,N_2237);
nand U2460 (N_2460,N_2348,N_2320);
nand U2461 (N_2461,N_2312,N_2362);
nand U2462 (N_2462,N_2327,N_2307);
nand U2463 (N_2463,N_2260,N_2216);
nand U2464 (N_2464,N_2268,N_2244);
nor U2465 (N_2465,N_2332,N_2367);
xnor U2466 (N_2466,N_2245,N_2346);
nand U2467 (N_2467,N_2201,N_2228);
xor U2468 (N_2468,N_2265,N_2270);
or U2469 (N_2469,N_2283,N_2276);
nor U2470 (N_2470,N_2306,N_2366);
xor U2471 (N_2471,N_2396,N_2398);
nand U2472 (N_2472,N_2397,N_2381);
nor U2473 (N_2473,N_2254,N_2384);
or U2474 (N_2474,N_2238,N_2331);
nand U2475 (N_2475,N_2219,N_2322);
nor U2476 (N_2476,N_2241,N_2354);
nor U2477 (N_2477,N_2212,N_2202);
or U2478 (N_2478,N_2305,N_2274);
and U2479 (N_2479,N_2298,N_2292);
nand U2480 (N_2480,N_2369,N_2205);
xor U2481 (N_2481,N_2215,N_2386);
xnor U2482 (N_2482,N_2342,N_2334);
xnor U2483 (N_2483,N_2223,N_2256);
nand U2484 (N_2484,N_2239,N_2393);
nand U2485 (N_2485,N_2269,N_2247);
xor U2486 (N_2486,N_2326,N_2344);
or U2487 (N_2487,N_2314,N_2353);
and U2488 (N_2488,N_2303,N_2206);
nand U2489 (N_2489,N_2337,N_2286);
and U2490 (N_2490,N_2261,N_2266);
or U2491 (N_2491,N_2357,N_2231);
and U2492 (N_2492,N_2389,N_2385);
or U2493 (N_2493,N_2243,N_2347);
nand U2494 (N_2494,N_2308,N_2203);
nand U2495 (N_2495,N_2394,N_2242);
and U2496 (N_2496,N_2258,N_2227);
nor U2497 (N_2497,N_2365,N_2304);
xnor U2498 (N_2498,N_2253,N_2391);
xnor U2499 (N_2499,N_2379,N_2220);
nand U2500 (N_2500,N_2313,N_2318);
nor U2501 (N_2501,N_2235,N_2398);
or U2502 (N_2502,N_2389,N_2218);
and U2503 (N_2503,N_2251,N_2347);
xnor U2504 (N_2504,N_2264,N_2321);
or U2505 (N_2505,N_2373,N_2269);
xor U2506 (N_2506,N_2230,N_2349);
and U2507 (N_2507,N_2271,N_2376);
or U2508 (N_2508,N_2291,N_2399);
nor U2509 (N_2509,N_2340,N_2218);
nor U2510 (N_2510,N_2336,N_2361);
xor U2511 (N_2511,N_2242,N_2393);
or U2512 (N_2512,N_2248,N_2350);
and U2513 (N_2513,N_2263,N_2218);
xnor U2514 (N_2514,N_2397,N_2302);
nand U2515 (N_2515,N_2360,N_2243);
or U2516 (N_2516,N_2382,N_2353);
nand U2517 (N_2517,N_2298,N_2380);
or U2518 (N_2518,N_2300,N_2318);
xnor U2519 (N_2519,N_2274,N_2389);
nand U2520 (N_2520,N_2340,N_2212);
or U2521 (N_2521,N_2268,N_2246);
or U2522 (N_2522,N_2230,N_2279);
xor U2523 (N_2523,N_2301,N_2249);
and U2524 (N_2524,N_2320,N_2208);
nor U2525 (N_2525,N_2321,N_2347);
nand U2526 (N_2526,N_2311,N_2281);
nor U2527 (N_2527,N_2302,N_2323);
xor U2528 (N_2528,N_2299,N_2366);
nand U2529 (N_2529,N_2337,N_2378);
and U2530 (N_2530,N_2307,N_2305);
xor U2531 (N_2531,N_2386,N_2364);
or U2532 (N_2532,N_2314,N_2267);
nand U2533 (N_2533,N_2326,N_2231);
xor U2534 (N_2534,N_2296,N_2245);
xnor U2535 (N_2535,N_2301,N_2297);
and U2536 (N_2536,N_2252,N_2393);
nor U2537 (N_2537,N_2241,N_2396);
nand U2538 (N_2538,N_2271,N_2309);
nand U2539 (N_2539,N_2366,N_2326);
nor U2540 (N_2540,N_2248,N_2302);
xor U2541 (N_2541,N_2293,N_2248);
and U2542 (N_2542,N_2275,N_2325);
xor U2543 (N_2543,N_2223,N_2293);
xor U2544 (N_2544,N_2330,N_2219);
xor U2545 (N_2545,N_2202,N_2353);
xnor U2546 (N_2546,N_2271,N_2312);
nor U2547 (N_2547,N_2350,N_2317);
or U2548 (N_2548,N_2322,N_2229);
nor U2549 (N_2549,N_2375,N_2370);
or U2550 (N_2550,N_2230,N_2276);
nand U2551 (N_2551,N_2336,N_2210);
or U2552 (N_2552,N_2375,N_2319);
xor U2553 (N_2553,N_2269,N_2240);
xor U2554 (N_2554,N_2203,N_2358);
nand U2555 (N_2555,N_2250,N_2351);
xor U2556 (N_2556,N_2250,N_2312);
nor U2557 (N_2557,N_2393,N_2275);
nand U2558 (N_2558,N_2263,N_2220);
nor U2559 (N_2559,N_2387,N_2338);
xor U2560 (N_2560,N_2335,N_2347);
nand U2561 (N_2561,N_2380,N_2235);
nand U2562 (N_2562,N_2255,N_2338);
nand U2563 (N_2563,N_2320,N_2371);
nand U2564 (N_2564,N_2340,N_2219);
xnor U2565 (N_2565,N_2281,N_2357);
or U2566 (N_2566,N_2358,N_2363);
and U2567 (N_2567,N_2265,N_2227);
nor U2568 (N_2568,N_2203,N_2281);
nand U2569 (N_2569,N_2306,N_2215);
xnor U2570 (N_2570,N_2365,N_2228);
xnor U2571 (N_2571,N_2222,N_2261);
and U2572 (N_2572,N_2309,N_2356);
and U2573 (N_2573,N_2201,N_2334);
and U2574 (N_2574,N_2270,N_2383);
or U2575 (N_2575,N_2324,N_2262);
and U2576 (N_2576,N_2377,N_2329);
xnor U2577 (N_2577,N_2201,N_2373);
and U2578 (N_2578,N_2351,N_2239);
xnor U2579 (N_2579,N_2261,N_2327);
and U2580 (N_2580,N_2357,N_2218);
nand U2581 (N_2581,N_2350,N_2327);
xnor U2582 (N_2582,N_2264,N_2237);
nor U2583 (N_2583,N_2345,N_2208);
nand U2584 (N_2584,N_2305,N_2252);
nor U2585 (N_2585,N_2239,N_2238);
or U2586 (N_2586,N_2316,N_2358);
xnor U2587 (N_2587,N_2265,N_2381);
nand U2588 (N_2588,N_2356,N_2228);
nand U2589 (N_2589,N_2262,N_2351);
nor U2590 (N_2590,N_2395,N_2376);
or U2591 (N_2591,N_2240,N_2276);
nand U2592 (N_2592,N_2212,N_2356);
nor U2593 (N_2593,N_2202,N_2277);
xor U2594 (N_2594,N_2282,N_2281);
or U2595 (N_2595,N_2209,N_2216);
nand U2596 (N_2596,N_2200,N_2267);
and U2597 (N_2597,N_2222,N_2317);
nor U2598 (N_2598,N_2265,N_2203);
nand U2599 (N_2599,N_2335,N_2224);
and U2600 (N_2600,N_2560,N_2420);
or U2601 (N_2601,N_2503,N_2489);
or U2602 (N_2602,N_2491,N_2576);
nor U2603 (N_2603,N_2413,N_2557);
nor U2604 (N_2604,N_2407,N_2554);
or U2605 (N_2605,N_2467,N_2493);
nor U2606 (N_2606,N_2505,N_2518);
nand U2607 (N_2607,N_2444,N_2516);
xnor U2608 (N_2608,N_2547,N_2578);
xnor U2609 (N_2609,N_2598,N_2488);
xor U2610 (N_2610,N_2404,N_2574);
or U2611 (N_2611,N_2590,N_2446);
nand U2612 (N_2612,N_2411,N_2566);
and U2613 (N_2613,N_2401,N_2545);
and U2614 (N_2614,N_2421,N_2573);
or U2615 (N_2615,N_2432,N_2502);
nor U2616 (N_2616,N_2452,N_2497);
nor U2617 (N_2617,N_2408,N_2400);
nor U2618 (N_2618,N_2461,N_2539);
nand U2619 (N_2619,N_2559,N_2438);
nor U2620 (N_2620,N_2422,N_2546);
or U2621 (N_2621,N_2511,N_2485);
nand U2622 (N_2622,N_2577,N_2477);
or U2623 (N_2623,N_2439,N_2427);
xnor U2624 (N_2624,N_2522,N_2478);
nand U2625 (N_2625,N_2445,N_2558);
nand U2626 (N_2626,N_2454,N_2423);
and U2627 (N_2627,N_2563,N_2464);
nand U2628 (N_2628,N_2580,N_2415);
nor U2629 (N_2629,N_2515,N_2528);
or U2630 (N_2630,N_2517,N_2429);
nor U2631 (N_2631,N_2537,N_2500);
nand U2632 (N_2632,N_2523,N_2410);
xor U2633 (N_2633,N_2456,N_2565);
xnor U2634 (N_2634,N_2584,N_2442);
or U2635 (N_2635,N_2530,N_2586);
xnor U2636 (N_2636,N_2469,N_2552);
nand U2637 (N_2637,N_2480,N_2436);
and U2638 (N_2638,N_2506,N_2431);
nor U2639 (N_2639,N_2570,N_2510);
nand U2640 (N_2640,N_2450,N_2443);
or U2641 (N_2641,N_2426,N_2593);
xor U2642 (N_2642,N_2466,N_2541);
nand U2643 (N_2643,N_2476,N_2535);
nand U2644 (N_2644,N_2462,N_2409);
xnor U2645 (N_2645,N_2588,N_2504);
xor U2646 (N_2646,N_2428,N_2441);
and U2647 (N_2647,N_2542,N_2499);
xnor U2648 (N_2648,N_2472,N_2507);
and U2649 (N_2649,N_2587,N_2481);
xnor U2650 (N_2650,N_2520,N_2457);
xor U2651 (N_2651,N_2549,N_2406);
or U2652 (N_2652,N_2562,N_2583);
nand U2653 (N_2653,N_2434,N_2596);
or U2654 (N_2654,N_2575,N_2448);
xnor U2655 (N_2655,N_2526,N_2533);
or U2656 (N_2656,N_2459,N_2498);
and U2657 (N_2657,N_2585,N_2550);
nand U2658 (N_2658,N_2468,N_2402);
nand U2659 (N_2659,N_2571,N_2403);
nand U2660 (N_2660,N_2569,N_2555);
nor U2661 (N_2661,N_2465,N_2484);
and U2662 (N_2662,N_2486,N_2433);
xor U2663 (N_2663,N_2591,N_2492);
xor U2664 (N_2664,N_2473,N_2599);
nor U2665 (N_2665,N_2544,N_2471);
or U2666 (N_2666,N_2487,N_2412);
or U2667 (N_2667,N_2567,N_2532);
xor U2668 (N_2668,N_2548,N_2536);
xor U2669 (N_2669,N_2538,N_2531);
and U2670 (N_2670,N_2579,N_2509);
and U2671 (N_2671,N_2524,N_2551);
and U2672 (N_2672,N_2460,N_2529);
nor U2673 (N_2673,N_2474,N_2458);
nor U2674 (N_2674,N_2494,N_2597);
xnor U2675 (N_2675,N_2540,N_2495);
xor U2676 (N_2676,N_2534,N_2514);
or U2677 (N_2677,N_2483,N_2424);
nor U2678 (N_2678,N_2525,N_2453);
nor U2679 (N_2679,N_2418,N_2527);
xnor U2680 (N_2680,N_2589,N_2508);
or U2681 (N_2681,N_2572,N_2419);
and U2682 (N_2682,N_2553,N_2496);
nor U2683 (N_2683,N_2564,N_2512);
xnor U2684 (N_2684,N_2581,N_2519);
xor U2685 (N_2685,N_2592,N_2447);
and U2686 (N_2686,N_2425,N_2435);
xor U2687 (N_2687,N_2451,N_2455);
or U2688 (N_2688,N_2437,N_2595);
nand U2689 (N_2689,N_2417,N_2405);
nand U2690 (N_2690,N_2470,N_2561);
or U2691 (N_2691,N_2543,N_2521);
nand U2692 (N_2692,N_2594,N_2513);
and U2693 (N_2693,N_2463,N_2416);
nor U2694 (N_2694,N_2449,N_2430);
or U2695 (N_2695,N_2582,N_2440);
nand U2696 (N_2696,N_2501,N_2479);
nand U2697 (N_2697,N_2414,N_2556);
nand U2698 (N_2698,N_2482,N_2490);
nor U2699 (N_2699,N_2568,N_2475);
or U2700 (N_2700,N_2578,N_2462);
xnor U2701 (N_2701,N_2447,N_2556);
and U2702 (N_2702,N_2471,N_2445);
and U2703 (N_2703,N_2488,N_2450);
and U2704 (N_2704,N_2400,N_2482);
nand U2705 (N_2705,N_2411,N_2414);
nor U2706 (N_2706,N_2521,N_2441);
xnor U2707 (N_2707,N_2528,N_2561);
or U2708 (N_2708,N_2414,N_2475);
xor U2709 (N_2709,N_2501,N_2523);
and U2710 (N_2710,N_2462,N_2546);
xor U2711 (N_2711,N_2506,N_2481);
xor U2712 (N_2712,N_2477,N_2530);
nand U2713 (N_2713,N_2553,N_2508);
xnor U2714 (N_2714,N_2441,N_2565);
or U2715 (N_2715,N_2508,N_2415);
xnor U2716 (N_2716,N_2456,N_2427);
xnor U2717 (N_2717,N_2411,N_2582);
nor U2718 (N_2718,N_2565,N_2526);
or U2719 (N_2719,N_2516,N_2543);
nand U2720 (N_2720,N_2527,N_2405);
nor U2721 (N_2721,N_2579,N_2590);
and U2722 (N_2722,N_2474,N_2532);
or U2723 (N_2723,N_2454,N_2555);
or U2724 (N_2724,N_2470,N_2499);
or U2725 (N_2725,N_2569,N_2507);
nor U2726 (N_2726,N_2454,N_2584);
or U2727 (N_2727,N_2534,N_2559);
nor U2728 (N_2728,N_2524,N_2572);
or U2729 (N_2729,N_2504,N_2561);
or U2730 (N_2730,N_2429,N_2553);
nand U2731 (N_2731,N_2568,N_2488);
and U2732 (N_2732,N_2440,N_2563);
nor U2733 (N_2733,N_2405,N_2524);
nor U2734 (N_2734,N_2495,N_2511);
or U2735 (N_2735,N_2420,N_2552);
xnor U2736 (N_2736,N_2471,N_2440);
nor U2737 (N_2737,N_2572,N_2582);
and U2738 (N_2738,N_2536,N_2483);
nand U2739 (N_2739,N_2441,N_2561);
or U2740 (N_2740,N_2527,N_2431);
and U2741 (N_2741,N_2599,N_2516);
or U2742 (N_2742,N_2598,N_2529);
xor U2743 (N_2743,N_2564,N_2458);
or U2744 (N_2744,N_2578,N_2566);
and U2745 (N_2745,N_2474,N_2443);
nand U2746 (N_2746,N_2596,N_2546);
xor U2747 (N_2747,N_2432,N_2459);
nor U2748 (N_2748,N_2538,N_2588);
nand U2749 (N_2749,N_2579,N_2448);
nor U2750 (N_2750,N_2454,N_2464);
or U2751 (N_2751,N_2520,N_2538);
nor U2752 (N_2752,N_2421,N_2542);
and U2753 (N_2753,N_2470,N_2587);
nor U2754 (N_2754,N_2405,N_2476);
nor U2755 (N_2755,N_2478,N_2559);
nor U2756 (N_2756,N_2505,N_2455);
xor U2757 (N_2757,N_2572,N_2502);
or U2758 (N_2758,N_2481,N_2441);
xnor U2759 (N_2759,N_2418,N_2465);
nor U2760 (N_2760,N_2487,N_2448);
nor U2761 (N_2761,N_2437,N_2569);
nand U2762 (N_2762,N_2527,N_2594);
nand U2763 (N_2763,N_2495,N_2488);
xnor U2764 (N_2764,N_2412,N_2406);
or U2765 (N_2765,N_2537,N_2521);
nand U2766 (N_2766,N_2524,N_2434);
or U2767 (N_2767,N_2545,N_2539);
and U2768 (N_2768,N_2555,N_2455);
or U2769 (N_2769,N_2536,N_2440);
nor U2770 (N_2770,N_2599,N_2458);
nor U2771 (N_2771,N_2477,N_2459);
or U2772 (N_2772,N_2483,N_2433);
or U2773 (N_2773,N_2460,N_2579);
and U2774 (N_2774,N_2403,N_2564);
and U2775 (N_2775,N_2480,N_2460);
nor U2776 (N_2776,N_2491,N_2543);
or U2777 (N_2777,N_2549,N_2419);
or U2778 (N_2778,N_2507,N_2578);
or U2779 (N_2779,N_2449,N_2411);
and U2780 (N_2780,N_2409,N_2469);
and U2781 (N_2781,N_2413,N_2446);
nor U2782 (N_2782,N_2534,N_2464);
or U2783 (N_2783,N_2411,N_2487);
xor U2784 (N_2784,N_2426,N_2512);
or U2785 (N_2785,N_2522,N_2590);
or U2786 (N_2786,N_2477,N_2441);
nand U2787 (N_2787,N_2468,N_2462);
xor U2788 (N_2788,N_2459,N_2404);
or U2789 (N_2789,N_2420,N_2530);
nor U2790 (N_2790,N_2592,N_2402);
and U2791 (N_2791,N_2471,N_2541);
nor U2792 (N_2792,N_2467,N_2423);
nand U2793 (N_2793,N_2536,N_2546);
or U2794 (N_2794,N_2433,N_2575);
xor U2795 (N_2795,N_2479,N_2540);
xor U2796 (N_2796,N_2460,N_2555);
nand U2797 (N_2797,N_2584,N_2554);
xor U2798 (N_2798,N_2537,N_2485);
nor U2799 (N_2799,N_2426,N_2535);
nand U2800 (N_2800,N_2746,N_2695);
nor U2801 (N_2801,N_2782,N_2671);
and U2802 (N_2802,N_2771,N_2692);
and U2803 (N_2803,N_2730,N_2648);
nor U2804 (N_2804,N_2630,N_2742);
xnor U2805 (N_2805,N_2796,N_2716);
nor U2806 (N_2806,N_2772,N_2732);
nand U2807 (N_2807,N_2646,N_2724);
nand U2808 (N_2808,N_2634,N_2609);
or U2809 (N_2809,N_2779,N_2709);
nand U2810 (N_2810,N_2715,N_2728);
nor U2811 (N_2811,N_2721,N_2623);
or U2812 (N_2812,N_2621,N_2668);
nand U2813 (N_2813,N_2613,N_2679);
nand U2814 (N_2814,N_2693,N_2641);
xor U2815 (N_2815,N_2615,N_2770);
xor U2816 (N_2816,N_2755,N_2708);
or U2817 (N_2817,N_2763,N_2751);
nor U2818 (N_2818,N_2774,N_2685);
or U2819 (N_2819,N_2794,N_2756);
and U2820 (N_2820,N_2778,N_2667);
or U2821 (N_2821,N_2665,N_2786);
nor U2822 (N_2822,N_2725,N_2745);
and U2823 (N_2823,N_2768,N_2645);
or U2824 (N_2824,N_2792,N_2678);
xor U2825 (N_2825,N_2717,N_2736);
nand U2826 (N_2826,N_2636,N_2686);
and U2827 (N_2827,N_2750,N_2602);
or U2828 (N_2828,N_2601,N_2637);
and U2829 (N_2829,N_2731,N_2694);
or U2830 (N_2830,N_2647,N_2787);
or U2831 (N_2831,N_2690,N_2656);
or U2832 (N_2832,N_2780,N_2722);
xnor U2833 (N_2833,N_2767,N_2727);
or U2834 (N_2834,N_2799,N_2652);
nor U2835 (N_2835,N_2669,N_2775);
and U2836 (N_2836,N_2655,N_2748);
nor U2837 (N_2837,N_2659,N_2657);
or U2838 (N_2838,N_2705,N_2714);
or U2839 (N_2839,N_2629,N_2624);
and U2840 (N_2840,N_2710,N_2622);
nand U2841 (N_2841,N_2631,N_2611);
nand U2842 (N_2842,N_2712,N_2612);
or U2843 (N_2843,N_2762,N_2761);
or U2844 (N_2844,N_2789,N_2711);
or U2845 (N_2845,N_2610,N_2688);
xnor U2846 (N_2846,N_2749,N_2600);
nand U2847 (N_2847,N_2639,N_2733);
nor U2848 (N_2848,N_2752,N_2700);
and U2849 (N_2849,N_2698,N_2619);
nor U2850 (N_2850,N_2654,N_2642);
nand U2851 (N_2851,N_2798,N_2633);
nor U2852 (N_2852,N_2726,N_2741);
or U2853 (N_2853,N_2754,N_2765);
xnor U2854 (N_2854,N_2651,N_2662);
and U2855 (N_2855,N_2674,N_2660);
xnor U2856 (N_2856,N_2672,N_2643);
and U2857 (N_2857,N_2777,N_2735);
and U2858 (N_2858,N_2653,N_2719);
or U2859 (N_2859,N_2783,N_2743);
and U2860 (N_2860,N_2720,N_2682);
xnor U2861 (N_2861,N_2784,N_2677);
xor U2862 (N_2862,N_2625,N_2627);
nand U2863 (N_2863,N_2684,N_2753);
nor U2864 (N_2864,N_2683,N_2607);
xnor U2865 (N_2865,N_2758,N_2680);
xnor U2866 (N_2866,N_2616,N_2704);
nand U2867 (N_2867,N_2666,N_2790);
xor U2868 (N_2868,N_2744,N_2797);
xor U2869 (N_2869,N_2661,N_2632);
or U2870 (N_2870,N_2729,N_2608);
or U2871 (N_2871,N_2658,N_2793);
or U2872 (N_2872,N_2785,N_2764);
or U2873 (N_2873,N_2603,N_2617);
xor U2874 (N_2874,N_2697,N_2740);
or U2875 (N_2875,N_2759,N_2675);
nor U2876 (N_2876,N_2673,N_2644);
nor U2877 (N_2877,N_2618,N_2663);
nand U2878 (N_2878,N_2649,N_2626);
xor U2879 (N_2879,N_2606,N_2769);
or U2880 (N_2880,N_2773,N_2687);
or U2881 (N_2881,N_2718,N_2691);
or U2882 (N_2882,N_2676,N_2635);
and U2883 (N_2883,N_2734,N_2737);
nor U2884 (N_2884,N_2670,N_2620);
or U2885 (N_2885,N_2604,N_2791);
xnor U2886 (N_2886,N_2706,N_2605);
xnor U2887 (N_2887,N_2713,N_2707);
and U2888 (N_2888,N_2788,N_2723);
nor U2889 (N_2889,N_2640,N_2766);
or U2890 (N_2890,N_2638,N_2703);
and U2891 (N_2891,N_2650,N_2702);
or U2892 (N_2892,N_2760,N_2701);
or U2893 (N_2893,N_2699,N_2696);
and U2894 (N_2894,N_2628,N_2776);
nor U2895 (N_2895,N_2689,N_2781);
nor U2896 (N_2896,N_2757,N_2739);
xnor U2897 (N_2897,N_2795,N_2614);
nand U2898 (N_2898,N_2747,N_2681);
or U2899 (N_2899,N_2664,N_2738);
or U2900 (N_2900,N_2608,N_2713);
xnor U2901 (N_2901,N_2684,N_2754);
nor U2902 (N_2902,N_2710,N_2749);
nand U2903 (N_2903,N_2785,N_2628);
and U2904 (N_2904,N_2623,N_2768);
or U2905 (N_2905,N_2798,N_2651);
nor U2906 (N_2906,N_2700,N_2796);
xor U2907 (N_2907,N_2769,N_2637);
nor U2908 (N_2908,N_2715,N_2662);
or U2909 (N_2909,N_2727,N_2698);
nand U2910 (N_2910,N_2734,N_2774);
nand U2911 (N_2911,N_2764,N_2690);
nor U2912 (N_2912,N_2794,N_2752);
nor U2913 (N_2913,N_2611,N_2650);
nor U2914 (N_2914,N_2744,N_2756);
and U2915 (N_2915,N_2628,N_2696);
nand U2916 (N_2916,N_2612,N_2711);
nor U2917 (N_2917,N_2779,N_2677);
or U2918 (N_2918,N_2631,N_2626);
and U2919 (N_2919,N_2658,N_2784);
or U2920 (N_2920,N_2728,N_2635);
and U2921 (N_2921,N_2733,N_2718);
and U2922 (N_2922,N_2636,N_2667);
nand U2923 (N_2923,N_2678,N_2766);
nand U2924 (N_2924,N_2757,N_2603);
nand U2925 (N_2925,N_2641,N_2723);
or U2926 (N_2926,N_2782,N_2606);
nand U2927 (N_2927,N_2741,N_2688);
nor U2928 (N_2928,N_2791,N_2601);
nor U2929 (N_2929,N_2747,N_2787);
xnor U2930 (N_2930,N_2655,N_2606);
xnor U2931 (N_2931,N_2630,N_2635);
or U2932 (N_2932,N_2724,N_2786);
and U2933 (N_2933,N_2660,N_2617);
and U2934 (N_2934,N_2614,N_2633);
nand U2935 (N_2935,N_2758,N_2694);
or U2936 (N_2936,N_2763,N_2654);
nor U2937 (N_2937,N_2693,N_2616);
nand U2938 (N_2938,N_2629,N_2614);
nor U2939 (N_2939,N_2693,N_2666);
and U2940 (N_2940,N_2751,N_2748);
or U2941 (N_2941,N_2721,N_2766);
and U2942 (N_2942,N_2634,N_2670);
nand U2943 (N_2943,N_2646,N_2757);
nor U2944 (N_2944,N_2723,N_2681);
and U2945 (N_2945,N_2610,N_2736);
nor U2946 (N_2946,N_2750,N_2686);
nand U2947 (N_2947,N_2706,N_2610);
and U2948 (N_2948,N_2683,N_2692);
nor U2949 (N_2949,N_2662,N_2778);
nor U2950 (N_2950,N_2686,N_2711);
nand U2951 (N_2951,N_2789,N_2738);
xor U2952 (N_2952,N_2666,N_2773);
or U2953 (N_2953,N_2678,N_2697);
or U2954 (N_2954,N_2624,N_2791);
and U2955 (N_2955,N_2671,N_2742);
or U2956 (N_2956,N_2718,N_2658);
nor U2957 (N_2957,N_2750,N_2743);
nor U2958 (N_2958,N_2626,N_2711);
and U2959 (N_2959,N_2608,N_2789);
nor U2960 (N_2960,N_2725,N_2681);
and U2961 (N_2961,N_2614,N_2654);
and U2962 (N_2962,N_2600,N_2623);
nand U2963 (N_2963,N_2786,N_2687);
nand U2964 (N_2964,N_2632,N_2642);
nand U2965 (N_2965,N_2660,N_2600);
nor U2966 (N_2966,N_2768,N_2701);
or U2967 (N_2967,N_2678,N_2603);
nand U2968 (N_2968,N_2693,N_2639);
nor U2969 (N_2969,N_2749,N_2664);
and U2970 (N_2970,N_2671,N_2711);
xnor U2971 (N_2971,N_2636,N_2755);
nor U2972 (N_2972,N_2724,N_2687);
and U2973 (N_2973,N_2787,N_2604);
and U2974 (N_2974,N_2662,N_2614);
or U2975 (N_2975,N_2636,N_2662);
nand U2976 (N_2976,N_2676,N_2652);
nand U2977 (N_2977,N_2623,N_2788);
and U2978 (N_2978,N_2789,N_2754);
nor U2979 (N_2979,N_2765,N_2793);
or U2980 (N_2980,N_2609,N_2765);
nand U2981 (N_2981,N_2768,N_2784);
and U2982 (N_2982,N_2692,N_2682);
xnor U2983 (N_2983,N_2745,N_2677);
xnor U2984 (N_2984,N_2793,N_2603);
and U2985 (N_2985,N_2751,N_2798);
nand U2986 (N_2986,N_2604,N_2642);
xor U2987 (N_2987,N_2780,N_2651);
xnor U2988 (N_2988,N_2718,N_2665);
and U2989 (N_2989,N_2658,N_2743);
nor U2990 (N_2990,N_2628,N_2608);
xor U2991 (N_2991,N_2777,N_2786);
nor U2992 (N_2992,N_2690,N_2785);
xor U2993 (N_2993,N_2729,N_2710);
nand U2994 (N_2994,N_2694,N_2705);
and U2995 (N_2995,N_2701,N_2611);
nor U2996 (N_2996,N_2684,N_2662);
or U2997 (N_2997,N_2737,N_2763);
nor U2998 (N_2998,N_2769,N_2742);
nand U2999 (N_2999,N_2680,N_2666);
nand UO_0 (O_0,N_2952,N_2869);
and UO_1 (O_1,N_2822,N_2821);
and UO_2 (O_2,N_2941,N_2917);
and UO_3 (O_3,N_2824,N_2925);
nor UO_4 (O_4,N_2988,N_2995);
or UO_5 (O_5,N_2963,N_2845);
or UO_6 (O_6,N_2889,N_2851);
and UO_7 (O_7,N_2826,N_2872);
and UO_8 (O_8,N_2998,N_2823);
and UO_9 (O_9,N_2965,N_2959);
nand UO_10 (O_10,N_2895,N_2996);
or UO_11 (O_11,N_2841,N_2816);
and UO_12 (O_12,N_2871,N_2942);
xor UO_13 (O_13,N_2979,N_2908);
or UO_14 (O_14,N_2849,N_2968);
nand UO_15 (O_15,N_2837,N_2804);
nor UO_16 (O_16,N_2880,N_2852);
and UO_17 (O_17,N_2817,N_2948);
xor UO_18 (O_18,N_2801,N_2812);
nand UO_19 (O_19,N_2805,N_2915);
nand UO_20 (O_20,N_2928,N_2904);
or UO_21 (O_21,N_2985,N_2836);
nand UO_22 (O_22,N_2840,N_2947);
nand UO_23 (O_23,N_2974,N_2819);
nand UO_24 (O_24,N_2896,N_2926);
nor UO_25 (O_25,N_2954,N_2961);
and UO_26 (O_26,N_2914,N_2986);
or UO_27 (O_27,N_2936,N_2885);
nor UO_28 (O_28,N_2982,N_2859);
and UO_29 (O_29,N_2879,N_2883);
xor UO_30 (O_30,N_2861,N_2981);
and UO_31 (O_31,N_2960,N_2882);
xnor UO_32 (O_32,N_2847,N_2910);
nand UO_33 (O_33,N_2802,N_2903);
or UO_34 (O_34,N_2943,N_2976);
or UO_35 (O_35,N_2810,N_2829);
nor UO_36 (O_36,N_2980,N_2811);
nor UO_37 (O_37,N_2983,N_2935);
and UO_38 (O_38,N_2843,N_2956);
and UO_39 (O_39,N_2932,N_2833);
and UO_40 (O_40,N_2828,N_2875);
and UO_41 (O_41,N_2938,N_2940);
and UO_42 (O_42,N_2993,N_2884);
xnor UO_43 (O_43,N_2853,N_2806);
nand UO_44 (O_44,N_2870,N_2962);
nor UO_45 (O_45,N_2873,N_2838);
xor UO_46 (O_46,N_2808,N_2860);
or UO_47 (O_47,N_2957,N_2975);
and UO_48 (O_48,N_2877,N_2930);
and UO_49 (O_49,N_2858,N_2892);
xor UO_50 (O_50,N_2803,N_2978);
nor UO_51 (O_51,N_2813,N_2815);
or UO_52 (O_52,N_2835,N_2920);
nor UO_53 (O_53,N_2929,N_2951);
xnor UO_54 (O_54,N_2878,N_2814);
or UO_55 (O_55,N_2827,N_2839);
and UO_56 (O_56,N_2939,N_2832);
nor UO_57 (O_57,N_2970,N_2863);
nor UO_58 (O_58,N_2987,N_2866);
nor UO_59 (O_59,N_2900,N_2830);
and UO_60 (O_60,N_2897,N_2992);
xnor UO_61 (O_61,N_2967,N_2955);
nor UO_62 (O_62,N_2906,N_2977);
nor UO_63 (O_63,N_2807,N_2902);
nor UO_64 (O_64,N_2831,N_2958);
and UO_65 (O_65,N_2834,N_2887);
and UO_66 (O_66,N_2850,N_2891);
or UO_67 (O_67,N_2905,N_2874);
nand UO_68 (O_68,N_2944,N_2886);
nand UO_69 (O_69,N_2950,N_2933);
xnor UO_70 (O_70,N_2818,N_2997);
nand UO_71 (O_71,N_2964,N_2868);
xnor UO_72 (O_72,N_2898,N_2862);
nor UO_73 (O_73,N_2894,N_2972);
or UO_74 (O_74,N_2876,N_2909);
nor UO_75 (O_75,N_2984,N_2971);
xnor UO_76 (O_76,N_2888,N_2922);
or UO_77 (O_77,N_2969,N_2800);
and UO_78 (O_78,N_2867,N_2890);
nand UO_79 (O_79,N_2991,N_2927);
or UO_80 (O_80,N_2809,N_2848);
or UO_81 (O_81,N_2913,N_2973);
or UO_82 (O_82,N_2923,N_2899);
nand UO_83 (O_83,N_2953,N_2855);
nor UO_84 (O_84,N_2966,N_2989);
and UO_85 (O_85,N_2911,N_2916);
nor UO_86 (O_86,N_2994,N_2999);
or UO_87 (O_87,N_2912,N_2934);
and UO_88 (O_88,N_2901,N_2842);
nor UO_89 (O_89,N_2921,N_2893);
nor UO_90 (O_90,N_2946,N_2924);
and UO_91 (O_91,N_2820,N_2881);
nor UO_92 (O_92,N_2931,N_2937);
nand UO_93 (O_93,N_2918,N_2864);
and UO_94 (O_94,N_2854,N_2857);
and UO_95 (O_95,N_2945,N_2949);
nand UO_96 (O_96,N_2865,N_2907);
nor UO_97 (O_97,N_2846,N_2844);
and UO_98 (O_98,N_2856,N_2919);
nand UO_99 (O_99,N_2825,N_2990);
xor UO_100 (O_100,N_2932,N_2940);
and UO_101 (O_101,N_2848,N_2804);
nor UO_102 (O_102,N_2989,N_2994);
xor UO_103 (O_103,N_2870,N_2868);
nor UO_104 (O_104,N_2959,N_2920);
and UO_105 (O_105,N_2817,N_2992);
nor UO_106 (O_106,N_2907,N_2843);
xnor UO_107 (O_107,N_2890,N_2934);
or UO_108 (O_108,N_2800,N_2866);
nand UO_109 (O_109,N_2940,N_2931);
and UO_110 (O_110,N_2822,N_2865);
or UO_111 (O_111,N_2801,N_2879);
nand UO_112 (O_112,N_2849,N_2863);
and UO_113 (O_113,N_2951,N_2804);
and UO_114 (O_114,N_2871,N_2892);
nor UO_115 (O_115,N_2867,N_2922);
nor UO_116 (O_116,N_2832,N_2993);
and UO_117 (O_117,N_2829,N_2921);
and UO_118 (O_118,N_2827,N_2804);
nand UO_119 (O_119,N_2980,N_2948);
xnor UO_120 (O_120,N_2961,N_2886);
or UO_121 (O_121,N_2964,N_2811);
or UO_122 (O_122,N_2806,N_2803);
and UO_123 (O_123,N_2988,N_2922);
xor UO_124 (O_124,N_2818,N_2866);
nand UO_125 (O_125,N_2951,N_2802);
or UO_126 (O_126,N_2925,N_2847);
and UO_127 (O_127,N_2994,N_2812);
nand UO_128 (O_128,N_2849,N_2813);
xnor UO_129 (O_129,N_2988,N_2816);
nand UO_130 (O_130,N_2842,N_2925);
or UO_131 (O_131,N_2972,N_2819);
nand UO_132 (O_132,N_2913,N_2901);
nand UO_133 (O_133,N_2971,N_2975);
and UO_134 (O_134,N_2948,N_2859);
and UO_135 (O_135,N_2979,N_2806);
nand UO_136 (O_136,N_2947,N_2826);
or UO_137 (O_137,N_2973,N_2810);
or UO_138 (O_138,N_2942,N_2935);
or UO_139 (O_139,N_2989,N_2992);
nand UO_140 (O_140,N_2813,N_2963);
xor UO_141 (O_141,N_2921,N_2823);
nand UO_142 (O_142,N_2807,N_2812);
and UO_143 (O_143,N_2944,N_2907);
xor UO_144 (O_144,N_2915,N_2845);
and UO_145 (O_145,N_2933,N_2972);
or UO_146 (O_146,N_2964,N_2923);
nor UO_147 (O_147,N_2897,N_2953);
xnor UO_148 (O_148,N_2982,N_2996);
nand UO_149 (O_149,N_2815,N_2909);
and UO_150 (O_150,N_2998,N_2979);
nor UO_151 (O_151,N_2925,N_2912);
and UO_152 (O_152,N_2805,N_2925);
or UO_153 (O_153,N_2984,N_2895);
and UO_154 (O_154,N_2836,N_2897);
nand UO_155 (O_155,N_2998,N_2988);
or UO_156 (O_156,N_2839,N_2846);
xnor UO_157 (O_157,N_2987,N_2920);
and UO_158 (O_158,N_2958,N_2851);
nand UO_159 (O_159,N_2940,N_2959);
nor UO_160 (O_160,N_2914,N_2919);
and UO_161 (O_161,N_2800,N_2835);
and UO_162 (O_162,N_2846,N_2976);
xnor UO_163 (O_163,N_2962,N_2969);
or UO_164 (O_164,N_2963,N_2835);
nand UO_165 (O_165,N_2998,N_2914);
and UO_166 (O_166,N_2831,N_2994);
xnor UO_167 (O_167,N_2806,N_2908);
nand UO_168 (O_168,N_2998,N_2919);
nand UO_169 (O_169,N_2801,N_2996);
nor UO_170 (O_170,N_2816,N_2918);
and UO_171 (O_171,N_2822,N_2874);
or UO_172 (O_172,N_2884,N_2976);
nor UO_173 (O_173,N_2911,N_2950);
or UO_174 (O_174,N_2849,N_2930);
nor UO_175 (O_175,N_2855,N_2829);
xor UO_176 (O_176,N_2809,N_2814);
nor UO_177 (O_177,N_2939,N_2871);
and UO_178 (O_178,N_2980,N_2834);
nand UO_179 (O_179,N_2922,N_2941);
and UO_180 (O_180,N_2835,N_2857);
nand UO_181 (O_181,N_2802,N_2878);
nand UO_182 (O_182,N_2972,N_2801);
nor UO_183 (O_183,N_2963,N_2853);
nor UO_184 (O_184,N_2988,N_2978);
nor UO_185 (O_185,N_2876,N_2967);
xor UO_186 (O_186,N_2948,N_2993);
xor UO_187 (O_187,N_2893,N_2843);
nand UO_188 (O_188,N_2905,N_2894);
xnor UO_189 (O_189,N_2800,N_2862);
nand UO_190 (O_190,N_2992,N_2844);
nor UO_191 (O_191,N_2861,N_2927);
nand UO_192 (O_192,N_2891,N_2999);
nor UO_193 (O_193,N_2845,N_2953);
xor UO_194 (O_194,N_2917,N_2956);
nand UO_195 (O_195,N_2989,N_2932);
nor UO_196 (O_196,N_2868,N_2861);
and UO_197 (O_197,N_2992,N_2907);
nand UO_198 (O_198,N_2864,N_2972);
or UO_199 (O_199,N_2814,N_2945);
or UO_200 (O_200,N_2972,N_2960);
nand UO_201 (O_201,N_2846,N_2966);
or UO_202 (O_202,N_2863,N_2831);
or UO_203 (O_203,N_2826,N_2959);
xor UO_204 (O_204,N_2904,N_2948);
xnor UO_205 (O_205,N_2912,N_2980);
nand UO_206 (O_206,N_2925,N_2969);
nand UO_207 (O_207,N_2874,N_2910);
and UO_208 (O_208,N_2993,N_2867);
nand UO_209 (O_209,N_2974,N_2806);
xnor UO_210 (O_210,N_2907,N_2949);
nand UO_211 (O_211,N_2847,N_2998);
and UO_212 (O_212,N_2809,N_2872);
nand UO_213 (O_213,N_2863,N_2972);
xor UO_214 (O_214,N_2828,N_2889);
and UO_215 (O_215,N_2865,N_2913);
or UO_216 (O_216,N_2860,N_2929);
nor UO_217 (O_217,N_2967,N_2809);
nand UO_218 (O_218,N_2802,N_2996);
nor UO_219 (O_219,N_2811,N_2805);
xor UO_220 (O_220,N_2918,N_2970);
nand UO_221 (O_221,N_2938,N_2979);
nand UO_222 (O_222,N_2800,N_2854);
nor UO_223 (O_223,N_2875,N_2919);
and UO_224 (O_224,N_2959,N_2955);
nor UO_225 (O_225,N_2801,N_2952);
nor UO_226 (O_226,N_2820,N_2857);
or UO_227 (O_227,N_2822,N_2885);
xor UO_228 (O_228,N_2918,N_2977);
nand UO_229 (O_229,N_2985,N_2961);
nor UO_230 (O_230,N_2848,N_2830);
nor UO_231 (O_231,N_2950,N_2803);
or UO_232 (O_232,N_2922,N_2878);
nand UO_233 (O_233,N_2861,N_2891);
nor UO_234 (O_234,N_2834,N_2974);
nor UO_235 (O_235,N_2875,N_2918);
or UO_236 (O_236,N_2906,N_2997);
or UO_237 (O_237,N_2995,N_2975);
and UO_238 (O_238,N_2955,N_2803);
nand UO_239 (O_239,N_2870,N_2957);
or UO_240 (O_240,N_2951,N_2874);
and UO_241 (O_241,N_2837,N_2913);
nor UO_242 (O_242,N_2941,N_2834);
and UO_243 (O_243,N_2980,N_2850);
nand UO_244 (O_244,N_2858,N_2946);
and UO_245 (O_245,N_2987,N_2843);
xnor UO_246 (O_246,N_2952,N_2826);
xor UO_247 (O_247,N_2963,N_2842);
xor UO_248 (O_248,N_2894,N_2901);
or UO_249 (O_249,N_2814,N_2991);
or UO_250 (O_250,N_2848,N_2930);
nand UO_251 (O_251,N_2979,N_2869);
nor UO_252 (O_252,N_2892,N_2925);
nand UO_253 (O_253,N_2931,N_2921);
nor UO_254 (O_254,N_2936,N_2914);
xor UO_255 (O_255,N_2927,N_2948);
xor UO_256 (O_256,N_2837,N_2819);
nand UO_257 (O_257,N_2966,N_2801);
and UO_258 (O_258,N_2951,N_2938);
nor UO_259 (O_259,N_2811,N_2927);
and UO_260 (O_260,N_2997,N_2846);
and UO_261 (O_261,N_2916,N_2938);
or UO_262 (O_262,N_2992,N_2973);
or UO_263 (O_263,N_2952,N_2948);
nand UO_264 (O_264,N_2913,N_2897);
or UO_265 (O_265,N_2968,N_2921);
xnor UO_266 (O_266,N_2878,N_2875);
or UO_267 (O_267,N_2804,N_2845);
or UO_268 (O_268,N_2936,N_2979);
nand UO_269 (O_269,N_2976,N_2892);
and UO_270 (O_270,N_2976,N_2912);
or UO_271 (O_271,N_2892,N_2855);
nand UO_272 (O_272,N_2883,N_2989);
or UO_273 (O_273,N_2930,N_2955);
nand UO_274 (O_274,N_2935,N_2846);
nor UO_275 (O_275,N_2986,N_2828);
xnor UO_276 (O_276,N_2868,N_2967);
nor UO_277 (O_277,N_2949,N_2852);
nand UO_278 (O_278,N_2969,N_2900);
nand UO_279 (O_279,N_2823,N_2853);
and UO_280 (O_280,N_2844,N_2824);
nand UO_281 (O_281,N_2814,N_2946);
xnor UO_282 (O_282,N_2885,N_2824);
and UO_283 (O_283,N_2951,N_2871);
nand UO_284 (O_284,N_2820,N_2824);
xnor UO_285 (O_285,N_2926,N_2893);
xnor UO_286 (O_286,N_2970,N_2931);
xnor UO_287 (O_287,N_2935,N_2840);
nand UO_288 (O_288,N_2974,N_2966);
and UO_289 (O_289,N_2868,N_2895);
nor UO_290 (O_290,N_2977,N_2931);
or UO_291 (O_291,N_2803,N_2985);
and UO_292 (O_292,N_2867,N_2932);
xnor UO_293 (O_293,N_2808,N_2986);
or UO_294 (O_294,N_2881,N_2855);
nand UO_295 (O_295,N_2808,N_2991);
nand UO_296 (O_296,N_2994,N_2998);
xnor UO_297 (O_297,N_2993,N_2998);
xor UO_298 (O_298,N_2884,N_2920);
nand UO_299 (O_299,N_2842,N_2992);
xnor UO_300 (O_300,N_2968,N_2816);
nor UO_301 (O_301,N_2945,N_2873);
and UO_302 (O_302,N_2824,N_2936);
nor UO_303 (O_303,N_2988,N_2823);
xor UO_304 (O_304,N_2866,N_2840);
xnor UO_305 (O_305,N_2826,N_2999);
nor UO_306 (O_306,N_2844,N_2826);
xor UO_307 (O_307,N_2817,N_2823);
and UO_308 (O_308,N_2980,N_2824);
xnor UO_309 (O_309,N_2806,N_2877);
nand UO_310 (O_310,N_2938,N_2902);
or UO_311 (O_311,N_2924,N_2872);
xor UO_312 (O_312,N_2847,N_2826);
nor UO_313 (O_313,N_2855,N_2818);
nor UO_314 (O_314,N_2970,N_2841);
and UO_315 (O_315,N_2900,N_2909);
nor UO_316 (O_316,N_2932,N_2915);
or UO_317 (O_317,N_2878,N_2931);
xnor UO_318 (O_318,N_2941,N_2811);
or UO_319 (O_319,N_2833,N_2889);
or UO_320 (O_320,N_2969,N_2887);
nand UO_321 (O_321,N_2890,N_2956);
and UO_322 (O_322,N_2979,N_2993);
nand UO_323 (O_323,N_2886,N_2909);
nand UO_324 (O_324,N_2934,N_2867);
nand UO_325 (O_325,N_2920,N_2882);
or UO_326 (O_326,N_2945,N_2829);
nor UO_327 (O_327,N_2976,N_2864);
and UO_328 (O_328,N_2926,N_2920);
nand UO_329 (O_329,N_2994,N_2859);
and UO_330 (O_330,N_2827,N_2835);
nand UO_331 (O_331,N_2839,N_2961);
nor UO_332 (O_332,N_2806,N_2983);
and UO_333 (O_333,N_2941,N_2887);
xnor UO_334 (O_334,N_2845,N_2882);
nand UO_335 (O_335,N_2963,N_2887);
nand UO_336 (O_336,N_2956,N_2972);
nor UO_337 (O_337,N_2933,N_2923);
or UO_338 (O_338,N_2894,N_2828);
and UO_339 (O_339,N_2942,N_2829);
and UO_340 (O_340,N_2929,N_2930);
or UO_341 (O_341,N_2904,N_2911);
nor UO_342 (O_342,N_2854,N_2875);
and UO_343 (O_343,N_2928,N_2890);
nor UO_344 (O_344,N_2962,N_2804);
and UO_345 (O_345,N_2979,N_2933);
xnor UO_346 (O_346,N_2849,N_2909);
nand UO_347 (O_347,N_2849,N_2864);
xnor UO_348 (O_348,N_2954,N_2876);
xnor UO_349 (O_349,N_2938,N_2983);
or UO_350 (O_350,N_2932,N_2875);
and UO_351 (O_351,N_2878,N_2991);
nand UO_352 (O_352,N_2824,N_2890);
xor UO_353 (O_353,N_2936,N_2886);
or UO_354 (O_354,N_2813,N_2960);
and UO_355 (O_355,N_2830,N_2837);
xnor UO_356 (O_356,N_2964,N_2873);
nand UO_357 (O_357,N_2824,N_2831);
xor UO_358 (O_358,N_2937,N_2929);
nor UO_359 (O_359,N_2913,N_2860);
and UO_360 (O_360,N_2866,N_2958);
or UO_361 (O_361,N_2950,N_2997);
and UO_362 (O_362,N_2942,N_2895);
xnor UO_363 (O_363,N_2900,N_2847);
or UO_364 (O_364,N_2806,N_2823);
nand UO_365 (O_365,N_2997,N_2873);
nor UO_366 (O_366,N_2933,N_2998);
xor UO_367 (O_367,N_2926,N_2871);
or UO_368 (O_368,N_2909,N_2820);
or UO_369 (O_369,N_2846,N_2953);
nor UO_370 (O_370,N_2883,N_2956);
nor UO_371 (O_371,N_2978,N_2977);
nand UO_372 (O_372,N_2977,N_2961);
and UO_373 (O_373,N_2912,N_2809);
or UO_374 (O_374,N_2961,N_2810);
xor UO_375 (O_375,N_2927,N_2804);
or UO_376 (O_376,N_2979,N_2894);
nand UO_377 (O_377,N_2964,N_2865);
xor UO_378 (O_378,N_2912,N_2817);
nor UO_379 (O_379,N_2897,N_2810);
nand UO_380 (O_380,N_2925,N_2806);
xnor UO_381 (O_381,N_2980,N_2894);
xor UO_382 (O_382,N_2983,N_2844);
xor UO_383 (O_383,N_2887,N_2829);
nor UO_384 (O_384,N_2954,N_2807);
and UO_385 (O_385,N_2911,N_2867);
nand UO_386 (O_386,N_2843,N_2982);
or UO_387 (O_387,N_2925,N_2926);
nor UO_388 (O_388,N_2923,N_2850);
or UO_389 (O_389,N_2955,N_2931);
or UO_390 (O_390,N_2912,N_2873);
xor UO_391 (O_391,N_2889,N_2944);
nor UO_392 (O_392,N_2826,N_2879);
or UO_393 (O_393,N_2845,N_2935);
nand UO_394 (O_394,N_2911,N_2913);
or UO_395 (O_395,N_2928,N_2906);
and UO_396 (O_396,N_2938,N_2851);
or UO_397 (O_397,N_2964,N_2921);
or UO_398 (O_398,N_2872,N_2959);
nor UO_399 (O_399,N_2860,N_2951);
nor UO_400 (O_400,N_2953,N_2892);
or UO_401 (O_401,N_2813,N_2900);
nand UO_402 (O_402,N_2809,N_2803);
or UO_403 (O_403,N_2873,N_2905);
xnor UO_404 (O_404,N_2969,N_2913);
or UO_405 (O_405,N_2895,N_2809);
and UO_406 (O_406,N_2864,N_2946);
or UO_407 (O_407,N_2881,N_2987);
nor UO_408 (O_408,N_2995,N_2938);
nand UO_409 (O_409,N_2854,N_2991);
xnor UO_410 (O_410,N_2850,N_2953);
xnor UO_411 (O_411,N_2827,N_2864);
or UO_412 (O_412,N_2929,N_2975);
nand UO_413 (O_413,N_2802,N_2946);
and UO_414 (O_414,N_2912,N_2871);
xor UO_415 (O_415,N_2886,N_2866);
and UO_416 (O_416,N_2880,N_2820);
or UO_417 (O_417,N_2907,N_2885);
or UO_418 (O_418,N_2968,N_2820);
or UO_419 (O_419,N_2934,N_2961);
nand UO_420 (O_420,N_2967,N_2855);
and UO_421 (O_421,N_2981,N_2920);
nor UO_422 (O_422,N_2958,N_2870);
xor UO_423 (O_423,N_2872,N_2985);
or UO_424 (O_424,N_2909,N_2920);
nand UO_425 (O_425,N_2944,N_2989);
and UO_426 (O_426,N_2975,N_2819);
or UO_427 (O_427,N_2987,N_2930);
or UO_428 (O_428,N_2987,N_2968);
or UO_429 (O_429,N_2833,N_2914);
nand UO_430 (O_430,N_2882,N_2925);
xnor UO_431 (O_431,N_2919,N_2833);
or UO_432 (O_432,N_2863,N_2899);
nand UO_433 (O_433,N_2815,N_2888);
nand UO_434 (O_434,N_2804,N_2902);
or UO_435 (O_435,N_2958,N_2934);
xnor UO_436 (O_436,N_2942,N_2989);
or UO_437 (O_437,N_2994,N_2980);
and UO_438 (O_438,N_2805,N_2946);
nand UO_439 (O_439,N_2855,N_2911);
or UO_440 (O_440,N_2904,N_2810);
nand UO_441 (O_441,N_2972,N_2853);
nand UO_442 (O_442,N_2982,N_2887);
or UO_443 (O_443,N_2949,N_2804);
or UO_444 (O_444,N_2976,N_2839);
or UO_445 (O_445,N_2894,N_2830);
and UO_446 (O_446,N_2867,N_2808);
nor UO_447 (O_447,N_2813,N_2950);
nor UO_448 (O_448,N_2872,N_2828);
and UO_449 (O_449,N_2945,N_2988);
xnor UO_450 (O_450,N_2979,N_2901);
or UO_451 (O_451,N_2913,N_2932);
nand UO_452 (O_452,N_2960,N_2990);
nand UO_453 (O_453,N_2941,N_2810);
xnor UO_454 (O_454,N_2803,N_2946);
nand UO_455 (O_455,N_2886,N_2985);
or UO_456 (O_456,N_2931,N_2853);
nor UO_457 (O_457,N_2965,N_2991);
xor UO_458 (O_458,N_2945,N_2866);
xor UO_459 (O_459,N_2964,N_2840);
and UO_460 (O_460,N_2825,N_2961);
xnor UO_461 (O_461,N_2906,N_2870);
xor UO_462 (O_462,N_2941,N_2816);
nor UO_463 (O_463,N_2896,N_2802);
or UO_464 (O_464,N_2863,N_2874);
and UO_465 (O_465,N_2810,N_2919);
and UO_466 (O_466,N_2858,N_2937);
and UO_467 (O_467,N_2871,N_2961);
nand UO_468 (O_468,N_2899,N_2853);
and UO_469 (O_469,N_2867,N_2972);
or UO_470 (O_470,N_2967,N_2988);
or UO_471 (O_471,N_2984,N_2867);
nor UO_472 (O_472,N_2864,N_2928);
and UO_473 (O_473,N_2823,N_2931);
nand UO_474 (O_474,N_2803,N_2899);
nor UO_475 (O_475,N_2979,N_2839);
and UO_476 (O_476,N_2821,N_2976);
nor UO_477 (O_477,N_2859,N_2836);
or UO_478 (O_478,N_2970,N_2844);
and UO_479 (O_479,N_2846,N_2824);
nor UO_480 (O_480,N_2801,N_2898);
and UO_481 (O_481,N_2953,N_2951);
nor UO_482 (O_482,N_2991,N_2915);
nand UO_483 (O_483,N_2849,N_2832);
and UO_484 (O_484,N_2868,N_2968);
nand UO_485 (O_485,N_2981,N_2954);
nand UO_486 (O_486,N_2865,N_2984);
and UO_487 (O_487,N_2959,N_2923);
nor UO_488 (O_488,N_2886,N_2981);
nand UO_489 (O_489,N_2826,N_2988);
nand UO_490 (O_490,N_2879,N_2928);
or UO_491 (O_491,N_2913,N_2958);
xnor UO_492 (O_492,N_2983,N_2867);
or UO_493 (O_493,N_2823,N_2839);
nor UO_494 (O_494,N_2943,N_2935);
xor UO_495 (O_495,N_2884,N_2918);
or UO_496 (O_496,N_2914,N_2979);
xor UO_497 (O_497,N_2809,N_2800);
nor UO_498 (O_498,N_2868,N_2950);
xor UO_499 (O_499,N_2908,N_2996);
endmodule