module basic_1500_15000_2000_60_levels_2xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_1208,In_545);
and U1 (N_1,In_363,In_313);
and U2 (N_2,In_1388,In_1365);
or U3 (N_3,In_128,In_929);
and U4 (N_4,In_1477,In_639);
and U5 (N_5,In_1368,In_1154);
nand U6 (N_6,In_1246,In_856);
nor U7 (N_7,In_1138,In_346);
or U8 (N_8,In_329,In_1047);
or U9 (N_9,In_456,In_982);
or U10 (N_10,In_1226,In_1397);
and U11 (N_11,In_523,In_1189);
and U12 (N_12,In_719,In_315);
and U13 (N_13,In_890,In_349);
or U14 (N_14,In_1309,In_1006);
or U15 (N_15,In_692,In_861);
nand U16 (N_16,In_742,In_1143);
or U17 (N_17,In_538,In_828);
nand U18 (N_18,In_1360,In_498);
nor U19 (N_19,In_628,In_1135);
nor U20 (N_20,In_1450,In_940);
and U21 (N_21,In_995,In_761);
nor U22 (N_22,In_864,In_223);
nand U23 (N_23,In_948,In_829);
nand U24 (N_24,In_1499,In_1111);
nand U25 (N_25,In_801,In_426);
nand U26 (N_26,In_563,In_1324);
or U27 (N_27,In_731,In_808);
nor U28 (N_28,In_1392,In_720);
nand U29 (N_29,In_1056,In_1485);
nand U30 (N_30,In_521,In_1473);
and U31 (N_31,In_1380,In_832);
xor U32 (N_32,In_125,In_508);
nor U33 (N_33,In_875,In_1156);
or U34 (N_34,In_1093,In_1136);
or U35 (N_35,In_1005,In_863);
nor U36 (N_36,In_942,In_941);
and U37 (N_37,In_693,In_17);
nand U38 (N_38,In_705,In_1104);
nand U39 (N_39,In_500,In_499);
nand U40 (N_40,In_371,In_596);
or U41 (N_41,In_709,In_526);
nand U42 (N_42,In_542,In_320);
or U43 (N_43,In_1078,In_572);
and U44 (N_44,In_974,In_1417);
or U45 (N_45,In_484,In_25);
nor U46 (N_46,In_360,In_520);
or U47 (N_47,In_338,In_215);
nand U48 (N_48,In_1454,In_385);
and U49 (N_49,In_1086,In_1200);
and U50 (N_50,In_1446,In_454);
nor U51 (N_51,In_1455,In_1404);
nand U52 (N_52,In_253,In_522);
and U53 (N_53,In_1140,In_684);
or U54 (N_54,In_1002,In_1399);
nor U55 (N_55,In_785,In_568);
nand U56 (N_56,In_581,In_1354);
nand U57 (N_57,In_159,In_462);
nand U58 (N_58,In_886,In_778);
nand U59 (N_59,In_1031,In_840);
and U60 (N_60,In_1234,In_765);
xor U61 (N_61,In_1028,In_6);
or U62 (N_62,In_798,In_1306);
nand U63 (N_63,In_1277,In_656);
or U64 (N_64,In_1456,In_300);
nand U65 (N_65,In_431,In_1264);
and U66 (N_66,In_979,In_1307);
or U67 (N_67,In_584,In_347);
nand U68 (N_68,In_540,In_463);
nand U69 (N_69,In_1411,In_615);
and U70 (N_70,In_734,In_1459);
nand U71 (N_71,In_108,In_192);
nand U72 (N_72,In_1363,In_1290);
or U73 (N_73,In_1162,In_1339);
nand U74 (N_74,In_1438,In_1160);
and U75 (N_75,In_983,In_583);
or U76 (N_76,In_268,In_167);
and U77 (N_77,In_1487,In_1071);
and U78 (N_78,In_344,In_1118);
nand U79 (N_79,In_1284,In_473);
and U80 (N_80,In_1391,In_397);
nor U81 (N_81,In_551,In_851);
or U82 (N_82,In_968,In_988);
and U83 (N_83,In_891,In_562);
and U84 (N_84,In_123,In_1068);
or U85 (N_85,In_97,In_52);
nor U86 (N_86,In_809,In_303);
and U87 (N_87,In_477,In_1451);
xnor U88 (N_88,In_844,In_712);
or U89 (N_89,In_1225,In_1389);
nand U90 (N_90,In_670,In_1094);
and U91 (N_91,In_800,In_488);
or U92 (N_92,In_150,In_1345);
and U93 (N_93,In_920,In_47);
and U94 (N_94,In_603,In_39);
or U95 (N_95,In_737,In_241);
nor U96 (N_96,In_835,In_1466);
or U97 (N_97,In_117,In_365);
or U98 (N_98,In_298,In_1039);
and U99 (N_99,In_1432,In_1010);
nor U100 (N_100,In_1413,In_62);
nand U101 (N_101,In_1341,In_1132);
or U102 (N_102,In_55,In_1333);
nor U103 (N_103,In_1161,In_1030);
and U104 (N_104,In_28,In_779);
or U105 (N_105,In_502,In_1114);
or U106 (N_106,In_773,In_37);
or U107 (N_107,In_1350,In_1097);
nand U108 (N_108,In_1169,In_1175);
nor U109 (N_109,In_607,In_1270);
or U110 (N_110,In_814,In_435);
and U111 (N_111,In_725,In_304);
nor U112 (N_112,In_1149,In_1240);
nor U113 (N_113,In_683,In_1023);
and U114 (N_114,In_1322,In_513);
nor U115 (N_115,In_1167,In_357);
xor U116 (N_116,In_1362,In_1089);
or U117 (N_117,In_753,In_514);
xnor U118 (N_118,In_557,In_63);
nand U119 (N_119,In_86,In_222);
nor U120 (N_120,In_1045,In_1281);
and U121 (N_121,In_51,In_590);
nor U122 (N_122,In_1422,In_1124);
nor U123 (N_123,In_918,In_789);
and U124 (N_124,In_270,In_868);
or U125 (N_125,In_254,In_366);
nor U126 (N_126,In_1382,In_1106);
nand U127 (N_127,In_805,In_944);
or U128 (N_128,In_442,In_375);
nand U129 (N_129,In_361,In_1013);
and U130 (N_130,In_448,In_194);
and U131 (N_131,In_642,In_565);
nand U132 (N_132,In_1024,In_310);
and U133 (N_133,In_790,In_662);
nand U134 (N_134,In_962,In_1112);
xnor U135 (N_135,In_438,In_763);
and U136 (N_136,In_1427,In_978);
nand U137 (N_137,In_1332,In_1424);
nand U138 (N_138,In_493,In_700);
nand U139 (N_139,In_1077,In_73);
nand U140 (N_140,In_1107,In_322);
and U141 (N_141,In_959,In_611);
or U142 (N_142,In_1387,In_1130);
or U143 (N_143,In_1174,In_1458);
and U144 (N_144,In_1054,In_24);
and U145 (N_145,In_1445,In_393);
nand U146 (N_146,In_119,In_202);
nand U147 (N_147,In_876,In_1471);
or U148 (N_148,In_674,In_470);
nor U149 (N_149,In_1377,In_364);
or U150 (N_150,In_976,In_1295);
nor U151 (N_151,In_911,In_122);
and U152 (N_152,In_286,In_403);
nor U153 (N_153,In_1251,In_1479);
or U154 (N_154,In_1376,In_496);
nor U155 (N_155,In_1425,In_530);
nand U156 (N_156,In_193,In_1053);
and U157 (N_157,In_277,In_446);
and U158 (N_158,In_1117,In_199);
or U159 (N_159,In_1325,In_115);
nor U160 (N_160,In_923,In_1201);
and U161 (N_161,In_750,In_987);
or U162 (N_162,In_1082,In_850);
and U163 (N_163,In_695,In_782);
nor U164 (N_164,In_1063,In_296);
or U165 (N_165,In_955,In_291);
nand U166 (N_166,In_749,In_796);
or U167 (N_167,In_821,In_1032);
nand U168 (N_168,In_458,In_579);
or U169 (N_169,In_981,In_533);
or U170 (N_170,In_26,In_265);
nor U171 (N_171,In_90,In_612);
nor U172 (N_172,In_1249,In_101);
nand U173 (N_173,In_636,In_586);
nor U174 (N_174,In_998,In_707);
nand U175 (N_175,In_675,In_418);
nand U176 (N_176,In_339,In_627);
nand U177 (N_177,In_895,In_1492);
and U178 (N_178,In_149,In_299);
nand U179 (N_179,In_1034,In_1393);
nor U180 (N_180,In_1470,In_44);
and U181 (N_181,In_316,In_1493);
and U182 (N_182,In_260,In_135);
nand U183 (N_183,In_61,In_984);
and U184 (N_184,In_1357,In_1283);
nor U185 (N_185,In_387,In_1321);
or U186 (N_186,In_497,In_1462);
nand U187 (N_187,In_281,In_525);
or U188 (N_188,In_686,In_1179);
and U189 (N_189,In_1108,In_614);
nor U190 (N_190,In_1449,In_141);
or U191 (N_191,In_1057,In_921);
nor U192 (N_192,In_951,In_328);
and U193 (N_193,In_186,In_1323);
nand U194 (N_194,In_966,In_494);
nor U195 (N_195,In_1415,In_1308);
and U196 (N_196,In_218,In_587);
and U197 (N_197,In_384,In_818);
and U198 (N_198,In_871,In_174);
and U199 (N_199,In_532,In_757);
nand U200 (N_200,In_635,In_196);
and U201 (N_201,In_466,In_990);
and U202 (N_202,In_1434,In_1443);
nor U203 (N_203,In_495,In_931);
and U204 (N_204,In_593,In_893);
nand U205 (N_205,In_678,In_489);
nand U206 (N_206,In_114,In_973);
or U207 (N_207,In_263,In_1300);
nand U208 (N_208,In_820,In_843);
nand U209 (N_209,In_509,In_791);
or U210 (N_210,In_1352,In_716);
nand U211 (N_211,In_107,In_246);
nand U212 (N_212,In_696,In_608);
nor U213 (N_213,In_120,In_1369);
and U214 (N_214,In_1441,In_345);
and U215 (N_215,In_1334,In_118);
or U216 (N_216,In_1199,In_439);
nand U217 (N_217,In_1159,In_985);
nor U218 (N_218,In_297,In_578);
nor U219 (N_219,In_585,In_155);
and U220 (N_220,In_837,In_162);
and U221 (N_221,In_1347,In_802);
nor U222 (N_222,In_666,In_130);
and U223 (N_223,In_145,In_1327);
and U224 (N_224,In_516,In_331);
nand U225 (N_225,In_20,In_680);
and U226 (N_226,In_306,In_1266);
nand U227 (N_227,In_1361,In_434);
nand U228 (N_228,In_208,In_48);
and U229 (N_229,In_374,In_1280);
nor U230 (N_230,In_916,In_1469);
or U231 (N_231,In_710,In_838);
nor U232 (N_232,In_1355,In_225);
nor U233 (N_233,In_970,In_354);
nand U234 (N_234,In_899,In_652);
nor U235 (N_235,In_410,In_474);
nor U236 (N_236,In_1440,In_566);
nand U237 (N_237,In_1285,In_1095);
nor U238 (N_238,In_877,In_1027);
and U239 (N_239,In_836,In_1085);
and U240 (N_240,In_478,In_659);
xnor U241 (N_241,In_278,In_1079);
nor U242 (N_242,In_592,In_1405);
or U243 (N_243,In_1131,In_146);
nand U244 (N_244,In_1273,In_834);
or U245 (N_245,In_232,In_904);
or U246 (N_246,In_730,In_274);
or U247 (N_247,In_950,In_799);
or U248 (N_248,In_1489,In_792);
nor U249 (N_249,In_243,In_53);
or U250 (N_250,In_394,In_482);
nand U251 (N_251,N_153,N_249);
nand U252 (N_252,In_1409,In_164);
nand U253 (N_253,In_571,In_401);
nand U254 (N_254,In_109,In_70);
nand U255 (N_255,In_370,In_1435);
xor U256 (N_256,In_1315,N_29);
nand U257 (N_257,In_351,In_867);
nor U258 (N_258,In_65,In_846);
nand U259 (N_259,In_913,N_81);
and U260 (N_260,In_43,In_1292);
or U261 (N_261,In_1069,In_1074);
and U262 (N_262,In_423,In_112);
and U263 (N_263,In_1457,In_1326);
nand U264 (N_264,In_1330,In_1491);
nor U265 (N_265,In_175,In_1364);
nor U266 (N_266,In_1172,In_134);
nand U267 (N_267,In_142,In_632);
or U268 (N_268,N_193,In_945);
or U269 (N_269,In_250,In_810);
nand U270 (N_270,In_217,In_84);
nand U271 (N_271,In_244,In_546);
and U272 (N_272,In_391,In_1373);
nor U273 (N_273,In_986,In_1168);
or U274 (N_274,N_229,In_1171);
nor U275 (N_275,N_126,In_881);
and U276 (N_276,In_755,In_667);
and U277 (N_277,In_768,In_1142);
nand U278 (N_278,In_885,In_87);
nand U279 (N_279,In_342,In_1206);
and U280 (N_280,N_56,In_859);
and U281 (N_281,In_631,In_1119);
and U282 (N_282,In_1188,In_637);
and U283 (N_283,N_125,In_511);
nand U284 (N_284,In_884,In_1298);
or U285 (N_285,In_946,In_1163);
xnor U286 (N_286,In_902,N_103);
or U287 (N_287,In_177,In_855);
nand U288 (N_288,In_1060,In_1213);
or U289 (N_289,In_714,In_152);
xnor U290 (N_290,In_564,In_616);
or U291 (N_291,In_599,In_415);
nor U292 (N_292,In_273,In_1239);
nand U293 (N_293,In_78,N_36);
and U294 (N_294,In_404,In_132);
and U295 (N_295,N_182,In_1379);
nand U296 (N_296,In_234,In_1328);
nor U297 (N_297,In_1312,In_1205);
nor U298 (N_298,In_251,N_12);
and U299 (N_299,In_503,In_433);
and U300 (N_300,N_236,In_1083);
nand U301 (N_301,In_770,In_219);
and U302 (N_302,In_1,In_949);
nand U303 (N_303,In_1252,In_957);
nor U304 (N_304,In_623,In_266);
or U305 (N_305,In_455,In_327);
and U306 (N_306,In_29,In_34);
nor U307 (N_307,In_9,In_1180);
xnor U308 (N_308,In_704,In_1040);
and U309 (N_309,In_994,N_49);
nand U310 (N_310,In_823,In_75);
and U311 (N_311,N_232,N_119);
nor U312 (N_312,In_421,N_231);
or U313 (N_313,In_788,In_1406);
and U314 (N_314,In_292,N_108);
nor U315 (N_315,In_172,N_85);
or U316 (N_316,N_190,In_919);
nor U317 (N_317,In_558,N_166);
or U318 (N_318,N_3,In_1091);
or U319 (N_319,In_491,In_336);
and U320 (N_320,In_870,In_335);
and U321 (N_321,In_77,In_826);
nand U322 (N_322,In_1288,In_967);
nor U323 (N_323,In_103,N_104);
and U324 (N_324,In_379,In_1297);
nand U325 (N_325,In_181,In_42);
or U326 (N_326,In_928,In_325);
or U327 (N_327,N_110,N_170);
nor U328 (N_328,In_227,N_1);
nor U329 (N_329,In_582,N_226);
and U330 (N_330,N_169,In_1497);
and U331 (N_331,In_515,In_965);
or U332 (N_332,In_728,In_643);
and U333 (N_333,In_248,In_1222);
nor U334 (N_334,In_262,N_39);
and U335 (N_335,In_58,In_204);
and U336 (N_336,In_781,N_227);
nor U337 (N_337,In_408,In_1099);
or U338 (N_338,N_53,N_149);
and U339 (N_339,In_1049,N_130);
or U340 (N_340,In_89,In_348);
nor U341 (N_341,In_191,In_386);
nand U342 (N_342,In_673,In_1467);
nor U343 (N_343,In_203,N_142);
or U344 (N_344,In_852,In_280);
or U345 (N_345,In_68,N_102);
and U346 (N_346,In_355,In_72);
and U347 (N_347,In_1113,In_302);
nand U348 (N_348,N_38,In_909);
and U349 (N_349,In_595,In_1088);
and U350 (N_350,In_560,N_44);
nor U351 (N_351,In_685,In_1311);
and U352 (N_352,In_567,In_690);
nor U353 (N_353,In_1029,In_92);
and U354 (N_354,In_1274,In_897);
and U355 (N_355,N_105,In_486);
or U356 (N_356,In_1204,In_1148);
nand U357 (N_357,N_148,In_189);
and U358 (N_358,In_570,N_222);
or U359 (N_359,In_57,N_192);
and U360 (N_360,N_189,In_179);
nand U361 (N_361,N_160,In_747);
nand U362 (N_362,In_1367,In_1007);
and U363 (N_363,In_736,In_1102);
or U364 (N_364,In_1058,In_943);
xnor U365 (N_365,In_1145,In_1395);
or U366 (N_366,In_519,In_1253);
and U367 (N_367,In_432,In_399);
nand U368 (N_368,In_334,In_771);
nand U369 (N_369,In_1176,In_934);
nand U370 (N_370,In_1242,In_447);
or U371 (N_371,In_1337,N_186);
nand U372 (N_372,In_190,In_1052);
nand U373 (N_373,In_1202,In_16);
or U374 (N_374,In_343,In_769);
or U375 (N_375,In_975,In_1016);
and U376 (N_376,In_718,In_1394);
or U377 (N_377,In_549,In_318);
and U378 (N_378,In_1262,In_1316);
nor U379 (N_379,In_1084,N_176);
and U380 (N_380,In_723,In_527);
and U381 (N_381,In_660,In_1408);
nor U382 (N_382,In_1123,In_210);
and U383 (N_383,In_1258,In_1268);
xnor U384 (N_384,In_1439,In_472);
or U385 (N_385,In_59,In_1139);
nand U386 (N_386,In_479,In_839);
nand U387 (N_387,N_15,In_1155);
nand U388 (N_388,In_989,N_201);
nand U389 (N_389,N_30,In_668);
nand U390 (N_390,In_517,In_1259);
and U391 (N_391,In_1335,N_70);
nor U392 (N_392,In_409,In_849);
and U393 (N_393,N_99,In_15);
nor U394 (N_394,In_293,In_738);
nand U395 (N_395,In_38,In_1320);
or U396 (N_396,In_1317,N_111);
or U397 (N_397,N_86,N_42);
or U398 (N_398,In_10,In_854);
xnor U399 (N_399,In_926,In_535);
nand U400 (N_400,N_181,In_997);
and U401 (N_401,N_74,In_443);
nand U402 (N_402,In_170,In_1375);
nor U403 (N_403,In_857,N_187);
nand U404 (N_404,In_767,In_1064);
nand U405 (N_405,In_1418,In_1051);
nand U406 (N_406,N_247,In_996);
and U407 (N_407,In_461,N_155);
nor U408 (N_408,N_107,In_1025);
nor U409 (N_409,In_312,In_137);
and U410 (N_410,In_294,N_173);
nor U411 (N_411,In_275,In_60);
nand U412 (N_412,In_883,N_67);
and U413 (N_413,In_157,N_89);
or U414 (N_414,In_41,In_1353);
nand U415 (N_415,In_12,In_1150);
or U416 (N_416,In_79,In_264);
nand U417 (N_417,In_1046,In_206);
or U418 (N_418,In_402,N_118);
or U419 (N_419,N_14,In_784);
nand U420 (N_420,In_681,In_598);
or U421 (N_421,In_452,In_1233);
nor U422 (N_422,N_138,In_597);
nand U423 (N_423,In_213,N_159);
nor U424 (N_424,In_317,In_419);
xnor U425 (N_425,In_694,In_780);
or U426 (N_426,N_100,In_1314);
nand U427 (N_427,In_436,In_21);
or U428 (N_428,N_143,In_1182);
nor U429 (N_429,In_156,In_400);
nand U430 (N_430,In_200,In_414);
and U431 (N_431,N_146,In_1127);
or U432 (N_432,In_441,In_703);
or U433 (N_433,N_233,In_1190);
nand U434 (N_434,In_269,In_676);
or U435 (N_435,N_195,N_242);
nor U436 (N_436,In_613,In_480);
nand U437 (N_437,In_127,In_552);
and U438 (N_438,In_764,In_732);
nor U439 (N_439,In_2,In_1336);
nand U440 (N_440,In_1291,N_124);
and U441 (N_441,In_209,In_661);
and U442 (N_442,In_1444,N_180);
and U443 (N_443,In_879,N_127);
nor U444 (N_444,In_187,In_900);
and U445 (N_445,N_208,In_1230);
and U446 (N_446,In_1217,In_464);
or U447 (N_447,In_717,In_23);
xnor U448 (N_448,N_52,In_610);
nand U449 (N_449,N_31,In_13);
nand U450 (N_450,In_1228,In_618);
nand U451 (N_451,N_51,In_1236);
and U452 (N_452,N_71,N_234);
xor U453 (N_453,In_104,In_367);
or U454 (N_454,N_194,In_1048);
nor U455 (N_455,In_912,In_425);
and U456 (N_456,In_1196,N_140);
and U457 (N_457,In_1478,In_759);
xor U458 (N_458,N_79,N_235);
nand U459 (N_459,In_1223,In_1126);
and U460 (N_460,N_152,In_1219);
or U461 (N_461,In_1214,N_225);
and U462 (N_462,In_1100,In_1000);
or U463 (N_463,In_1338,In_1460);
nor U464 (N_464,In_1301,In_359);
and U465 (N_465,In_787,In_163);
or U466 (N_466,In_368,In_501);
and U467 (N_467,In_139,In_953);
xnor U468 (N_468,In_1304,N_240);
nand U469 (N_469,In_1423,In_350);
and U470 (N_470,In_381,In_1194);
nand U471 (N_471,In_467,In_76);
nor U472 (N_472,In_589,In_547);
nor U473 (N_473,In_847,In_252);
nand U474 (N_474,In_1157,In_1310);
nand U475 (N_475,In_11,In_138);
nand U476 (N_476,In_1019,In_963);
nor U477 (N_477,In_93,N_122);
nor U478 (N_478,N_179,N_59);
nand U479 (N_479,In_289,In_766);
or U480 (N_480,In_1475,In_775);
nand U481 (N_481,In_1381,In_1015);
nand U482 (N_482,In_556,N_230);
nor U483 (N_483,In_1426,In_45);
or U484 (N_484,In_326,In_153);
and U485 (N_485,In_842,In_1279);
or U486 (N_486,In_624,N_114);
and U487 (N_487,In_812,In_935);
nand U488 (N_488,In_947,In_288);
nor U489 (N_489,N_244,In_151);
or U490 (N_490,In_183,In_1203);
or U491 (N_491,In_1125,In_468);
or U492 (N_492,In_3,In_1390);
nand U493 (N_493,In_1076,In_301);
or U494 (N_494,In_1191,In_116);
and U495 (N_495,In_195,N_207);
nand U496 (N_496,In_641,N_75);
and U497 (N_497,In_1416,In_762);
and U498 (N_498,N_174,N_238);
nand U499 (N_499,In_860,N_72);
nand U500 (N_500,N_168,In_362);
or U501 (N_501,N_256,In_64);
nor U502 (N_502,N_129,In_481);
and U503 (N_503,N_325,In_650);
or U504 (N_504,N_498,In_569);
or U505 (N_505,In_960,In_1488);
or U506 (N_506,In_1141,N_396);
nand U507 (N_507,In_1216,In_1173);
nand U508 (N_508,In_1062,N_422);
nand U509 (N_509,In_444,N_395);
nand U510 (N_510,In_1366,In_740);
and U511 (N_511,N_477,In_1134);
or U512 (N_512,In_1181,In_1192);
and U513 (N_513,In_311,In_475);
or U514 (N_514,In_110,N_183);
nor U515 (N_515,In_358,N_19);
nand U516 (N_516,In_233,In_83);
nor U517 (N_517,N_454,N_447);
or U518 (N_518,In_617,In_405);
nand U519 (N_519,In_111,In_305);
and U520 (N_520,N_281,In_1043);
or U521 (N_521,In_952,N_414);
nand U522 (N_522,N_254,N_94);
and U523 (N_523,N_315,N_18);
nand U524 (N_524,N_48,In_460);
or U525 (N_525,N_175,N_445);
nand U526 (N_526,N_6,In_1463);
nand U527 (N_527,In_848,In_1021);
nand U528 (N_528,In_82,N_434);
xor U529 (N_529,In_231,In_910);
and U530 (N_530,N_339,N_449);
nand U531 (N_531,N_76,In_930);
and U532 (N_532,N_37,In_588);
and U533 (N_533,In_216,N_210);
or U534 (N_534,In_1067,N_453);
and U535 (N_535,In_553,In_1476);
xor U536 (N_536,In_185,In_756);
and U537 (N_537,In_1014,In_644);
nand U538 (N_538,In_698,N_496);
nor U539 (N_539,N_215,In_869);
nor U540 (N_540,In_437,N_369);
nor U541 (N_541,In_1044,In_36);
nand U542 (N_542,N_112,In_417);
nor U543 (N_543,In_1374,In_284);
or U544 (N_544,N_115,N_20);
nand U545 (N_545,In_1461,In_49);
nand U546 (N_546,N_465,In_98);
nand U547 (N_547,N_161,N_471);
nand U548 (N_548,N_352,N_224);
and U549 (N_549,N_408,In_14);
and U550 (N_550,N_144,In_74);
or U551 (N_551,In_1420,N_459);
nand U552 (N_552,N_337,N_484);
and U553 (N_553,N_332,N_277);
or U554 (N_554,In_548,In_1371);
and U555 (N_555,In_806,N_318);
nor U556 (N_556,N_415,In_54);
or U557 (N_557,In_1185,N_172);
nand U558 (N_558,In_543,N_432);
nor U559 (N_559,In_971,In_154);
nand U560 (N_560,In_201,In_748);
nand U561 (N_561,N_397,In_131);
nand U562 (N_562,In_182,N_24);
or U563 (N_563,N_316,N_188);
nor U564 (N_564,In_1319,In_715);
and U565 (N_565,In_198,In_729);
or U566 (N_566,In_671,In_276);
nand U567 (N_567,In_819,In_892);
and U568 (N_568,N_317,In_121);
and U569 (N_569,In_4,In_746);
or U570 (N_570,N_62,N_421);
nand U571 (N_571,N_402,In_1229);
and U572 (N_572,N_109,In_1209);
and U573 (N_573,N_329,N_248);
nor U574 (N_574,N_394,In_999);
and U575 (N_575,In_1147,N_295);
nor U576 (N_576,N_45,In_1260);
and U577 (N_577,N_268,N_426);
nand U578 (N_578,In_908,N_286);
or U579 (N_579,In_898,N_58);
nor U580 (N_580,In_295,In_1278);
nor U581 (N_581,In_831,N_483);
nand U582 (N_582,In_880,In_1359);
and U583 (N_583,N_346,In_1495);
and U584 (N_584,In_309,In_1221);
and U585 (N_585,In_1263,N_458);
nor U586 (N_586,N_360,In_412);
nor U587 (N_587,N_150,In_1087);
or U588 (N_588,N_391,N_185);
or U589 (N_589,In_240,N_17);
or U590 (N_590,N_425,In_100);
nand U591 (N_591,In_324,In_786);
nor U592 (N_592,In_938,In_1358);
nand U593 (N_593,In_1401,N_451);
or U594 (N_594,N_2,In_554);
nand U595 (N_595,In_372,In_711);
nor U596 (N_596,N_485,In_449);
and U597 (N_597,N_265,In_845);
and U598 (N_598,N_243,In_81);
nor U599 (N_599,N_353,In_657);
and U600 (N_600,In_1096,N_23);
or U601 (N_601,N_211,In_922);
nand U602 (N_602,In_1286,N_213);
or U603 (N_603,In_95,N_384);
or U604 (N_604,N_43,N_78);
nor U605 (N_605,In_1122,N_272);
nand U606 (N_606,In_1340,In_972);
xnor U607 (N_607,N_418,In_258);
nand U608 (N_608,N_223,N_25);
nand U609 (N_609,In_722,In_245);
and U610 (N_610,In_754,In_1215);
nor U611 (N_611,N_91,In_144);
xnor U612 (N_612,In_529,In_862);
nand U613 (N_613,In_1498,In_625);
nor U614 (N_614,N_263,In_380);
or U615 (N_615,N_209,In_1407);
nand U616 (N_616,In_713,In_1305);
or U617 (N_617,In_888,In_1486);
nor U618 (N_618,In_1346,N_488);
or U619 (N_619,N_64,N_375);
nor U620 (N_620,In_422,In_469);
and U621 (N_621,In_212,In_804);
nand U622 (N_622,N_252,N_216);
or U623 (N_623,N_361,N_139);
and U624 (N_624,N_377,In_314);
or U625 (N_625,In_825,In_143);
nand U626 (N_626,In_1020,In_451);
nand U627 (N_627,N_264,N_26);
nand U628 (N_628,In_106,In_230);
and U629 (N_629,N_164,N_0);
nand U630 (N_630,In_1433,N_8);
and U631 (N_631,N_294,N_492);
and U632 (N_632,N_357,In_369);
or U633 (N_633,In_1403,N_178);
or U634 (N_634,N_101,In_382);
and U635 (N_635,In_777,In_88);
and U636 (N_636,N_301,In_356);
or U637 (N_637,N_203,In_776);
nor U638 (N_638,In_691,N_269);
nor U639 (N_639,In_1081,In_440);
and U640 (N_640,N_288,In_858);
nor U641 (N_641,In_1245,N_393);
or U642 (N_642,In_701,N_433);
and U643 (N_643,In_1303,N_307);
nor U644 (N_644,N_7,In_133);
xor U645 (N_645,N_366,In_1244);
or U646 (N_646,N_333,In_1022);
nand U647 (N_647,In_1080,In_259);
and U648 (N_648,In_1329,In_99);
nor U649 (N_649,N_276,In_50);
nand U650 (N_650,N_350,In_609);
or U651 (N_651,In_697,N_372);
nand U652 (N_652,In_993,In_1421);
nor U653 (N_653,N_334,N_310);
nor U654 (N_654,N_359,N_162);
nor U655 (N_655,In_31,N_84);
nor U656 (N_656,N_311,In_518);
or U657 (N_657,In_1276,In_457);
nor U658 (N_658,N_57,In_1255);
xor U659 (N_659,N_431,In_1009);
nand U660 (N_660,N_260,In_573);
or U661 (N_661,N_378,N_167);
nand U662 (N_662,N_406,N_499);
nand U663 (N_663,N_61,In_1004);
or U664 (N_664,In_1452,In_465);
nor U665 (N_665,In_505,In_665);
nor U666 (N_666,N_98,In_158);
and U667 (N_667,N_371,N_219);
nand U668 (N_668,N_305,In_574);
nor U669 (N_669,N_368,N_13);
nor U670 (N_670,N_482,N_428);
nand U671 (N_671,In_229,N_171);
nand U672 (N_672,N_448,N_338);
nor U673 (N_673,N_47,In_169);
and U674 (N_674,N_218,In_648);
or U675 (N_675,In_272,In_430);
nor U676 (N_676,In_424,N_60);
nor U677 (N_677,N_135,N_355);
or U678 (N_678,In_224,In_1496);
or U679 (N_679,N_312,In_396);
nor U680 (N_680,In_383,In_1267);
or U681 (N_681,In_816,In_1494);
nor U682 (N_682,In_180,N_380);
and U683 (N_683,N_356,N_92);
and U684 (N_684,In_807,N_494);
and U685 (N_685,In_1059,In_677);
nand U686 (N_686,N_340,N_306);
nand U687 (N_687,In_992,N_293);
nor U688 (N_688,In_964,In_905);
nand U689 (N_689,In_173,N_95);
or U690 (N_690,In_353,In_1247);
nor U691 (N_691,N_34,In_450);
or U692 (N_692,In_654,N_399);
or U693 (N_693,In_492,In_878);
nand U694 (N_694,In_1207,N_370);
or U695 (N_695,N_489,In_471);
xnor U696 (N_696,In_866,N_478);
nand U697 (N_697,In_420,In_1098);
nor U698 (N_698,N_96,In_903);
or U699 (N_699,In_774,In_961);
nor U700 (N_700,In_794,N_141);
nand U701 (N_701,N_11,In_1349);
or U702 (N_702,N_486,N_320);
or U703 (N_703,In_0,N_466);
or U704 (N_704,In_165,In_22);
and U705 (N_705,N_21,N_5);
nand U706 (N_706,In_1003,N_351);
nor U707 (N_707,N_376,In_407);
or U708 (N_708,In_188,N_358);
nor U709 (N_709,N_237,In_1152);
or U710 (N_710,N_476,In_506);
nand U711 (N_711,In_1256,In_124);
nor U712 (N_712,In_1248,In_214);
and U713 (N_713,N_438,In_679);
nor U714 (N_714,In_46,N_284);
xnor U715 (N_715,In_1356,In_1195);
or U716 (N_716,N_65,In_1115);
and U717 (N_717,In_1158,N_267);
or U718 (N_718,In_1110,N_364);
or U719 (N_719,N_324,In_333);
and U720 (N_720,In_1133,In_1447);
nand U721 (N_721,In_321,N_120);
and U722 (N_722,N_349,In_490);
and U723 (N_723,In_32,In_865);
nor U724 (N_724,In_1414,N_28);
nor U725 (N_725,In_1254,N_322);
and U726 (N_726,In_682,In_1116);
nand U727 (N_727,In_1128,In_933);
nor U728 (N_728,N_151,N_417);
and U729 (N_729,In_969,In_932);
or U730 (N_730,In_1105,In_739);
or U731 (N_731,N_410,In_1250);
nor U732 (N_732,In_751,In_282);
nor U733 (N_733,In_1121,In_833);
and U734 (N_734,N_83,In_319);
nor U735 (N_735,N_354,In_102);
nand U736 (N_736,In_1429,In_1035);
and U737 (N_737,In_1269,N_16);
or U738 (N_738,In_1101,In_824);
nand U739 (N_739,In_1061,N_257);
xor U740 (N_740,N_419,In_395);
nand U741 (N_741,In_1066,In_271);
and U742 (N_742,In_5,In_80);
nand U743 (N_743,In_30,In_629);
and U744 (N_744,In_1484,In_140);
nor U745 (N_745,In_1026,In_1342);
nand U746 (N_746,In_7,In_1055);
nand U747 (N_747,N_467,In_221);
nand U748 (N_748,In_1235,In_69);
nor U749 (N_749,In_337,N_132);
or U750 (N_750,N_68,In_184);
nor U751 (N_751,N_409,N_740);
and U752 (N_752,N_572,N_666);
nand U753 (N_753,N_693,In_872);
nand U754 (N_754,In_663,N_570);
nor U755 (N_755,N_435,N_493);
and U756 (N_756,In_783,N_479);
nor U757 (N_757,N_335,N_626);
nand U758 (N_758,N_596,N_574);
or U759 (N_759,N_270,In_1187);
nor U760 (N_760,N_163,N_594);
and U761 (N_761,N_323,N_695);
or U762 (N_762,N_620,N_562);
nor U763 (N_763,In_1400,N_382);
or U764 (N_764,N_536,N_627);
and U765 (N_765,In_561,N_46);
nor U766 (N_766,In_483,In_594);
and U767 (N_767,N_722,N_581);
nand U768 (N_768,In_56,In_1237);
nand U769 (N_769,In_1184,N_551);
nand U770 (N_770,N_670,N_713);
nand U771 (N_771,In_958,In_249);
nor U772 (N_772,In_619,N_654);
nor U773 (N_773,In_874,In_176);
nand U774 (N_774,In_1383,In_290);
and U775 (N_775,N_196,N_158);
nand U776 (N_776,N_663,N_689);
nand U777 (N_777,N_633,N_720);
nor U778 (N_778,N_487,In_803);
or U779 (N_779,In_1398,N_582);
nor U780 (N_780,In_1351,N_735);
nor U781 (N_781,N_724,In_1033);
or U782 (N_782,N_711,N_212);
nand U783 (N_783,In_745,N_560);
or U784 (N_784,N_446,N_480);
or U785 (N_785,N_253,In_689);
and U786 (N_786,N_652,N_495);
nor U787 (N_787,N_259,N_610);
nand U788 (N_788,N_676,In_1198);
or U789 (N_789,N_512,N_10);
nor U790 (N_790,N_398,N_748);
nand U791 (N_791,N_688,N_539);
and U792 (N_792,In_1299,In_1017);
and U793 (N_793,N_66,In_459);
and U794 (N_794,N_113,In_33);
xnor U795 (N_795,N_401,N_714);
nand U796 (N_796,N_621,N_653);
and U797 (N_797,N_412,In_936);
nand U798 (N_798,In_1243,N_535);
nand U799 (N_799,N_643,In_1072);
nor U800 (N_800,N_374,N_623);
or U801 (N_801,N_440,In_917);
and U802 (N_802,N_747,N_734);
and U803 (N_803,N_647,N_228);
and U804 (N_804,N_439,N_522);
nor U805 (N_805,N_658,N_456);
nor U806 (N_806,N_93,In_1227);
or U807 (N_807,In_1490,In_487);
and U808 (N_808,In_1448,N_514);
or U809 (N_809,In_1465,In_1442);
and U810 (N_810,N_634,N_586);
and U811 (N_811,In_1293,N_661);
nor U812 (N_812,N_664,In_620);
nor U813 (N_813,N_615,N_441);
or U814 (N_814,In_330,In_1065);
xor U815 (N_815,In_724,In_925);
xor U816 (N_816,In_27,In_822);
nor U817 (N_817,In_752,In_1436);
or U818 (N_818,In_1294,N_733);
nand U819 (N_819,N_404,N_157);
and U820 (N_820,In_1075,N_423);
or U821 (N_821,N_255,N_199);
and U822 (N_822,In_389,N_655);
nor U823 (N_823,In_416,N_745);
nor U824 (N_824,N_386,N_690);
nand U825 (N_825,N_565,In_1343);
nor U826 (N_826,In_261,N_575);
nor U827 (N_827,N_497,N_552);
or U828 (N_828,N_200,In_772);
and U829 (N_829,N_579,N_90);
nand U830 (N_830,In_1372,In_129);
nand U831 (N_831,In_1385,N_573);
nor U832 (N_832,In_1231,N_662);
or U833 (N_833,In_332,N_667);
nand U834 (N_834,In_1178,N_413);
nand U835 (N_835,In_601,In_373);
or U836 (N_836,In_1164,N_541);
nor U837 (N_837,N_283,N_650);
and U838 (N_838,N_22,N_279);
nor U839 (N_839,N_80,In_1193);
nand U840 (N_840,N_721,N_612);
nand U841 (N_841,N_591,In_544);
nor U842 (N_842,N_282,N_603);
or U843 (N_843,In_664,N_385);
nand U844 (N_844,N_692,In_1431);
or U845 (N_845,N_569,In_1018);
and U846 (N_846,N_258,N_526);
or U847 (N_847,N_500,N_33);
or U848 (N_848,N_698,N_702);
nand U849 (N_849,In_1313,N_639);
nor U850 (N_850,In_602,N_624);
nor U851 (N_851,N_55,N_595);
nor U852 (N_852,N_297,N_668);
or U853 (N_853,N_473,In_1090);
and U854 (N_854,In_429,In_1129);
nand U855 (N_855,N_275,In_1177);
nand U856 (N_856,N_629,N_345);
nor U857 (N_857,In_699,N_450);
nand U858 (N_858,In_937,In_980);
and U859 (N_859,In_797,In_147);
nand U860 (N_860,In_352,N_642);
nand U861 (N_861,N_580,In_647);
nand U862 (N_862,In_485,N_558);
and U863 (N_863,N_608,In_18);
nor U864 (N_864,In_1483,In_605);
nor U865 (N_865,In_827,N_604);
nor U866 (N_866,N_468,In_646);
nor U867 (N_867,In_1186,N_429);
nor U868 (N_868,In_537,In_1287);
and U869 (N_869,N_88,In_1302);
and U870 (N_870,N_469,In_977);
nor U871 (N_871,N_326,In_622);
or U872 (N_872,N_470,In_1480);
nand U873 (N_873,In_1275,N_730);
nor U874 (N_874,In_1344,N_716);
nor U875 (N_875,In_793,In_8);
nor U876 (N_876,N_527,N_602);
or U877 (N_877,In_392,In_411);
nand U878 (N_878,N_533,N_736);
and U879 (N_879,In_1468,In_1144);
and U880 (N_880,In_1428,N_553);
nand U881 (N_881,N_121,N_50);
and U882 (N_882,In_171,N_544);
nor U883 (N_883,N_381,N_137);
nand U884 (N_884,N_563,N_327);
and U885 (N_885,N_308,N_532);
and U886 (N_886,N_274,N_640);
nor U887 (N_887,In_604,In_853);
and U888 (N_888,N_35,N_638);
nor U889 (N_889,N_600,In_1137);
and U890 (N_890,In_1272,N_217);
nor U891 (N_891,N_675,In_1153);
or U892 (N_892,N_519,N_645);
nor U893 (N_893,In_927,N_221);
and U894 (N_894,N_529,N_681);
xnor U895 (N_895,N_266,N_707);
or U896 (N_896,In_1041,N_660);
nand U897 (N_897,N_490,N_584);
or U898 (N_898,In_1464,N_246);
nor U899 (N_899,N_649,In_283);
and U900 (N_900,N_475,In_228);
and U901 (N_901,In_1348,In_19);
nand U902 (N_902,In_896,N_696);
and U903 (N_903,In_105,N_136);
nand U904 (N_904,N_299,In_815);
nor U905 (N_905,N_723,N_708);
or U906 (N_906,N_509,N_147);
and U907 (N_907,N_619,N_717);
and U908 (N_908,In_1042,In_1038);
nand U909 (N_909,In_247,In_887);
nor U910 (N_910,In_649,N_705);
nand U911 (N_911,In_220,In_341);
and U912 (N_912,N_592,N_69);
nand U913 (N_913,In_507,N_641);
or U914 (N_914,In_94,N_564);
nand U915 (N_915,In_1241,N_197);
nand U916 (N_916,N_133,N_285);
and U917 (N_917,N_328,In_901);
and U918 (N_918,N_697,In_376);
or U919 (N_919,N_191,N_715);
or U920 (N_920,N_607,In_841);
nand U921 (N_921,In_197,In_555);
nand U922 (N_922,In_640,N_727);
and U923 (N_923,N_644,In_66);
nor U924 (N_924,N_296,N_87);
nor U925 (N_925,In_760,In_1073);
xor U926 (N_926,In_915,N_726);
or U927 (N_927,N_463,N_403);
or U928 (N_928,N_672,In_1070);
nor U929 (N_929,N_452,In_161);
nand U930 (N_930,N_491,N_206);
and U931 (N_931,In_1224,In_817);
or U932 (N_932,In_238,N_289);
xnor U933 (N_933,N_712,In_528);
nand U934 (N_934,In_1001,N_342);
and U935 (N_935,In_1282,N_348);
or U936 (N_936,N_32,In_1296);
nor U937 (N_937,N_184,N_290);
nor U938 (N_938,In_1410,In_453);
or U939 (N_939,N_550,In_1036);
nand U940 (N_940,N_749,N_204);
xnor U941 (N_941,N_525,N_543);
nor U942 (N_942,N_617,N_77);
nor U943 (N_943,N_4,In_67);
nor U944 (N_944,N_576,N_568);
and U945 (N_945,In_1453,N_220);
or U946 (N_946,N_388,In_136);
nand U947 (N_947,In_1378,N_513);
and U948 (N_948,In_1474,N_508);
and U949 (N_949,N_379,N_518);
nor U950 (N_950,N_321,In_889);
and U951 (N_951,N_743,N_362);
and U952 (N_952,In_160,In_939);
nor U953 (N_953,N_630,N_411);
and U954 (N_954,N_515,N_154);
and U955 (N_955,In_655,N_251);
nor U956 (N_956,In_906,N_442);
and U957 (N_957,In_308,In_1120);
or U958 (N_958,In_882,In_427);
and U959 (N_959,In_621,In_669);
nor U960 (N_960,In_924,N_462);
and U961 (N_961,N_738,In_830);
nor U962 (N_962,In_873,In_524);
or U963 (N_963,In_1165,N_40);
nand U964 (N_964,In_1146,N_117);
or U965 (N_965,N_506,N_673);
nor U966 (N_966,N_566,N_202);
nand U967 (N_967,N_545,In_559);
nor U968 (N_968,In_510,N_648);
nand U969 (N_969,N_646,N_656);
and U970 (N_970,N_389,N_504);
nand U971 (N_971,N_686,In_658);
and U972 (N_972,N_436,In_256);
or U973 (N_973,N_63,N_241);
or U974 (N_974,N_347,In_377);
nand U975 (N_975,N_367,N_737);
and U976 (N_976,In_504,In_991);
nand U977 (N_977,N_742,In_71);
or U978 (N_978,In_390,N_319);
and U979 (N_979,N_444,N_671);
nand U980 (N_980,In_1103,N_416);
nand U981 (N_981,In_1331,In_907);
and U982 (N_982,N_387,N_145);
nand U983 (N_983,N_651,N_198);
xor U984 (N_984,In_1011,N_637);
or U985 (N_985,In_536,In_476);
nand U986 (N_986,In_914,In_626);
nand U987 (N_987,N_505,In_706);
or U988 (N_988,N_392,In_1370);
nor U989 (N_989,In_688,In_576);
and U990 (N_990,N_549,N_622);
and U991 (N_991,N_588,N_701);
and U992 (N_992,In_1289,N_239);
and U993 (N_993,N_177,In_744);
and U994 (N_994,N_691,In_1232);
or U995 (N_995,In_1218,N_593);
and U996 (N_996,N_511,In_35);
and U997 (N_997,N_390,N_273);
nand U998 (N_998,N_344,N_632);
and U999 (N_999,N_82,In_687);
nor U1000 (N_1000,N_280,In_428);
nand U1001 (N_1001,N_775,N_945);
and U1002 (N_1002,In_413,In_645);
nor U1003 (N_1003,N_287,N_810);
and U1004 (N_1004,In_733,N_894);
and U1005 (N_1005,In_285,In_91);
or U1006 (N_1006,N_474,In_956);
nor U1007 (N_1007,In_1220,N_933);
or U1008 (N_1008,N_920,In_653);
or U1009 (N_1009,N_540,N_41);
nand U1010 (N_1010,N_719,N_261);
nor U1011 (N_1011,N_771,N_457);
or U1012 (N_1012,N_802,In_166);
nor U1013 (N_1013,In_1257,In_378);
and U1014 (N_1014,N_903,N_782);
or U1015 (N_1015,N_801,In_307);
or U1016 (N_1016,N_9,N_599);
and U1017 (N_1017,N_868,N_165);
or U1018 (N_1018,N_985,N_537);
nor U1019 (N_1019,In_1261,N_878);
and U1020 (N_1020,N_843,N_823);
nand U1021 (N_1021,N_501,N_924);
or U1022 (N_1022,N_732,N_997);
and U1023 (N_1023,N_926,N_704);
and U1024 (N_1024,N_787,N_785);
or U1025 (N_1025,N_883,N_958);
nand U1026 (N_1026,In_708,N_790);
nand U1027 (N_1027,In_1166,N_245);
and U1028 (N_1028,N_796,N_824);
nand U1029 (N_1029,N_892,N_865);
nor U1030 (N_1030,N_729,N_461);
nor U1031 (N_1031,N_761,N_262);
nor U1032 (N_1032,N_866,N_601);
or U1033 (N_1033,N_957,N_822);
nor U1034 (N_1034,N_901,N_935);
and U1035 (N_1035,In_168,N_995);
and U1036 (N_1036,N_762,N_860);
nand U1037 (N_1037,N_97,N_943);
nor U1038 (N_1038,In_340,N_590);
or U1039 (N_1039,N_993,N_982);
or U1040 (N_1040,N_784,N_521);
nand U1041 (N_1041,In_795,N_942);
and U1042 (N_1042,N_950,In_702);
and U1043 (N_1043,N_583,N_864);
and U1044 (N_1044,In_205,N_967);
nand U1045 (N_1045,N_460,N_871);
and U1046 (N_1046,N_777,N_304);
nor U1047 (N_1047,N_953,N_800);
nor U1048 (N_1048,N_928,N_365);
or U1049 (N_1049,N_818,N_834);
nor U1050 (N_1050,N_812,N_988);
nand U1051 (N_1051,N_867,N_839);
nor U1052 (N_1052,N_611,N_794);
or U1053 (N_1053,In_758,N_757);
and U1054 (N_1054,N_841,In_1265);
and U1055 (N_1055,N_559,In_606);
or U1056 (N_1056,N_857,N_628);
and U1057 (N_1057,N_430,N_940);
nor U1058 (N_1058,N_992,N_846);
and U1059 (N_1059,N_587,In_741);
nor U1060 (N_1060,N_905,N_976);
or U1061 (N_1061,N_832,N_911);
or U1062 (N_1062,N_917,N_847);
and U1063 (N_1063,N_766,N_927);
and U1064 (N_1064,N_977,N_636);
nand U1065 (N_1065,N_939,In_239);
or U1066 (N_1066,N_776,N_614);
xor U1067 (N_1067,In_1482,N_659);
nor U1068 (N_1068,N_922,N_826);
or U1069 (N_1069,In_255,In_651);
nand U1070 (N_1070,N_817,N_585);
nor U1071 (N_1071,N_764,In_1402);
nor U1072 (N_1072,N_542,N_530);
or U1073 (N_1073,N_804,N_899);
or U1074 (N_1074,N_768,In_211);
xor U1075 (N_1075,In_1472,N_870);
or U1076 (N_1076,N_968,N_685);
or U1077 (N_1077,N_703,N_872);
or U1078 (N_1078,N_665,N_278);
nor U1079 (N_1079,N_844,N_835);
xnor U1080 (N_1080,N_214,In_1412);
or U1081 (N_1081,N_657,N_930);
and U1082 (N_1082,N_767,N_959);
and U1083 (N_1083,N_578,N_741);
nor U1084 (N_1084,N_309,N_756);
or U1085 (N_1085,N_885,N_808);
and U1086 (N_1086,N_773,N_123);
nand U1087 (N_1087,N_884,In_1212);
nor U1088 (N_1088,N_948,N_972);
or U1089 (N_1089,N_966,N_793);
or U1090 (N_1090,N_427,N_850);
or U1091 (N_1091,N_861,N_887);
and U1092 (N_1092,N_472,N_994);
and U1093 (N_1093,N_728,N_852);
or U1094 (N_1094,N_814,N_916);
nor U1095 (N_1095,In_1197,N_987);
nor U1096 (N_1096,N_999,N_531);
or U1097 (N_1097,N_900,N_400);
nor U1098 (N_1098,N_975,N_528);
nand U1099 (N_1099,N_684,N_313);
nand U1100 (N_1100,N_464,N_205);
or U1101 (N_1101,N_991,N_840);
or U1102 (N_1102,In_85,N_718);
nor U1103 (N_1103,In_577,N_910);
and U1104 (N_1104,N_271,N_407);
and U1105 (N_1105,In_575,In_445);
nor U1106 (N_1106,N_303,N_792);
nand U1107 (N_1107,In_388,N_547);
and U1108 (N_1108,In_398,In_634);
nand U1109 (N_1109,N_954,N_330);
nand U1110 (N_1110,N_783,In_541);
and U1111 (N_1111,In_512,N_813);
or U1112 (N_1112,N_556,N_778);
and U1113 (N_1113,N_797,N_538);
nand U1114 (N_1114,In_1396,N_828);
and U1115 (N_1115,N_709,N_669);
and U1116 (N_1116,N_825,N_921);
and U1117 (N_1117,N_481,N_710);
and U1118 (N_1118,N_786,N_909);
nand U1119 (N_1119,N_331,N_609);
nand U1120 (N_1120,N_848,N_424);
nor U1121 (N_1121,In_96,N_534);
or U1122 (N_1122,N_915,N_986);
nand U1123 (N_1123,N_934,In_148);
nor U1124 (N_1124,In_1271,N_908);
and U1125 (N_1125,N_862,N_970);
or U1126 (N_1126,N_964,N_962);
or U1127 (N_1127,N_886,N_54);
nor U1128 (N_1128,N_302,In_894);
nor U1129 (N_1129,In_1238,In_267);
or U1130 (N_1130,In_1008,N_739);
nand U1131 (N_1131,N_455,N_789);
or U1132 (N_1132,N_983,N_875);
or U1133 (N_1133,N_73,N_827);
and U1134 (N_1134,In_591,In_1386);
or U1135 (N_1135,N_597,In_1092);
and U1136 (N_1136,N_753,In_539);
and U1137 (N_1137,In_237,N_780);
nor U1138 (N_1138,N_838,N_156);
or U1139 (N_1139,In_1109,N_567);
nor U1140 (N_1140,N_912,In_721);
or U1141 (N_1141,N_980,N_589);
and U1142 (N_1142,In_287,N_856);
or U1143 (N_1143,In_726,N_863);
or U1144 (N_1144,In_531,N_605);
and U1145 (N_1145,In_735,N_744);
or U1146 (N_1146,In_406,In_1170);
and U1147 (N_1147,N_517,N_700);
nand U1148 (N_1148,In_1210,N_755);
and U1149 (N_1149,N_938,N_754);
nand U1150 (N_1150,N_405,N_961);
nand U1151 (N_1151,N_363,N_341);
or U1152 (N_1152,N_677,N_851);
xor U1153 (N_1153,N_420,N_791);
or U1154 (N_1154,N_606,N_443);
nand U1155 (N_1155,N_516,N_869);
and U1156 (N_1156,N_769,N_974);
or U1157 (N_1157,N_781,In_1183);
or U1158 (N_1158,N_963,N_971);
xnor U1159 (N_1159,In_1151,N_557);
and U1160 (N_1160,N_694,N_795);
and U1161 (N_1161,N_131,N_805);
and U1162 (N_1162,N_343,N_751);
nand U1163 (N_1163,N_837,In_1012);
nand U1164 (N_1164,N_830,N_770);
nand U1165 (N_1165,In_672,N_699);
and U1166 (N_1166,N_678,N_949);
and U1167 (N_1167,N_849,N_891);
nand U1168 (N_1168,N_779,N_815);
or U1169 (N_1169,In_743,N_811);
nor U1170 (N_1170,N_881,N_845);
nand U1171 (N_1171,N_577,N_888);
nor U1172 (N_1172,N_929,In_1481);
and U1173 (N_1173,In_1050,N_725);
nor U1174 (N_1174,N_882,N_524);
and U1175 (N_1175,N_502,N_616);
or U1176 (N_1176,N_858,In_40);
nand U1177 (N_1177,N_874,In_113);
and U1178 (N_1178,In_257,N_631);
or U1179 (N_1179,N_907,N_932);
nor U1180 (N_1180,In_1430,N_880);
or U1181 (N_1181,N_746,N_925);
or U1182 (N_1182,N_956,In_279);
xor U1183 (N_1183,N_760,N_680);
nand U1184 (N_1184,N_683,N_859);
or U1185 (N_1185,N_682,N_772);
or U1186 (N_1186,In_1384,N_520);
or U1187 (N_1187,N_955,In_580);
nand U1188 (N_1188,N_876,N_990);
nand U1189 (N_1189,In_813,N_829);
nor U1190 (N_1190,N_836,N_820);
or U1191 (N_1191,N_437,N_546);
and U1192 (N_1192,N_906,N_854);
nor U1193 (N_1193,N_763,N_635);
or U1194 (N_1194,In_600,N_889);
nor U1195 (N_1195,N_300,N_919);
nand U1196 (N_1196,N_613,In_534);
nor U1197 (N_1197,N_996,In_633);
nor U1198 (N_1198,N_952,N_931);
xor U1199 (N_1199,In_630,N_116);
or U1200 (N_1200,N_314,N_913);
and U1201 (N_1201,N_336,N_618);
nor U1202 (N_1202,N_960,In_242);
nand U1203 (N_1203,N_799,N_853);
nor U1204 (N_1204,N_946,N_873);
and U1205 (N_1205,In_126,In_207);
and U1206 (N_1206,In_638,N_855);
and U1207 (N_1207,N_510,In_954);
nand U1208 (N_1208,N_914,N_944);
or U1209 (N_1209,N_554,In_323);
and U1210 (N_1210,N_877,N_973);
nor U1211 (N_1211,N_806,N_291);
xor U1212 (N_1212,N_809,In_811);
nor U1213 (N_1213,N_788,N_902);
nand U1214 (N_1214,N_833,N_798);
or U1215 (N_1215,N_298,N_897);
nor U1216 (N_1216,N_758,N_383);
nor U1217 (N_1217,N_890,N_106);
nand U1218 (N_1218,N_674,In_1318);
and U1219 (N_1219,In_550,N_941);
and U1220 (N_1220,N_947,N_896);
or U1221 (N_1221,N_895,N_981);
or U1222 (N_1222,N_625,N_687);
or U1223 (N_1223,N_134,N_561);
and U1224 (N_1224,N_965,N_969);
or U1225 (N_1225,N_807,N_979);
nor U1226 (N_1226,N_373,N_752);
nor U1227 (N_1227,N_842,N_555);
nor U1228 (N_1228,N_879,N_978);
xor U1229 (N_1229,In_1437,N_128);
or U1230 (N_1230,N_731,N_706);
or U1231 (N_1231,N_989,N_750);
or U1232 (N_1232,N_951,N_571);
nor U1233 (N_1233,N_765,N_893);
nor U1234 (N_1234,N_898,N_923);
nor U1235 (N_1235,N_503,In_727);
nor U1236 (N_1236,N_250,N_679);
nand U1237 (N_1237,N_904,N_774);
nand U1238 (N_1238,In_235,In_1211);
and U1239 (N_1239,In_236,N_831);
nor U1240 (N_1240,N_816,N_918);
or U1241 (N_1241,N_548,N_759);
and U1242 (N_1242,N_292,In_226);
or U1243 (N_1243,N_819,N_984);
nand U1244 (N_1244,In_1419,N_803);
xnor U1245 (N_1245,N_937,N_27);
nand U1246 (N_1246,N_507,In_178);
nand U1247 (N_1247,N_936,In_1037);
or U1248 (N_1248,N_821,N_598);
and U1249 (N_1249,N_998,N_523);
xor U1250 (N_1250,N_1133,N_1006);
or U1251 (N_1251,N_1164,N_1249);
nor U1252 (N_1252,N_1203,N_1029);
nand U1253 (N_1253,N_1054,N_1047);
or U1254 (N_1254,N_1013,N_1210);
or U1255 (N_1255,N_1243,N_1145);
nand U1256 (N_1256,N_1128,N_1095);
nor U1257 (N_1257,N_1184,N_1126);
or U1258 (N_1258,N_1120,N_1223);
nor U1259 (N_1259,N_1053,N_1017);
or U1260 (N_1260,N_1228,N_1079);
and U1261 (N_1261,N_1211,N_1022);
or U1262 (N_1262,N_1192,N_1058);
nand U1263 (N_1263,N_1106,N_1207);
or U1264 (N_1264,N_1160,N_1169);
nor U1265 (N_1265,N_1062,N_1048);
or U1266 (N_1266,N_1246,N_1125);
nand U1267 (N_1267,N_1052,N_1086);
and U1268 (N_1268,N_1072,N_1123);
and U1269 (N_1269,N_1209,N_1194);
nor U1270 (N_1270,N_1204,N_1028);
xnor U1271 (N_1271,N_1186,N_1015);
and U1272 (N_1272,N_1027,N_1105);
xor U1273 (N_1273,N_1153,N_1036);
and U1274 (N_1274,N_1221,N_1127);
nand U1275 (N_1275,N_1011,N_1099);
nand U1276 (N_1276,N_1137,N_1044);
nor U1277 (N_1277,N_1213,N_1037);
or U1278 (N_1278,N_1232,N_1103);
and U1279 (N_1279,N_1091,N_1073);
xor U1280 (N_1280,N_1076,N_1132);
and U1281 (N_1281,N_1012,N_1090);
nand U1282 (N_1282,N_1189,N_1144);
nand U1283 (N_1283,N_1063,N_1065);
nor U1284 (N_1284,N_1059,N_1094);
or U1285 (N_1285,N_1046,N_1206);
nand U1286 (N_1286,N_1110,N_1051);
and U1287 (N_1287,N_1116,N_1122);
nor U1288 (N_1288,N_1101,N_1240);
and U1289 (N_1289,N_1118,N_1066);
and U1290 (N_1290,N_1085,N_1139);
or U1291 (N_1291,N_1010,N_1035);
nand U1292 (N_1292,N_1107,N_1092);
nor U1293 (N_1293,N_1142,N_1138);
or U1294 (N_1294,N_1061,N_1119);
nor U1295 (N_1295,N_1055,N_1177);
and U1296 (N_1296,N_1014,N_1057);
nand U1297 (N_1297,N_1007,N_1175);
nand U1298 (N_1298,N_1140,N_1056);
nand U1299 (N_1299,N_1236,N_1042);
nor U1300 (N_1300,N_1087,N_1187);
or U1301 (N_1301,N_1088,N_1024);
and U1302 (N_1302,N_1136,N_1161);
nand U1303 (N_1303,N_1016,N_1159);
nor U1304 (N_1304,N_1157,N_1067);
xor U1305 (N_1305,N_1039,N_1131);
nor U1306 (N_1306,N_1176,N_1166);
and U1307 (N_1307,N_1178,N_1075);
or U1308 (N_1308,N_1050,N_1069);
and U1309 (N_1309,N_1196,N_1023);
nand U1310 (N_1310,N_1233,N_1004);
or U1311 (N_1311,N_1245,N_1114);
nor U1312 (N_1312,N_1241,N_1020);
and U1313 (N_1313,N_1163,N_1235);
nor U1314 (N_1314,N_1038,N_1225);
or U1315 (N_1315,N_1064,N_1195);
or U1316 (N_1316,N_1185,N_1068);
nor U1317 (N_1317,N_1183,N_1190);
nand U1318 (N_1318,N_1170,N_1089);
or U1319 (N_1319,N_1108,N_1019);
nor U1320 (N_1320,N_1074,N_1081);
nor U1321 (N_1321,N_1165,N_1174);
nor U1322 (N_1322,N_1148,N_1151);
and U1323 (N_1323,N_1239,N_1030);
nor U1324 (N_1324,N_1231,N_1156);
and U1325 (N_1325,N_1003,N_1021);
nand U1326 (N_1326,N_1155,N_1043);
nand U1327 (N_1327,N_1134,N_1147);
or U1328 (N_1328,N_1179,N_1005);
nand U1329 (N_1329,N_1100,N_1129);
or U1330 (N_1330,N_1109,N_1244);
or U1331 (N_1331,N_1197,N_1049);
nand U1332 (N_1332,N_1070,N_1115);
nor U1333 (N_1333,N_1009,N_1117);
and U1334 (N_1334,N_1242,N_1083);
nor U1335 (N_1335,N_1078,N_1025);
nand U1336 (N_1336,N_1130,N_1198);
nand U1337 (N_1337,N_1172,N_1082);
or U1338 (N_1338,N_1121,N_1031);
nand U1339 (N_1339,N_1199,N_1216);
or U1340 (N_1340,N_1219,N_1224);
or U1341 (N_1341,N_1226,N_1201);
nor U1342 (N_1342,N_1162,N_1146);
nand U1343 (N_1343,N_1032,N_1098);
nand U1344 (N_1344,N_1045,N_1214);
and U1345 (N_1345,N_1248,N_1208);
nor U1346 (N_1346,N_1084,N_1182);
or U1347 (N_1347,N_1200,N_1222);
xnor U1348 (N_1348,N_1041,N_1077);
nor U1349 (N_1349,N_1071,N_1141);
nand U1350 (N_1350,N_1215,N_1002);
and U1351 (N_1351,N_1181,N_1113);
and U1352 (N_1352,N_1001,N_1173);
or U1353 (N_1353,N_1227,N_1237);
nor U1354 (N_1354,N_1111,N_1143);
nor U1355 (N_1355,N_1191,N_1188);
xnor U1356 (N_1356,N_1096,N_1008);
or U1357 (N_1357,N_1180,N_1168);
and U1358 (N_1358,N_1060,N_1104);
nand U1359 (N_1359,N_1124,N_1149);
nand U1360 (N_1360,N_1018,N_1220);
or U1361 (N_1361,N_1229,N_1152);
and U1362 (N_1362,N_1158,N_1230);
nand U1363 (N_1363,N_1218,N_1234);
nand U1364 (N_1364,N_1093,N_1171);
and U1365 (N_1365,N_1193,N_1212);
or U1366 (N_1366,N_1202,N_1080);
nand U1367 (N_1367,N_1167,N_1097);
nand U1368 (N_1368,N_1205,N_1217);
xor U1369 (N_1369,N_1135,N_1150);
and U1370 (N_1370,N_1033,N_1000);
or U1371 (N_1371,N_1238,N_1026);
nand U1372 (N_1372,N_1102,N_1154);
nand U1373 (N_1373,N_1112,N_1247);
or U1374 (N_1374,N_1034,N_1040);
nor U1375 (N_1375,N_1236,N_1048);
and U1376 (N_1376,N_1144,N_1194);
and U1377 (N_1377,N_1221,N_1132);
and U1378 (N_1378,N_1057,N_1003);
or U1379 (N_1379,N_1030,N_1042);
or U1380 (N_1380,N_1129,N_1041);
nand U1381 (N_1381,N_1191,N_1199);
or U1382 (N_1382,N_1009,N_1087);
nand U1383 (N_1383,N_1085,N_1191);
nor U1384 (N_1384,N_1112,N_1003);
nor U1385 (N_1385,N_1010,N_1129);
and U1386 (N_1386,N_1240,N_1182);
xor U1387 (N_1387,N_1037,N_1019);
or U1388 (N_1388,N_1020,N_1143);
nand U1389 (N_1389,N_1248,N_1069);
nand U1390 (N_1390,N_1206,N_1015);
nand U1391 (N_1391,N_1110,N_1187);
nor U1392 (N_1392,N_1023,N_1043);
and U1393 (N_1393,N_1117,N_1047);
nor U1394 (N_1394,N_1132,N_1170);
nor U1395 (N_1395,N_1113,N_1092);
nand U1396 (N_1396,N_1116,N_1113);
nor U1397 (N_1397,N_1187,N_1193);
nand U1398 (N_1398,N_1130,N_1165);
and U1399 (N_1399,N_1207,N_1192);
xor U1400 (N_1400,N_1243,N_1039);
and U1401 (N_1401,N_1206,N_1051);
nor U1402 (N_1402,N_1103,N_1215);
nor U1403 (N_1403,N_1024,N_1249);
nor U1404 (N_1404,N_1078,N_1057);
nand U1405 (N_1405,N_1192,N_1163);
nand U1406 (N_1406,N_1135,N_1115);
nor U1407 (N_1407,N_1197,N_1189);
xnor U1408 (N_1408,N_1001,N_1188);
or U1409 (N_1409,N_1011,N_1107);
nor U1410 (N_1410,N_1007,N_1104);
or U1411 (N_1411,N_1184,N_1188);
or U1412 (N_1412,N_1186,N_1161);
nand U1413 (N_1413,N_1021,N_1143);
and U1414 (N_1414,N_1084,N_1089);
or U1415 (N_1415,N_1179,N_1145);
and U1416 (N_1416,N_1124,N_1243);
nand U1417 (N_1417,N_1099,N_1075);
nor U1418 (N_1418,N_1119,N_1063);
nand U1419 (N_1419,N_1036,N_1033);
xnor U1420 (N_1420,N_1176,N_1071);
and U1421 (N_1421,N_1075,N_1221);
and U1422 (N_1422,N_1055,N_1240);
nor U1423 (N_1423,N_1049,N_1145);
or U1424 (N_1424,N_1091,N_1106);
or U1425 (N_1425,N_1238,N_1152);
nand U1426 (N_1426,N_1143,N_1060);
and U1427 (N_1427,N_1107,N_1032);
nand U1428 (N_1428,N_1007,N_1185);
or U1429 (N_1429,N_1004,N_1232);
nand U1430 (N_1430,N_1236,N_1115);
nand U1431 (N_1431,N_1207,N_1203);
and U1432 (N_1432,N_1033,N_1046);
or U1433 (N_1433,N_1230,N_1044);
nand U1434 (N_1434,N_1206,N_1078);
and U1435 (N_1435,N_1104,N_1005);
nand U1436 (N_1436,N_1107,N_1165);
or U1437 (N_1437,N_1093,N_1164);
or U1438 (N_1438,N_1121,N_1153);
and U1439 (N_1439,N_1062,N_1173);
or U1440 (N_1440,N_1146,N_1177);
nor U1441 (N_1441,N_1139,N_1241);
nand U1442 (N_1442,N_1085,N_1242);
nand U1443 (N_1443,N_1201,N_1061);
nor U1444 (N_1444,N_1222,N_1063);
and U1445 (N_1445,N_1242,N_1027);
nor U1446 (N_1446,N_1063,N_1138);
nor U1447 (N_1447,N_1171,N_1218);
and U1448 (N_1448,N_1050,N_1191);
nor U1449 (N_1449,N_1079,N_1033);
nand U1450 (N_1450,N_1113,N_1206);
or U1451 (N_1451,N_1035,N_1023);
or U1452 (N_1452,N_1082,N_1015);
and U1453 (N_1453,N_1086,N_1065);
or U1454 (N_1454,N_1228,N_1237);
nand U1455 (N_1455,N_1228,N_1017);
or U1456 (N_1456,N_1099,N_1130);
and U1457 (N_1457,N_1006,N_1072);
or U1458 (N_1458,N_1087,N_1196);
or U1459 (N_1459,N_1097,N_1208);
or U1460 (N_1460,N_1011,N_1094);
and U1461 (N_1461,N_1169,N_1032);
and U1462 (N_1462,N_1136,N_1206);
nor U1463 (N_1463,N_1013,N_1067);
and U1464 (N_1464,N_1223,N_1162);
or U1465 (N_1465,N_1017,N_1098);
nor U1466 (N_1466,N_1230,N_1017);
or U1467 (N_1467,N_1032,N_1060);
and U1468 (N_1468,N_1068,N_1140);
and U1469 (N_1469,N_1002,N_1247);
nand U1470 (N_1470,N_1164,N_1238);
or U1471 (N_1471,N_1149,N_1130);
or U1472 (N_1472,N_1246,N_1028);
nand U1473 (N_1473,N_1178,N_1024);
or U1474 (N_1474,N_1101,N_1224);
or U1475 (N_1475,N_1134,N_1162);
and U1476 (N_1476,N_1173,N_1046);
nor U1477 (N_1477,N_1158,N_1085);
nor U1478 (N_1478,N_1087,N_1142);
and U1479 (N_1479,N_1121,N_1003);
nand U1480 (N_1480,N_1225,N_1060);
nor U1481 (N_1481,N_1069,N_1174);
or U1482 (N_1482,N_1203,N_1204);
nor U1483 (N_1483,N_1069,N_1149);
nor U1484 (N_1484,N_1141,N_1049);
nor U1485 (N_1485,N_1174,N_1022);
nor U1486 (N_1486,N_1015,N_1160);
nor U1487 (N_1487,N_1183,N_1139);
and U1488 (N_1488,N_1222,N_1012);
and U1489 (N_1489,N_1207,N_1052);
and U1490 (N_1490,N_1078,N_1080);
and U1491 (N_1491,N_1057,N_1198);
or U1492 (N_1492,N_1106,N_1095);
and U1493 (N_1493,N_1030,N_1026);
or U1494 (N_1494,N_1091,N_1017);
nor U1495 (N_1495,N_1135,N_1001);
and U1496 (N_1496,N_1226,N_1053);
or U1497 (N_1497,N_1239,N_1106);
and U1498 (N_1498,N_1163,N_1109);
and U1499 (N_1499,N_1044,N_1016);
xor U1500 (N_1500,N_1305,N_1322);
nor U1501 (N_1501,N_1488,N_1255);
and U1502 (N_1502,N_1463,N_1476);
nor U1503 (N_1503,N_1407,N_1478);
nand U1504 (N_1504,N_1369,N_1465);
nand U1505 (N_1505,N_1473,N_1297);
or U1506 (N_1506,N_1251,N_1292);
nand U1507 (N_1507,N_1446,N_1336);
nor U1508 (N_1508,N_1385,N_1471);
and U1509 (N_1509,N_1360,N_1491);
nor U1510 (N_1510,N_1278,N_1472);
or U1511 (N_1511,N_1361,N_1301);
nand U1512 (N_1512,N_1450,N_1328);
or U1513 (N_1513,N_1283,N_1495);
nand U1514 (N_1514,N_1417,N_1290);
nand U1515 (N_1515,N_1431,N_1497);
and U1516 (N_1516,N_1314,N_1250);
nor U1517 (N_1517,N_1440,N_1368);
nand U1518 (N_1518,N_1358,N_1258);
and U1519 (N_1519,N_1400,N_1470);
nor U1520 (N_1520,N_1316,N_1345);
nor U1521 (N_1521,N_1344,N_1296);
or U1522 (N_1522,N_1371,N_1408);
or U1523 (N_1523,N_1461,N_1370);
nand U1524 (N_1524,N_1354,N_1259);
or U1525 (N_1525,N_1393,N_1428);
nand U1526 (N_1526,N_1264,N_1413);
nand U1527 (N_1527,N_1362,N_1294);
nor U1528 (N_1528,N_1373,N_1422);
nand U1529 (N_1529,N_1423,N_1492);
nor U1530 (N_1530,N_1256,N_1269);
nor U1531 (N_1531,N_1451,N_1280);
and U1532 (N_1532,N_1490,N_1330);
and U1533 (N_1533,N_1483,N_1341);
and U1534 (N_1534,N_1279,N_1432);
or U1535 (N_1535,N_1399,N_1268);
or U1536 (N_1536,N_1282,N_1350);
or U1537 (N_1537,N_1469,N_1386);
nand U1538 (N_1538,N_1460,N_1315);
nor U1539 (N_1539,N_1479,N_1310);
nand U1540 (N_1540,N_1397,N_1477);
nand U1541 (N_1541,N_1396,N_1437);
and U1542 (N_1542,N_1349,N_1254);
xnor U1543 (N_1543,N_1257,N_1430);
nor U1544 (N_1544,N_1334,N_1485);
nor U1545 (N_1545,N_1415,N_1475);
or U1546 (N_1546,N_1391,N_1337);
or U1547 (N_1547,N_1442,N_1348);
or U1548 (N_1548,N_1436,N_1416);
xnor U1549 (N_1549,N_1409,N_1274);
nor U1550 (N_1550,N_1335,N_1447);
nor U1551 (N_1551,N_1452,N_1494);
and U1552 (N_1552,N_1387,N_1339);
xor U1553 (N_1553,N_1406,N_1390);
nor U1554 (N_1554,N_1394,N_1424);
nor U1555 (N_1555,N_1306,N_1455);
or U1556 (N_1556,N_1457,N_1359);
or U1557 (N_1557,N_1281,N_1449);
nor U1558 (N_1558,N_1352,N_1453);
xnor U1559 (N_1559,N_1275,N_1454);
or U1560 (N_1560,N_1493,N_1321);
or U1561 (N_1561,N_1462,N_1323);
and U1562 (N_1562,N_1418,N_1356);
and U1563 (N_1563,N_1333,N_1403);
nor U1564 (N_1564,N_1398,N_1340);
nor U1565 (N_1565,N_1327,N_1487);
or U1566 (N_1566,N_1468,N_1380);
and U1567 (N_1567,N_1338,N_1474);
nor U1568 (N_1568,N_1342,N_1270);
and U1569 (N_1569,N_1482,N_1467);
xnor U1570 (N_1570,N_1298,N_1411);
nand U1571 (N_1571,N_1420,N_1299);
and U1572 (N_1572,N_1374,N_1262);
xor U1573 (N_1573,N_1367,N_1355);
nor U1574 (N_1574,N_1263,N_1311);
nor U1575 (N_1575,N_1496,N_1346);
or U1576 (N_1576,N_1443,N_1302);
and U1577 (N_1577,N_1324,N_1267);
or U1578 (N_1578,N_1375,N_1419);
nor U1579 (N_1579,N_1319,N_1410);
and U1580 (N_1580,N_1427,N_1372);
nand U1581 (N_1581,N_1308,N_1309);
and U1582 (N_1582,N_1404,N_1395);
nor U1583 (N_1583,N_1286,N_1276);
nand U1584 (N_1584,N_1277,N_1265);
nor U1585 (N_1585,N_1441,N_1381);
nand U1586 (N_1586,N_1405,N_1253);
nor U1587 (N_1587,N_1464,N_1384);
nand U1588 (N_1588,N_1312,N_1377);
and U1589 (N_1589,N_1351,N_1444);
nor U1590 (N_1590,N_1439,N_1285);
and U1591 (N_1591,N_1261,N_1456);
and U1592 (N_1592,N_1401,N_1343);
nand U1593 (N_1593,N_1466,N_1388);
and U1594 (N_1594,N_1325,N_1288);
or U1595 (N_1595,N_1284,N_1421);
nand U1596 (N_1596,N_1266,N_1320);
or U1597 (N_1597,N_1295,N_1433);
and U1598 (N_1598,N_1434,N_1379);
and U1599 (N_1599,N_1425,N_1389);
and U1600 (N_1600,N_1499,N_1318);
nand U1601 (N_1601,N_1382,N_1272);
nor U1602 (N_1602,N_1332,N_1353);
and U1603 (N_1603,N_1412,N_1392);
nor U1604 (N_1604,N_1287,N_1448);
or U1605 (N_1605,N_1289,N_1459);
and U1606 (N_1606,N_1307,N_1313);
nand U1607 (N_1607,N_1260,N_1291);
and U1608 (N_1608,N_1364,N_1363);
and U1609 (N_1609,N_1414,N_1366);
nand U1610 (N_1610,N_1438,N_1480);
nor U1611 (N_1611,N_1365,N_1429);
and U1612 (N_1612,N_1300,N_1331);
nor U1613 (N_1613,N_1317,N_1458);
nor U1614 (N_1614,N_1383,N_1293);
and U1615 (N_1615,N_1326,N_1252);
nor U1616 (N_1616,N_1376,N_1498);
or U1617 (N_1617,N_1273,N_1303);
and U1618 (N_1618,N_1445,N_1378);
and U1619 (N_1619,N_1484,N_1271);
nand U1620 (N_1620,N_1347,N_1481);
nand U1621 (N_1621,N_1426,N_1304);
nor U1622 (N_1622,N_1435,N_1357);
nand U1623 (N_1623,N_1329,N_1402);
and U1624 (N_1624,N_1486,N_1489);
xnor U1625 (N_1625,N_1315,N_1483);
or U1626 (N_1626,N_1395,N_1380);
or U1627 (N_1627,N_1412,N_1470);
or U1628 (N_1628,N_1378,N_1497);
and U1629 (N_1629,N_1400,N_1388);
and U1630 (N_1630,N_1285,N_1350);
and U1631 (N_1631,N_1338,N_1494);
or U1632 (N_1632,N_1380,N_1295);
and U1633 (N_1633,N_1458,N_1335);
and U1634 (N_1634,N_1274,N_1495);
or U1635 (N_1635,N_1458,N_1417);
and U1636 (N_1636,N_1274,N_1355);
and U1637 (N_1637,N_1373,N_1342);
or U1638 (N_1638,N_1271,N_1409);
nor U1639 (N_1639,N_1351,N_1280);
nand U1640 (N_1640,N_1270,N_1427);
nand U1641 (N_1641,N_1431,N_1477);
or U1642 (N_1642,N_1271,N_1278);
nor U1643 (N_1643,N_1313,N_1252);
and U1644 (N_1644,N_1327,N_1285);
nor U1645 (N_1645,N_1381,N_1254);
and U1646 (N_1646,N_1488,N_1468);
nand U1647 (N_1647,N_1342,N_1291);
or U1648 (N_1648,N_1328,N_1268);
or U1649 (N_1649,N_1451,N_1365);
or U1650 (N_1650,N_1278,N_1411);
and U1651 (N_1651,N_1390,N_1264);
and U1652 (N_1652,N_1447,N_1495);
or U1653 (N_1653,N_1432,N_1337);
nor U1654 (N_1654,N_1331,N_1409);
nand U1655 (N_1655,N_1341,N_1425);
or U1656 (N_1656,N_1466,N_1495);
or U1657 (N_1657,N_1342,N_1262);
nand U1658 (N_1658,N_1397,N_1357);
or U1659 (N_1659,N_1280,N_1399);
nand U1660 (N_1660,N_1296,N_1425);
or U1661 (N_1661,N_1485,N_1474);
xnor U1662 (N_1662,N_1276,N_1253);
nor U1663 (N_1663,N_1383,N_1310);
and U1664 (N_1664,N_1429,N_1496);
and U1665 (N_1665,N_1304,N_1380);
nand U1666 (N_1666,N_1346,N_1407);
or U1667 (N_1667,N_1414,N_1427);
nand U1668 (N_1668,N_1300,N_1405);
nor U1669 (N_1669,N_1371,N_1423);
and U1670 (N_1670,N_1499,N_1384);
nand U1671 (N_1671,N_1257,N_1266);
or U1672 (N_1672,N_1343,N_1416);
nand U1673 (N_1673,N_1265,N_1418);
or U1674 (N_1674,N_1324,N_1387);
xor U1675 (N_1675,N_1495,N_1430);
xnor U1676 (N_1676,N_1339,N_1439);
nand U1677 (N_1677,N_1385,N_1428);
and U1678 (N_1678,N_1394,N_1386);
and U1679 (N_1679,N_1424,N_1270);
and U1680 (N_1680,N_1438,N_1277);
nand U1681 (N_1681,N_1387,N_1315);
nor U1682 (N_1682,N_1251,N_1405);
nand U1683 (N_1683,N_1370,N_1426);
nor U1684 (N_1684,N_1372,N_1392);
nand U1685 (N_1685,N_1368,N_1282);
nand U1686 (N_1686,N_1282,N_1340);
or U1687 (N_1687,N_1350,N_1430);
or U1688 (N_1688,N_1423,N_1256);
and U1689 (N_1689,N_1407,N_1460);
nor U1690 (N_1690,N_1426,N_1450);
and U1691 (N_1691,N_1472,N_1357);
or U1692 (N_1692,N_1315,N_1486);
and U1693 (N_1693,N_1275,N_1337);
nand U1694 (N_1694,N_1443,N_1396);
nor U1695 (N_1695,N_1457,N_1251);
or U1696 (N_1696,N_1297,N_1497);
xor U1697 (N_1697,N_1399,N_1362);
and U1698 (N_1698,N_1299,N_1298);
xor U1699 (N_1699,N_1494,N_1321);
or U1700 (N_1700,N_1280,N_1482);
nand U1701 (N_1701,N_1301,N_1434);
or U1702 (N_1702,N_1477,N_1486);
and U1703 (N_1703,N_1451,N_1488);
and U1704 (N_1704,N_1354,N_1451);
nand U1705 (N_1705,N_1336,N_1395);
nand U1706 (N_1706,N_1483,N_1406);
nor U1707 (N_1707,N_1379,N_1403);
nor U1708 (N_1708,N_1477,N_1415);
nor U1709 (N_1709,N_1451,N_1419);
and U1710 (N_1710,N_1387,N_1486);
and U1711 (N_1711,N_1408,N_1271);
xor U1712 (N_1712,N_1354,N_1427);
nor U1713 (N_1713,N_1346,N_1348);
nand U1714 (N_1714,N_1250,N_1270);
nand U1715 (N_1715,N_1491,N_1298);
and U1716 (N_1716,N_1266,N_1391);
or U1717 (N_1717,N_1419,N_1425);
and U1718 (N_1718,N_1352,N_1306);
or U1719 (N_1719,N_1467,N_1485);
nand U1720 (N_1720,N_1332,N_1440);
nor U1721 (N_1721,N_1391,N_1273);
xor U1722 (N_1722,N_1344,N_1474);
and U1723 (N_1723,N_1463,N_1374);
nor U1724 (N_1724,N_1388,N_1309);
and U1725 (N_1725,N_1300,N_1272);
xnor U1726 (N_1726,N_1354,N_1275);
xor U1727 (N_1727,N_1479,N_1262);
nor U1728 (N_1728,N_1441,N_1264);
or U1729 (N_1729,N_1364,N_1476);
nor U1730 (N_1730,N_1257,N_1420);
and U1731 (N_1731,N_1298,N_1489);
nor U1732 (N_1732,N_1370,N_1322);
nor U1733 (N_1733,N_1471,N_1355);
or U1734 (N_1734,N_1483,N_1357);
nand U1735 (N_1735,N_1344,N_1445);
and U1736 (N_1736,N_1360,N_1412);
and U1737 (N_1737,N_1352,N_1455);
and U1738 (N_1738,N_1461,N_1494);
and U1739 (N_1739,N_1333,N_1348);
nand U1740 (N_1740,N_1457,N_1298);
or U1741 (N_1741,N_1376,N_1258);
nand U1742 (N_1742,N_1372,N_1354);
and U1743 (N_1743,N_1443,N_1421);
nand U1744 (N_1744,N_1345,N_1462);
xnor U1745 (N_1745,N_1368,N_1353);
nand U1746 (N_1746,N_1372,N_1483);
nand U1747 (N_1747,N_1381,N_1486);
nand U1748 (N_1748,N_1395,N_1481);
nand U1749 (N_1749,N_1427,N_1379);
nor U1750 (N_1750,N_1592,N_1718);
and U1751 (N_1751,N_1649,N_1500);
nor U1752 (N_1752,N_1615,N_1535);
or U1753 (N_1753,N_1508,N_1548);
nor U1754 (N_1754,N_1536,N_1523);
or U1755 (N_1755,N_1555,N_1520);
and U1756 (N_1756,N_1614,N_1564);
nand U1757 (N_1757,N_1580,N_1665);
nand U1758 (N_1758,N_1747,N_1725);
nor U1759 (N_1759,N_1590,N_1559);
nor U1760 (N_1760,N_1558,N_1654);
or U1761 (N_1761,N_1687,N_1708);
nor U1762 (N_1762,N_1639,N_1678);
nand U1763 (N_1763,N_1749,N_1566);
nand U1764 (N_1764,N_1578,N_1632);
nor U1765 (N_1765,N_1547,N_1728);
nand U1766 (N_1766,N_1634,N_1664);
nand U1767 (N_1767,N_1703,N_1528);
and U1768 (N_1768,N_1530,N_1674);
and U1769 (N_1769,N_1618,N_1586);
nor U1770 (N_1770,N_1745,N_1638);
or U1771 (N_1771,N_1669,N_1613);
nand U1772 (N_1772,N_1581,N_1648);
or U1773 (N_1773,N_1720,N_1546);
nand U1774 (N_1774,N_1666,N_1604);
nand U1775 (N_1775,N_1606,N_1731);
or U1776 (N_1776,N_1732,N_1624);
nor U1777 (N_1777,N_1589,N_1599);
or U1778 (N_1778,N_1647,N_1710);
or U1779 (N_1779,N_1585,N_1743);
nand U1780 (N_1780,N_1537,N_1739);
nand U1781 (N_1781,N_1712,N_1680);
nand U1782 (N_1782,N_1736,N_1602);
nor U1783 (N_1783,N_1574,N_1646);
or U1784 (N_1784,N_1593,N_1697);
nor U1785 (N_1785,N_1700,N_1543);
nand U1786 (N_1786,N_1587,N_1716);
nand U1787 (N_1787,N_1635,N_1699);
or U1788 (N_1788,N_1529,N_1588);
nand U1789 (N_1789,N_1692,N_1730);
and U1790 (N_1790,N_1741,N_1531);
and U1791 (N_1791,N_1533,N_1696);
nor U1792 (N_1792,N_1518,N_1641);
or U1793 (N_1793,N_1659,N_1506);
and U1794 (N_1794,N_1622,N_1617);
or U1795 (N_1795,N_1527,N_1633);
nor U1796 (N_1796,N_1663,N_1693);
nand U1797 (N_1797,N_1541,N_1724);
or U1798 (N_1798,N_1517,N_1538);
or U1799 (N_1799,N_1683,N_1675);
or U1800 (N_1800,N_1723,N_1607);
nand U1801 (N_1801,N_1553,N_1577);
nor U1802 (N_1802,N_1576,N_1542);
and U1803 (N_1803,N_1704,N_1667);
and U1804 (N_1804,N_1544,N_1691);
or U1805 (N_1805,N_1706,N_1561);
nor U1806 (N_1806,N_1713,N_1524);
and U1807 (N_1807,N_1673,N_1568);
or U1808 (N_1808,N_1655,N_1511);
nand U1809 (N_1809,N_1603,N_1637);
nor U1810 (N_1810,N_1557,N_1554);
and U1811 (N_1811,N_1540,N_1643);
nor U1812 (N_1812,N_1682,N_1620);
nor U1813 (N_1813,N_1522,N_1549);
and U1814 (N_1814,N_1545,N_1668);
nand U1815 (N_1815,N_1616,N_1626);
or U1816 (N_1816,N_1630,N_1662);
or U1817 (N_1817,N_1658,N_1726);
or U1818 (N_1818,N_1645,N_1686);
and U1819 (N_1819,N_1514,N_1597);
or U1820 (N_1820,N_1516,N_1627);
or U1821 (N_1821,N_1619,N_1707);
and U1822 (N_1822,N_1521,N_1661);
and U1823 (N_1823,N_1660,N_1711);
and U1824 (N_1824,N_1701,N_1734);
and U1825 (N_1825,N_1628,N_1600);
and U1826 (N_1826,N_1575,N_1556);
nor U1827 (N_1827,N_1709,N_1740);
and U1828 (N_1828,N_1512,N_1735);
and U1829 (N_1829,N_1583,N_1567);
and U1830 (N_1830,N_1525,N_1507);
nor U1831 (N_1831,N_1656,N_1601);
nand U1832 (N_1832,N_1653,N_1676);
nand U1833 (N_1833,N_1717,N_1563);
and U1834 (N_1834,N_1591,N_1515);
nor U1835 (N_1835,N_1502,N_1519);
nor U1836 (N_1836,N_1623,N_1594);
or U1837 (N_1837,N_1650,N_1672);
nand U1838 (N_1838,N_1612,N_1631);
nor U1839 (N_1839,N_1610,N_1738);
nor U1840 (N_1840,N_1510,N_1582);
or U1841 (N_1841,N_1539,N_1677);
and U1842 (N_1842,N_1690,N_1695);
and U1843 (N_1843,N_1727,N_1551);
and U1844 (N_1844,N_1565,N_1694);
and U1845 (N_1845,N_1670,N_1552);
nor U1846 (N_1846,N_1596,N_1671);
and U1847 (N_1847,N_1513,N_1526);
or U1848 (N_1848,N_1609,N_1642);
or U1849 (N_1849,N_1729,N_1579);
nor U1850 (N_1850,N_1742,N_1685);
nand U1851 (N_1851,N_1573,N_1550);
and U1852 (N_1852,N_1688,N_1560);
and U1853 (N_1853,N_1621,N_1651);
and U1854 (N_1854,N_1721,N_1595);
and U1855 (N_1855,N_1503,N_1744);
nand U1856 (N_1856,N_1504,N_1652);
nand U1857 (N_1857,N_1702,N_1657);
xor U1858 (N_1858,N_1501,N_1698);
or U1859 (N_1859,N_1640,N_1733);
nand U1860 (N_1860,N_1722,N_1681);
and U1861 (N_1861,N_1584,N_1636);
and U1862 (N_1862,N_1509,N_1746);
nor U1863 (N_1863,N_1598,N_1737);
or U1864 (N_1864,N_1570,N_1715);
or U1865 (N_1865,N_1629,N_1505);
nor U1866 (N_1866,N_1611,N_1532);
and U1867 (N_1867,N_1608,N_1572);
or U1868 (N_1868,N_1705,N_1689);
and U1869 (N_1869,N_1534,N_1569);
nand U1870 (N_1870,N_1571,N_1684);
and U1871 (N_1871,N_1605,N_1625);
xnor U1872 (N_1872,N_1719,N_1679);
nor U1873 (N_1873,N_1562,N_1644);
and U1874 (N_1874,N_1714,N_1748);
nor U1875 (N_1875,N_1520,N_1661);
nor U1876 (N_1876,N_1622,N_1573);
and U1877 (N_1877,N_1614,N_1512);
nor U1878 (N_1878,N_1526,N_1742);
and U1879 (N_1879,N_1606,N_1738);
and U1880 (N_1880,N_1706,N_1727);
or U1881 (N_1881,N_1592,N_1606);
nor U1882 (N_1882,N_1693,N_1646);
or U1883 (N_1883,N_1691,N_1685);
and U1884 (N_1884,N_1598,N_1655);
or U1885 (N_1885,N_1503,N_1528);
or U1886 (N_1886,N_1630,N_1650);
nand U1887 (N_1887,N_1607,N_1680);
nand U1888 (N_1888,N_1501,N_1692);
and U1889 (N_1889,N_1590,N_1538);
nor U1890 (N_1890,N_1620,N_1630);
or U1891 (N_1891,N_1577,N_1588);
nand U1892 (N_1892,N_1652,N_1522);
nor U1893 (N_1893,N_1728,N_1658);
and U1894 (N_1894,N_1741,N_1519);
or U1895 (N_1895,N_1545,N_1698);
nand U1896 (N_1896,N_1528,N_1588);
nand U1897 (N_1897,N_1680,N_1614);
nand U1898 (N_1898,N_1527,N_1679);
nor U1899 (N_1899,N_1540,N_1617);
nor U1900 (N_1900,N_1527,N_1661);
nand U1901 (N_1901,N_1628,N_1549);
or U1902 (N_1902,N_1734,N_1585);
or U1903 (N_1903,N_1634,N_1621);
or U1904 (N_1904,N_1744,N_1701);
nand U1905 (N_1905,N_1704,N_1523);
or U1906 (N_1906,N_1514,N_1505);
nor U1907 (N_1907,N_1676,N_1514);
or U1908 (N_1908,N_1664,N_1650);
or U1909 (N_1909,N_1615,N_1555);
nor U1910 (N_1910,N_1525,N_1565);
and U1911 (N_1911,N_1588,N_1617);
nand U1912 (N_1912,N_1590,N_1655);
and U1913 (N_1913,N_1598,N_1615);
or U1914 (N_1914,N_1615,N_1668);
and U1915 (N_1915,N_1699,N_1628);
and U1916 (N_1916,N_1508,N_1515);
and U1917 (N_1917,N_1619,N_1602);
or U1918 (N_1918,N_1504,N_1606);
and U1919 (N_1919,N_1667,N_1749);
nor U1920 (N_1920,N_1550,N_1697);
nand U1921 (N_1921,N_1620,N_1529);
or U1922 (N_1922,N_1636,N_1604);
or U1923 (N_1923,N_1680,N_1644);
and U1924 (N_1924,N_1694,N_1686);
xor U1925 (N_1925,N_1558,N_1609);
and U1926 (N_1926,N_1645,N_1610);
nor U1927 (N_1927,N_1630,N_1562);
nor U1928 (N_1928,N_1596,N_1609);
xor U1929 (N_1929,N_1664,N_1573);
and U1930 (N_1930,N_1536,N_1510);
and U1931 (N_1931,N_1583,N_1738);
nand U1932 (N_1932,N_1628,N_1631);
nand U1933 (N_1933,N_1723,N_1572);
nand U1934 (N_1934,N_1523,N_1539);
nand U1935 (N_1935,N_1535,N_1587);
or U1936 (N_1936,N_1647,N_1676);
xnor U1937 (N_1937,N_1618,N_1583);
or U1938 (N_1938,N_1548,N_1624);
and U1939 (N_1939,N_1701,N_1584);
and U1940 (N_1940,N_1669,N_1527);
and U1941 (N_1941,N_1509,N_1532);
or U1942 (N_1942,N_1682,N_1520);
xor U1943 (N_1943,N_1548,N_1635);
and U1944 (N_1944,N_1590,N_1580);
nor U1945 (N_1945,N_1585,N_1537);
nor U1946 (N_1946,N_1561,N_1652);
nor U1947 (N_1947,N_1570,N_1564);
and U1948 (N_1948,N_1630,N_1505);
nand U1949 (N_1949,N_1527,N_1707);
or U1950 (N_1950,N_1574,N_1719);
and U1951 (N_1951,N_1668,N_1522);
and U1952 (N_1952,N_1594,N_1652);
nor U1953 (N_1953,N_1516,N_1623);
nand U1954 (N_1954,N_1681,N_1525);
or U1955 (N_1955,N_1509,N_1637);
nand U1956 (N_1956,N_1533,N_1520);
nor U1957 (N_1957,N_1671,N_1537);
or U1958 (N_1958,N_1645,N_1512);
or U1959 (N_1959,N_1743,N_1725);
and U1960 (N_1960,N_1528,N_1689);
nor U1961 (N_1961,N_1679,N_1542);
and U1962 (N_1962,N_1696,N_1534);
nor U1963 (N_1963,N_1626,N_1545);
and U1964 (N_1964,N_1609,N_1556);
nand U1965 (N_1965,N_1500,N_1593);
and U1966 (N_1966,N_1634,N_1527);
nand U1967 (N_1967,N_1517,N_1737);
or U1968 (N_1968,N_1646,N_1501);
and U1969 (N_1969,N_1550,N_1728);
nand U1970 (N_1970,N_1636,N_1576);
or U1971 (N_1971,N_1642,N_1619);
nand U1972 (N_1972,N_1597,N_1692);
and U1973 (N_1973,N_1562,N_1586);
and U1974 (N_1974,N_1624,N_1672);
nand U1975 (N_1975,N_1562,N_1642);
or U1976 (N_1976,N_1558,N_1542);
nor U1977 (N_1977,N_1685,N_1718);
nor U1978 (N_1978,N_1725,N_1712);
nor U1979 (N_1979,N_1519,N_1511);
or U1980 (N_1980,N_1670,N_1534);
nor U1981 (N_1981,N_1715,N_1507);
or U1982 (N_1982,N_1617,N_1740);
and U1983 (N_1983,N_1695,N_1737);
nor U1984 (N_1984,N_1722,N_1676);
and U1985 (N_1985,N_1634,N_1529);
and U1986 (N_1986,N_1560,N_1541);
or U1987 (N_1987,N_1695,N_1557);
and U1988 (N_1988,N_1657,N_1560);
nor U1989 (N_1989,N_1534,N_1515);
nand U1990 (N_1990,N_1555,N_1718);
or U1991 (N_1991,N_1681,N_1644);
xor U1992 (N_1992,N_1609,N_1693);
nand U1993 (N_1993,N_1695,N_1697);
nor U1994 (N_1994,N_1583,N_1745);
nand U1995 (N_1995,N_1691,N_1639);
nand U1996 (N_1996,N_1667,N_1583);
and U1997 (N_1997,N_1586,N_1593);
nand U1998 (N_1998,N_1506,N_1741);
nor U1999 (N_1999,N_1748,N_1552);
and U2000 (N_2000,N_1930,N_1903);
nor U2001 (N_2001,N_1957,N_1976);
or U2002 (N_2002,N_1829,N_1991);
nand U2003 (N_2003,N_1937,N_1926);
nor U2004 (N_2004,N_1972,N_1792);
and U2005 (N_2005,N_1954,N_1776);
and U2006 (N_2006,N_1783,N_1808);
nor U2007 (N_2007,N_1925,N_1941);
and U2008 (N_2008,N_1968,N_1813);
nor U2009 (N_2009,N_1870,N_1880);
or U2010 (N_2010,N_1781,N_1987);
or U2011 (N_2011,N_1990,N_1777);
or U2012 (N_2012,N_1786,N_1833);
nand U2013 (N_2013,N_1796,N_1890);
nand U2014 (N_2014,N_1966,N_1970);
and U2015 (N_2015,N_1846,N_1791);
nor U2016 (N_2016,N_1995,N_1801);
and U2017 (N_2017,N_1921,N_1996);
nor U2018 (N_2018,N_1894,N_1751);
nand U2019 (N_2019,N_1812,N_1784);
nand U2020 (N_2020,N_1797,N_1815);
or U2021 (N_2021,N_1851,N_1849);
or U2022 (N_2022,N_1963,N_1943);
and U2023 (N_2023,N_1762,N_1764);
nor U2024 (N_2024,N_1800,N_1848);
or U2025 (N_2025,N_1779,N_1872);
nand U2026 (N_2026,N_1765,N_1753);
nand U2027 (N_2027,N_1977,N_1854);
or U2028 (N_2028,N_1861,N_1757);
or U2029 (N_2029,N_1940,N_1806);
and U2030 (N_2030,N_1986,N_1874);
and U2031 (N_2031,N_1973,N_1799);
nand U2032 (N_2032,N_1975,N_1928);
nand U2033 (N_2033,N_1760,N_1898);
nor U2034 (N_2034,N_1924,N_1844);
or U2035 (N_2035,N_1879,N_1752);
nand U2036 (N_2036,N_1809,N_1814);
nand U2037 (N_2037,N_1978,N_1923);
or U2038 (N_2038,N_1980,N_1778);
and U2039 (N_2039,N_1878,N_1931);
or U2040 (N_2040,N_1821,N_1811);
nor U2041 (N_2041,N_1913,N_1858);
or U2042 (N_2042,N_1947,N_1877);
or U2043 (N_2043,N_1969,N_1911);
or U2044 (N_2044,N_1759,N_1998);
or U2045 (N_2045,N_1948,N_1847);
or U2046 (N_2046,N_1934,N_1962);
or U2047 (N_2047,N_1876,N_1852);
or U2048 (N_2048,N_1901,N_1896);
or U2049 (N_2049,N_1845,N_1782);
or U2050 (N_2050,N_1841,N_1804);
or U2051 (N_2051,N_1895,N_1971);
nor U2052 (N_2052,N_1956,N_1768);
and U2053 (N_2053,N_1824,N_1802);
nor U2054 (N_2054,N_1899,N_1827);
and U2055 (N_2055,N_1953,N_1793);
nand U2056 (N_2056,N_1774,N_1859);
and U2057 (N_2057,N_1974,N_1922);
nand U2058 (N_2058,N_1885,N_1871);
or U2059 (N_2059,N_1912,N_1839);
and U2060 (N_2060,N_1864,N_1881);
or U2061 (N_2061,N_1888,N_1788);
nand U2062 (N_2062,N_1886,N_1989);
or U2063 (N_2063,N_1767,N_1887);
nand U2064 (N_2064,N_1843,N_1761);
nor U2065 (N_2065,N_1900,N_1798);
nor U2066 (N_2066,N_1984,N_1772);
and U2067 (N_2067,N_1866,N_1840);
nor U2068 (N_2068,N_1983,N_1826);
and U2069 (N_2069,N_1938,N_1959);
nor U2070 (N_2070,N_1834,N_1936);
or U2071 (N_2071,N_1999,N_1914);
or U2072 (N_2072,N_1863,N_1891);
or U2073 (N_2073,N_1915,N_1951);
and U2074 (N_2074,N_1836,N_1960);
xnor U2075 (N_2075,N_1822,N_1916);
xnor U2076 (N_2076,N_1917,N_1869);
and U2077 (N_2077,N_1771,N_1985);
xor U2078 (N_2078,N_1944,N_1856);
or U2079 (N_2079,N_1997,N_1750);
nand U2080 (N_2080,N_1906,N_1904);
nand U2081 (N_2081,N_1754,N_1819);
nand U2082 (N_2082,N_1927,N_1865);
nor U2083 (N_2083,N_1908,N_1942);
nor U2084 (N_2084,N_1875,N_1860);
nand U2085 (N_2085,N_1823,N_1838);
and U2086 (N_2086,N_1805,N_1992);
nand U2087 (N_2087,N_1807,N_1817);
and U2088 (N_2088,N_1905,N_1945);
nor U2089 (N_2089,N_1850,N_1889);
or U2090 (N_2090,N_1785,N_1892);
or U2091 (N_2091,N_1935,N_1979);
or U2092 (N_2092,N_1756,N_1883);
and U2093 (N_2093,N_1918,N_1775);
nor U2094 (N_2094,N_1902,N_1820);
nand U2095 (N_2095,N_1946,N_1909);
nand U2096 (N_2096,N_1939,N_1949);
and U2097 (N_2097,N_1955,N_1929);
or U2098 (N_2098,N_1831,N_1832);
or U2099 (N_2099,N_1950,N_1964);
and U2100 (N_2100,N_1868,N_1994);
nor U2101 (N_2101,N_1780,N_1867);
and U2102 (N_2102,N_1988,N_1897);
or U2103 (N_2103,N_1816,N_1755);
or U2104 (N_2104,N_1795,N_1794);
or U2105 (N_2105,N_1773,N_1758);
or U2106 (N_2106,N_1769,N_1853);
nor U2107 (N_2107,N_1803,N_1857);
nor U2108 (N_2108,N_1958,N_1952);
nor U2109 (N_2109,N_1789,N_1933);
or U2110 (N_2110,N_1862,N_1810);
and U2111 (N_2111,N_1910,N_1818);
nand U2112 (N_2112,N_1884,N_1965);
nor U2113 (N_2113,N_1835,N_1981);
and U2114 (N_2114,N_1920,N_1993);
and U2115 (N_2115,N_1770,N_1961);
and U2116 (N_2116,N_1766,N_1873);
or U2117 (N_2117,N_1830,N_1882);
nand U2118 (N_2118,N_1967,N_1787);
nand U2119 (N_2119,N_1837,N_1893);
and U2120 (N_2120,N_1907,N_1932);
nand U2121 (N_2121,N_1982,N_1842);
or U2122 (N_2122,N_1790,N_1763);
nor U2123 (N_2123,N_1919,N_1855);
nand U2124 (N_2124,N_1825,N_1828);
and U2125 (N_2125,N_1805,N_1911);
nand U2126 (N_2126,N_1969,N_1795);
nand U2127 (N_2127,N_1856,N_1994);
nor U2128 (N_2128,N_1834,N_1796);
or U2129 (N_2129,N_1977,N_1919);
and U2130 (N_2130,N_1906,N_1899);
or U2131 (N_2131,N_1952,N_1804);
nor U2132 (N_2132,N_1788,N_1970);
nor U2133 (N_2133,N_1986,N_1879);
nand U2134 (N_2134,N_1830,N_1961);
and U2135 (N_2135,N_1962,N_1869);
or U2136 (N_2136,N_1985,N_1821);
or U2137 (N_2137,N_1940,N_1944);
nor U2138 (N_2138,N_1906,N_1897);
or U2139 (N_2139,N_1829,N_1864);
nor U2140 (N_2140,N_1815,N_1874);
or U2141 (N_2141,N_1911,N_1850);
nor U2142 (N_2142,N_1897,N_1892);
or U2143 (N_2143,N_1985,N_1818);
and U2144 (N_2144,N_1968,N_1788);
or U2145 (N_2145,N_1910,N_1782);
or U2146 (N_2146,N_1985,N_1974);
and U2147 (N_2147,N_1835,N_1964);
and U2148 (N_2148,N_1839,N_1936);
nand U2149 (N_2149,N_1780,N_1930);
nand U2150 (N_2150,N_1812,N_1852);
and U2151 (N_2151,N_1881,N_1833);
and U2152 (N_2152,N_1837,N_1804);
nand U2153 (N_2153,N_1908,N_1986);
and U2154 (N_2154,N_1928,N_1923);
nand U2155 (N_2155,N_1870,N_1764);
and U2156 (N_2156,N_1796,N_1947);
and U2157 (N_2157,N_1803,N_1766);
xnor U2158 (N_2158,N_1764,N_1950);
nand U2159 (N_2159,N_1853,N_1860);
nor U2160 (N_2160,N_1885,N_1880);
nand U2161 (N_2161,N_1806,N_1920);
nand U2162 (N_2162,N_1754,N_1825);
nor U2163 (N_2163,N_1823,N_1869);
nand U2164 (N_2164,N_1982,N_1788);
nor U2165 (N_2165,N_1885,N_1773);
nor U2166 (N_2166,N_1875,N_1994);
nor U2167 (N_2167,N_1795,N_1934);
or U2168 (N_2168,N_1866,N_1812);
and U2169 (N_2169,N_1757,N_1750);
nand U2170 (N_2170,N_1874,N_1991);
nand U2171 (N_2171,N_1822,N_1961);
and U2172 (N_2172,N_1790,N_1768);
or U2173 (N_2173,N_1859,N_1908);
nand U2174 (N_2174,N_1848,N_1798);
nand U2175 (N_2175,N_1976,N_1779);
nor U2176 (N_2176,N_1816,N_1785);
and U2177 (N_2177,N_1937,N_1921);
xor U2178 (N_2178,N_1951,N_1914);
nand U2179 (N_2179,N_1924,N_1760);
and U2180 (N_2180,N_1959,N_1961);
or U2181 (N_2181,N_1937,N_1933);
nor U2182 (N_2182,N_1765,N_1876);
or U2183 (N_2183,N_1859,N_1840);
nand U2184 (N_2184,N_1820,N_1861);
nor U2185 (N_2185,N_1782,N_1789);
nand U2186 (N_2186,N_1862,N_1837);
nor U2187 (N_2187,N_1867,N_1797);
nor U2188 (N_2188,N_1812,N_1854);
and U2189 (N_2189,N_1932,N_1834);
and U2190 (N_2190,N_1805,N_1813);
or U2191 (N_2191,N_1829,N_1948);
nor U2192 (N_2192,N_1949,N_1851);
nor U2193 (N_2193,N_1851,N_1906);
nor U2194 (N_2194,N_1953,N_1856);
nor U2195 (N_2195,N_1870,N_1922);
nor U2196 (N_2196,N_1855,N_1971);
nor U2197 (N_2197,N_1880,N_1757);
xor U2198 (N_2198,N_1832,N_1791);
nand U2199 (N_2199,N_1842,N_1985);
nand U2200 (N_2200,N_1928,N_1872);
nor U2201 (N_2201,N_1815,N_1937);
nor U2202 (N_2202,N_1908,N_1934);
nor U2203 (N_2203,N_1801,N_1796);
or U2204 (N_2204,N_1764,N_1977);
and U2205 (N_2205,N_1818,N_1988);
nor U2206 (N_2206,N_1794,N_1770);
and U2207 (N_2207,N_1948,N_1767);
nor U2208 (N_2208,N_1761,N_1990);
and U2209 (N_2209,N_1790,N_1793);
nor U2210 (N_2210,N_1828,N_1785);
nor U2211 (N_2211,N_1766,N_1775);
or U2212 (N_2212,N_1831,N_1794);
and U2213 (N_2213,N_1758,N_1991);
and U2214 (N_2214,N_1772,N_1768);
or U2215 (N_2215,N_1783,N_1997);
and U2216 (N_2216,N_1842,N_1756);
or U2217 (N_2217,N_1780,N_1852);
nand U2218 (N_2218,N_1790,N_1780);
nor U2219 (N_2219,N_1824,N_1969);
nand U2220 (N_2220,N_1885,N_1941);
nand U2221 (N_2221,N_1839,N_1948);
and U2222 (N_2222,N_1974,N_1849);
or U2223 (N_2223,N_1874,N_1916);
nor U2224 (N_2224,N_1894,N_1826);
nor U2225 (N_2225,N_1818,N_1959);
and U2226 (N_2226,N_1946,N_1767);
nor U2227 (N_2227,N_1801,N_1794);
nor U2228 (N_2228,N_1809,N_1962);
and U2229 (N_2229,N_1813,N_1926);
or U2230 (N_2230,N_1947,N_1807);
or U2231 (N_2231,N_1894,N_1795);
and U2232 (N_2232,N_1811,N_1764);
and U2233 (N_2233,N_1780,N_1925);
or U2234 (N_2234,N_1994,N_1906);
and U2235 (N_2235,N_1993,N_1840);
nand U2236 (N_2236,N_1941,N_1974);
nand U2237 (N_2237,N_1754,N_1916);
or U2238 (N_2238,N_1991,N_1801);
nand U2239 (N_2239,N_1900,N_1936);
or U2240 (N_2240,N_1880,N_1833);
and U2241 (N_2241,N_1831,N_1903);
or U2242 (N_2242,N_1910,N_1988);
and U2243 (N_2243,N_1808,N_1965);
nand U2244 (N_2244,N_1798,N_1876);
and U2245 (N_2245,N_1767,N_1896);
or U2246 (N_2246,N_1796,N_1995);
xnor U2247 (N_2247,N_1871,N_1985);
and U2248 (N_2248,N_1957,N_1841);
xor U2249 (N_2249,N_1910,N_1832);
and U2250 (N_2250,N_2117,N_2086);
nand U2251 (N_2251,N_2077,N_2042);
and U2252 (N_2252,N_2065,N_2079);
or U2253 (N_2253,N_2124,N_2146);
nand U2254 (N_2254,N_2031,N_2191);
or U2255 (N_2255,N_2026,N_2165);
nand U2256 (N_2256,N_2168,N_2123);
nand U2257 (N_2257,N_2135,N_2180);
and U2258 (N_2258,N_2138,N_2033);
and U2259 (N_2259,N_2015,N_2132);
nor U2260 (N_2260,N_2099,N_2006);
nor U2261 (N_2261,N_2136,N_2056);
and U2262 (N_2262,N_2218,N_2047);
nor U2263 (N_2263,N_2110,N_2237);
and U2264 (N_2264,N_2049,N_2075);
nor U2265 (N_2265,N_2161,N_2160);
or U2266 (N_2266,N_2131,N_2024);
or U2267 (N_2267,N_2121,N_2013);
nand U2268 (N_2268,N_2116,N_2078);
and U2269 (N_2269,N_2204,N_2183);
or U2270 (N_2270,N_2069,N_2130);
or U2271 (N_2271,N_2201,N_2186);
nand U2272 (N_2272,N_2192,N_2109);
nand U2273 (N_2273,N_2236,N_2137);
and U2274 (N_2274,N_2092,N_2173);
nand U2275 (N_2275,N_2213,N_2224);
and U2276 (N_2276,N_2220,N_2166);
nand U2277 (N_2277,N_2149,N_2145);
nand U2278 (N_2278,N_2052,N_2067);
or U2279 (N_2279,N_2097,N_2045);
or U2280 (N_2280,N_2207,N_2030);
nand U2281 (N_2281,N_2139,N_2029);
or U2282 (N_2282,N_2169,N_2004);
or U2283 (N_2283,N_2177,N_2023);
or U2284 (N_2284,N_2001,N_2032);
nor U2285 (N_2285,N_2200,N_2061);
or U2286 (N_2286,N_2028,N_2058);
and U2287 (N_2287,N_2104,N_2157);
nand U2288 (N_2288,N_2090,N_2159);
nand U2289 (N_2289,N_2122,N_2059);
or U2290 (N_2290,N_2231,N_2153);
or U2291 (N_2291,N_2084,N_2232);
nand U2292 (N_2292,N_2007,N_2020);
and U2293 (N_2293,N_2223,N_2158);
or U2294 (N_2294,N_2009,N_2202);
nand U2295 (N_2295,N_2053,N_2151);
and U2296 (N_2296,N_2071,N_2195);
and U2297 (N_2297,N_2176,N_2081);
nand U2298 (N_2298,N_2048,N_2147);
or U2299 (N_2299,N_2193,N_2243);
and U2300 (N_2300,N_2102,N_2235);
or U2301 (N_2301,N_2039,N_2096);
or U2302 (N_2302,N_2127,N_2154);
or U2303 (N_2303,N_2179,N_2227);
and U2304 (N_2304,N_2219,N_2228);
or U2305 (N_2305,N_2167,N_2172);
nor U2306 (N_2306,N_2196,N_2206);
and U2307 (N_2307,N_2155,N_2120);
and U2308 (N_2308,N_2197,N_2025);
xnor U2309 (N_2309,N_2082,N_2114);
and U2310 (N_2310,N_2134,N_2118);
nand U2311 (N_2311,N_2246,N_2247);
or U2312 (N_2312,N_2095,N_2072);
or U2313 (N_2313,N_2057,N_2036);
or U2314 (N_2314,N_2062,N_2093);
or U2315 (N_2315,N_2005,N_2211);
and U2316 (N_2316,N_2239,N_2019);
nand U2317 (N_2317,N_2229,N_2010);
and U2318 (N_2318,N_2226,N_2073);
and U2319 (N_2319,N_2016,N_2216);
and U2320 (N_2320,N_2022,N_2054);
and U2321 (N_2321,N_2174,N_2230);
nor U2322 (N_2322,N_2119,N_2008);
xor U2323 (N_2323,N_2194,N_2106);
or U2324 (N_2324,N_2181,N_2021);
xor U2325 (N_2325,N_2163,N_2209);
and U2326 (N_2326,N_2101,N_2064);
or U2327 (N_2327,N_2152,N_2066);
and U2328 (N_2328,N_2162,N_2189);
and U2329 (N_2329,N_2068,N_2244);
or U2330 (N_2330,N_2060,N_2070);
or U2331 (N_2331,N_2000,N_2002);
nand U2332 (N_2332,N_2012,N_2222);
nand U2333 (N_2333,N_2044,N_2217);
and U2334 (N_2334,N_2043,N_2143);
or U2335 (N_2335,N_2215,N_2037);
and U2336 (N_2336,N_2034,N_2040);
nand U2337 (N_2337,N_2150,N_2094);
nor U2338 (N_2338,N_2063,N_2188);
nand U2339 (N_2339,N_2103,N_2187);
nor U2340 (N_2340,N_2249,N_2126);
or U2341 (N_2341,N_2221,N_2156);
or U2342 (N_2342,N_2234,N_2238);
and U2343 (N_2343,N_2115,N_2128);
or U2344 (N_2344,N_2164,N_2248);
or U2345 (N_2345,N_2199,N_2113);
and U2346 (N_2346,N_2170,N_2014);
nand U2347 (N_2347,N_2089,N_2027);
nand U2348 (N_2348,N_2242,N_2011);
xor U2349 (N_2349,N_2003,N_2046);
nand U2350 (N_2350,N_2125,N_2041);
xnor U2351 (N_2351,N_2087,N_2076);
and U2352 (N_2352,N_2175,N_2085);
nor U2353 (N_2353,N_2198,N_2233);
xnor U2354 (N_2354,N_2142,N_2203);
nor U2355 (N_2355,N_2141,N_2171);
nand U2356 (N_2356,N_2108,N_2140);
or U2357 (N_2357,N_2182,N_2148);
xnor U2358 (N_2358,N_2035,N_2038);
or U2359 (N_2359,N_2105,N_2055);
or U2360 (N_2360,N_2083,N_2210);
nor U2361 (N_2361,N_2017,N_2178);
xor U2362 (N_2362,N_2098,N_2088);
nand U2363 (N_2363,N_2091,N_2074);
and U2364 (N_2364,N_2080,N_2185);
and U2365 (N_2365,N_2107,N_2129);
and U2366 (N_2366,N_2205,N_2208);
or U2367 (N_2367,N_2144,N_2245);
nor U2368 (N_2368,N_2212,N_2214);
or U2369 (N_2369,N_2190,N_2111);
or U2370 (N_2370,N_2241,N_2051);
and U2371 (N_2371,N_2184,N_2240);
nand U2372 (N_2372,N_2225,N_2050);
nor U2373 (N_2373,N_2100,N_2133);
or U2374 (N_2374,N_2112,N_2018);
and U2375 (N_2375,N_2225,N_2079);
or U2376 (N_2376,N_2231,N_2007);
nand U2377 (N_2377,N_2017,N_2046);
nor U2378 (N_2378,N_2039,N_2205);
nand U2379 (N_2379,N_2173,N_2241);
or U2380 (N_2380,N_2096,N_2013);
nand U2381 (N_2381,N_2095,N_2204);
or U2382 (N_2382,N_2128,N_2157);
nor U2383 (N_2383,N_2032,N_2234);
nand U2384 (N_2384,N_2010,N_2050);
nand U2385 (N_2385,N_2180,N_2235);
and U2386 (N_2386,N_2161,N_2134);
nor U2387 (N_2387,N_2220,N_2062);
and U2388 (N_2388,N_2017,N_2247);
and U2389 (N_2389,N_2204,N_2178);
nor U2390 (N_2390,N_2231,N_2193);
and U2391 (N_2391,N_2054,N_2152);
and U2392 (N_2392,N_2163,N_2101);
and U2393 (N_2393,N_2174,N_2019);
and U2394 (N_2394,N_2043,N_2059);
or U2395 (N_2395,N_2207,N_2005);
or U2396 (N_2396,N_2133,N_2104);
or U2397 (N_2397,N_2249,N_2186);
or U2398 (N_2398,N_2126,N_2245);
and U2399 (N_2399,N_2162,N_2006);
nand U2400 (N_2400,N_2008,N_2231);
or U2401 (N_2401,N_2101,N_2083);
or U2402 (N_2402,N_2054,N_2212);
or U2403 (N_2403,N_2134,N_2207);
nand U2404 (N_2404,N_2072,N_2032);
nor U2405 (N_2405,N_2046,N_2149);
nor U2406 (N_2406,N_2104,N_2065);
or U2407 (N_2407,N_2041,N_2055);
xor U2408 (N_2408,N_2046,N_2168);
or U2409 (N_2409,N_2011,N_2129);
nand U2410 (N_2410,N_2210,N_2231);
and U2411 (N_2411,N_2133,N_2174);
nand U2412 (N_2412,N_2072,N_2031);
nor U2413 (N_2413,N_2098,N_2117);
or U2414 (N_2414,N_2126,N_2201);
xor U2415 (N_2415,N_2026,N_2064);
or U2416 (N_2416,N_2176,N_2112);
and U2417 (N_2417,N_2166,N_2140);
nor U2418 (N_2418,N_2034,N_2112);
nand U2419 (N_2419,N_2177,N_2157);
and U2420 (N_2420,N_2095,N_2089);
and U2421 (N_2421,N_2174,N_2231);
and U2422 (N_2422,N_2092,N_2017);
nand U2423 (N_2423,N_2203,N_2138);
or U2424 (N_2424,N_2163,N_2116);
nor U2425 (N_2425,N_2215,N_2073);
nand U2426 (N_2426,N_2027,N_2082);
and U2427 (N_2427,N_2231,N_2229);
nand U2428 (N_2428,N_2090,N_2209);
xor U2429 (N_2429,N_2209,N_2164);
nand U2430 (N_2430,N_2189,N_2172);
nand U2431 (N_2431,N_2086,N_2120);
and U2432 (N_2432,N_2158,N_2238);
nor U2433 (N_2433,N_2173,N_2060);
and U2434 (N_2434,N_2089,N_2203);
nor U2435 (N_2435,N_2154,N_2068);
or U2436 (N_2436,N_2245,N_2182);
and U2437 (N_2437,N_2160,N_2246);
and U2438 (N_2438,N_2047,N_2214);
nor U2439 (N_2439,N_2172,N_2185);
nand U2440 (N_2440,N_2026,N_2051);
nor U2441 (N_2441,N_2177,N_2114);
nor U2442 (N_2442,N_2068,N_2200);
nor U2443 (N_2443,N_2202,N_2152);
and U2444 (N_2444,N_2186,N_2033);
nand U2445 (N_2445,N_2144,N_2176);
or U2446 (N_2446,N_2089,N_2115);
nand U2447 (N_2447,N_2087,N_2089);
or U2448 (N_2448,N_2157,N_2091);
nor U2449 (N_2449,N_2105,N_2102);
and U2450 (N_2450,N_2210,N_2103);
or U2451 (N_2451,N_2022,N_2246);
and U2452 (N_2452,N_2192,N_2193);
nand U2453 (N_2453,N_2193,N_2080);
nor U2454 (N_2454,N_2184,N_2177);
and U2455 (N_2455,N_2209,N_2011);
or U2456 (N_2456,N_2223,N_2226);
nand U2457 (N_2457,N_2181,N_2220);
and U2458 (N_2458,N_2131,N_2009);
or U2459 (N_2459,N_2197,N_2097);
nand U2460 (N_2460,N_2036,N_2092);
or U2461 (N_2461,N_2175,N_2158);
or U2462 (N_2462,N_2158,N_2189);
and U2463 (N_2463,N_2103,N_2177);
nand U2464 (N_2464,N_2105,N_2179);
or U2465 (N_2465,N_2226,N_2037);
or U2466 (N_2466,N_2117,N_2092);
xor U2467 (N_2467,N_2036,N_2169);
and U2468 (N_2468,N_2120,N_2217);
nand U2469 (N_2469,N_2149,N_2213);
nor U2470 (N_2470,N_2083,N_2053);
or U2471 (N_2471,N_2192,N_2022);
and U2472 (N_2472,N_2107,N_2092);
xnor U2473 (N_2473,N_2094,N_2177);
nand U2474 (N_2474,N_2194,N_2066);
or U2475 (N_2475,N_2155,N_2198);
and U2476 (N_2476,N_2057,N_2025);
nor U2477 (N_2477,N_2071,N_2016);
and U2478 (N_2478,N_2238,N_2156);
or U2479 (N_2479,N_2064,N_2062);
and U2480 (N_2480,N_2202,N_2179);
nand U2481 (N_2481,N_2052,N_2144);
or U2482 (N_2482,N_2121,N_2005);
nor U2483 (N_2483,N_2115,N_2105);
and U2484 (N_2484,N_2076,N_2230);
and U2485 (N_2485,N_2046,N_2123);
nor U2486 (N_2486,N_2134,N_2243);
and U2487 (N_2487,N_2177,N_2189);
nor U2488 (N_2488,N_2100,N_2082);
or U2489 (N_2489,N_2003,N_2215);
and U2490 (N_2490,N_2154,N_2077);
nand U2491 (N_2491,N_2235,N_2192);
or U2492 (N_2492,N_2200,N_2157);
nor U2493 (N_2493,N_2207,N_2066);
nand U2494 (N_2494,N_2126,N_2105);
or U2495 (N_2495,N_2050,N_2083);
and U2496 (N_2496,N_2018,N_2186);
nand U2497 (N_2497,N_2176,N_2047);
nor U2498 (N_2498,N_2134,N_2125);
and U2499 (N_2499,N_2233,N_2156);
nand U2500 (N_2500,N_2292,N_2308);
or U2501 (N_2501,N_2400,N_2337);
nand U2502 (N_2502,N_2475,N_2255);
and U2503 (N_2503,N_2464,N_2284);
and U2504 (N_2504,N_2455,N_2268);
and U2505 (N_2505,N_2376,N_2382);
nand U2506 (N_2506,N_2346,N_2494);
nand U2507 (N_2507,N_2277,N_2296);
xnor U2508 (N_2508,N_2351,N_2338);
and U2509 (N_2509,N_2413,N_2339);
nor U2510 (N_2510,N_2440,N_2332);
and U2511 (N_2511,N_2417,N_2407);
and U2512 (N_2512,N_2425,N_2428);
and U2513 (N_2513,N_2412,N_2435);
or U2514 (N_2514,N_2399,N_2409);
nor U2515 (N_2515,N_2433,N_2340);
nand U2516 (N_2516,N_2359,N_2327);
and U2517 (N_2517,N_2418,N_2343);
or U2518 (N_2518,N_2374,N_2401);
nand U2519 (N_2519,N_2426,N_2481);
nor U2520 (N_2520,N_2488,N_2270);
and U2521 (N_2521,N_2474,N_2442);
nor U2522 (N_2522,N_2469,N_2403);
nor U2523 (N_2523,N_2498,N_2257);
and U2524 (N_2524,N_2406,N_2321);
nor U2525 (N_2525,N_2457,N_2436);
nand U2526 (N_2526,N_2465,N_2405);
and U2527 (N_2527,N_2356,N_2253);
and U2528 (N_2528,N_2370,N_2458);
or U2529 (N_2529,N_2489,N_2303);
and U2530 (N_2530,N_2453,N_2306);
nor U2531 (N_2531,N_2463,N_2259);
nor U2532 (N_2532,N_2393,N_2483);
or U2533 (N_2533,N_2402,N_2291);
and U2534 (N_2534,N_2349,N_2362);
nor U2535 (N_2535,N_2477,N_2294);
nand U2536 (N_2536,N_2493,N_2383);
or U2537 (N_2537,N_2468,N_2431);
and U2538 (N_2538,N_2476,N_2318);
or U2539 (N_2539,N_2484,N_2454);
nor U2540 (N_2540,N_2288,N_2365);
nand U2541 (N_2541,N_2377,N_2471);
nand U2542 (N_2542,N_2446,N_2293);
nand U2543 (N_2543,N_2491,N_2368);
nor U2544 (N_2544,N_2312,N_2326);
nor U2545 (N_2545,N_2432,N_2279);
and U2546 (N_2546,N_2280,N_2492);
and U2547 (N_2547,N_2275,N_2396);
nor U2548 (N_2548,N_2381,N_2371);
nor U2549 (N_2549,N_2419,N_2414);
nor U2550 (N_2550,N_2366,N_2473);
nor U2551 (N_2551,N_2364,N_2490);
nand U2552 (N_2552,N_2252,N_2311);
nor U2553 (N_2553,N_2322,N_2415);
or U2554 (N_2554,N_2427,N_2324);
and U2555 (N_2555,N_2387,N_2314);
and U2556 (N_2556,N_2388,N_2444);
or U2557 (N_2557,N_2404,N_2301);
and U2558 (N_2558,N_2267,N_2251);
xor U2559 (N_2559,N_2485,N_2459);
and U2560 (N_2560,N_2335,N_2434);
nand U2561 (N_2561,N_2379,N_2304);
or U2562 (N_2562,N_2375,N_2445);
or U2563 (N_2563,N_2353,N_2384);
nor U2564 (N_2564,N_2341,N_2302);
or U2565 (N_2565,N_2348,N_2369);
nor U2566 (N_2566,N_2470,N_2452);
and U2567 (N_2567,N_2334,N_2422);
nor U2568 (N_2568,N_2397,N_2472);
nand U2569 (N_2569,N_2439,N_2347);
or U2570 (N_2570,N_2336,N_2297);
nand U2571 (N_2571,N_2299,N_2298);
nor U2572 (N_2572,N_2269,N_2367);
and U2573 (N_2573,N_2395,N_2315);
and U2574 (N_2574,N_2316,N_2256);
nand U2575 (N_2575,N_2263,N_2380);
nor U2576 (N_2576,N_2378,N_2286);
nand U2577 (N_2577,N_2386,N_2354);
and U2578 (N_2578,N_2250,N_2310);
and U2579 (N_2579,N_2420,N_2305);
and U2580 (N_2580,N_2271,N_2456);
nand U2581 (N_2581,N_2438,N_2295);
or U2582 (N_2582,N_2441,N_2258);
nor U2583 (N_2583,N_2276,N_2479);
and U2584 (N_2584,N_2342,N_2449);
and U2585 (N_2585,N_2429,N_2330);
or U2586 (N_2586,N_2352,N_2320);
nand U2587 (N_2587,N_2467,N_2462);
nor U2588 (N_2588,N_2265,N_2329);
xnor U2589 (N_2589,N_2482,N_2423);
and U2590 (N_2590,N_2272,N_2461);
or U2591 (N_2591,N_2283,N_2450);
and U2592 (N_2592,N_2478,N_2285);
and U2593 (N_2593,N_2430,N_2497);
nor U2594 (N_2594,N_2254,N_2460);
nand U2595 (N_2595,N_2421,N_2355);
or U2596 (N_2596,N_2281,N_2451);
or U2597 (N_2597,N_2373,N_2363);
or U2598 (N_2598,N_2448,N_2443);
xnor U2599 (N_2599,N_2390,N_2389);
and U2600 (N_2600,N_2410,N_2328);
nor U2601 (N_2601,N_2408,N_2411);
nor U2602 (N_2602,N_2344,N_2319);
nand U2603 (N_2603,N_2290,N_2307);
and U2604 (N_2604,N_2437,N_2260);
or U2605 (N_2605,N_2360,N_2278);
and U2606 (N_2606,N_2447,N_2274);
nor U2607 (N_2607,N_2499,N_2394);
and U2608 (N_2608,N_2466,N_2262);
nor U2609 (N_2609,N_2317,N_2416);
nor U2610 (N_2610,N_2273,N_2350);
nand U2611 (N_2611,N_2264,N_2289);
or U2612 (N_2612,N_2372,N_2261);
nand U2613 (N_2613,N_2323,N_2331);
nor U2614 (N_2614,N_2345,N_2325);
nor U2615 (N_2615,N_2398,N_2391);
or U2616 (N_2616,N_2282,N_2495);
nand U2617 (N_2617,N_2385,N_2487);
nand U2618 (N_2618,N_2300,N_2392);
nor U2619 (N_2619,N_2266,N_2358);
nand U2620 (N_2620,N_2496,N_2313);
or U2621 (N_2621,N_2424,N_2287);
and U2622 (N_2622,N_2309,N_2333);
nand U2623 (N_2623,N_2480,N_2357);
xnor U2624 (N_2624,N_2486,N_2361);
nor U2625 (N_2625,N_2422,N_2491);
or U2626 (N_2626,N_2394,N_2296);
or U2627 (N_2627,N_2375,N_2374);
and U2628 (N_2628,N_2437,N_2418);
and U2629 (N_2629,N_2265,N_2496);
and U2630 (N_2630,N_2357,N_2261);
and U2631 (N_2631,N_2274,N_2317);
and U2632 (N_2632,N_2337,N_2270);
nand U2633 (N_2633,N_2339,N_2414);
or U2634 (N_2634,N_2408,N_2491);
and U2635 (N_2635,N_2270,N_2394);
nor U2636 (N_2636,N_2364,N_2415);
or U2637 (N_2637,N_2316,N_2288);
nor U2638 (N_2638,N_2333,N_2431);
or U2639 (N_2639,N_2479,N_2343);
nor U2640 (N_2640,N_2288,N_2359);
or U2641 (N_2641,N_2402,N_2367);
or U2642 (N_2642,N_2393,N_2351);
or U2643 (N_2643,N_2298,N_2371);
and U2644 (N_2644,N_2369,N_2434);
nor U2645 (N_2645,N_2421,N_2425);
and U2646 (N_2646,N_2309,N_2384);
and U2647 (N_2647,N_2394,N_2322);
or U2648 (N_2648,N_2260,N_2477);
or U2649 (N_2649,N_2327,N_2294);
or U2650 (N_2650,N_2387,N_2352);
and U2651 (N_2651,N_2264,N_2297);
or U2652 (N_2652,N_2397,N_2453);
nor U2653 (N_2653,N_2284,N_2428);
and U2654 (N_2654,N_2486,N_2401);
nor U2655 (N_2655,N_2373,N_2381);
xor U2656 (N_2656,N_2496,N_2452);
and U2657 (N_2657,N_2492,N_2257);
or U2658 (N_2658,N_2335,N_2322);
nand U2659 (N_2659,N_2423,N_2492);
and U2660 (N_2660,N_2342,N_2310);
and U2661 (N_2661,N_2286,N_2435);
and U2662 (N_2662,N_2264,N_2321);
or U2663 (N_2663,N_2324,N_2330);
or U2664 (N_2664,N_2299,N_2270);
and U2665 (N_2665,N_2486,N_2431);
and U2666 (N_2666,N_2409,N_2280);
or U2667 (N_2667,N_2406,N_2400);
and U2668 (N_2668,N_2492,N_2363);
nand U2669 (N_2669,N_2297,N_2353);
and U2670 (N_2670,N_2435,N_2284);
and U2671 (N_2671,N_2334,N_2494);
or U2672 (N_2672,N_2360,N_2398);
and U2673 (N_2673,N_2491,N_2359);
nor U2674 (N_2674,N_2320,N_2262);
and U2675 (N_2675,N_2315,N_2454);
or U2676 (N_2676,N_2454,N_2496);
nor U2677 (N_2677,N_2410,N_2363);
nor U2678 (N_2678,N_2326,N_2306);
nor U2679 (N_2679,N_2352,N_2343);
and U2680 (N_2680,N_2334,N_2395);
or U2681 (N_2681,N_2261,N_2426);
nor U2682 (N_2682,N_2280,N_2415);
nand U2683 (N_2683,N_2385,N_2272);
nor U2684 (N_2684,N_2258,N_2359);
nand U2685 (N_2685,N_2489,N_2453);
nor U2686 (N_2686,N_2325,N_2450);
and U2687 (N_2687,N_2449,N_2430);
or U2688 (N_2688,N_2308,N_2486);
nand U2689 (N_2689,N_2253,N_2361);
nand U2690 (N_2690,N_2336,N_2485);
and U2691 (N_2691,N_2329,N_2467);
or U2692 (N_2692,N_2447,N_2303);
nand U2693 (N_2693,N_2396,N_2361);
nor U2694 (N_2694,N_2328,N_2285);
or U2695 (N_2695,N_2467,N_2396);
nand U2696 (N_2696,N_2371,N_2397);
and U2697 (N_2697,N_2331,N_2452);
and U2698 (N_2698,N_2492,N_2289);
nor U2699 (N_2699,N_2333,N_2328);
or U2700 (N_2700,N_2391,N_2491);
or U2701 (N_2701,N_2380,N_2309);
nor U2702 (N_2702,N_2492,N_2286);
and U2703 (N_2703,N_2320,N_2484);
nand U2704 (N_2704,N_2395,N_2316);
nor U2705 (N_2705,N_2430,N_2446);
and U2706 (N_2706,N_2471,N_2397);
and U2707 (N_2707,N_2270,N_2498);
nand U2708 (N_2708,N_2454,N_2277);
nand U2709 (N_2709,N_2448,N_2289);
and U2710 (N_2710,N_2491,N_2381);
xnor U2711 (N_2711,N_2361,N_2462);
or U2712 (N_2712,N_2332,N_2471);
nor U2713 (N_2713,N_2389,N_2320);
and U2714 (N_2714,N_2484,N_2334);
or U2715 (N_2715,N_2460,N_2379);
and U2716 (N_2716,N_2282,N_2373);
or U2717 (N_2717,N_2331,N_2289);
or U2718 (N_2718,N_2316,N_2340);
and U2719 (N_2719,N_2424,N_2455);
or U2720 (N_2720,N_2251,N_2444);
and U2721 (N_2721,N_2334,N_2477);
or U2722 (N_2722,N_2395,N_2279);
or U2723 (N_2723,N_2322,N_2468);
nand U2724 (N_2724,N_2315,N_2334);
or U2725 (N_2725,N_2277,N_2378);
nand U2726 (N_2726,N_2272,N_2387);
nor U2727 (N_2727,N_2263,N_2462);
or U2728 (N_2728,N_2250,N_2362);
nand U2729 (N_2729,N_2450,N_2467);
or U2730 (N_2730,N_2360,N_2299);
and U2731 (N_2731,N_2380,N_2356);
nand U2732 (N_2732,N_2394,N_2496);
nand U2733 (N_2733,N_2416,N_2418);
or U2734 (N_2734,N_2373,N_2263);
nor U2735 (N_2735,N_2347,N_2252);
and U2736 (N_2736,N_2388,N_2412);
nor U2737 (N_2737,N_2356,N_2454);
and U2738 (N_2738,N_2475,N_2489);
nand U2739 (N_2739,N_2361,N_2269);
and U2740 (N_2740,N_2355,N_2433);
or U2741 (N_2741,N_2424,N_2428);
nand U2742 (N_2742,N_2348,N_2489);
or U2743 (N_2743,N_2441,N_2288);
nand U2744 (N_2744,N_2297,N_2398);
nand U2745 (N_2745,N_2309,N_2408);
or U2746 (N_2746,N_2270,N_2402);
nor U2747 (N_2747,N_2298,N_2319);
nor U2748 (N_2748,N_2487,N_2388);
nand U2749 (N_2749,N_2476,N_2378);
nand U2750 (N_2750,N_2619,N_2616);
nand U2751 (N_2751,N_2704,N_2567);
or U2752 (N_2752,N_2581,N_2516);
nand U2753 (N_2753,N_2720,N_2590);
nor U2754 (N_2754,N_2549,N_2710);
nand U2755 (N_2755,N_2733,N_2657);
or U2756 (N_2756,N_2559,N_2613);
nand U2757 (N_2757,N_2614,N_2682);
and U2758 (N_2758,N_2659,N_2635);
nand U2759 (N_2759,N_2738,N_2622);
nor U2760 (N_2760,N_2700,N_2637);
or U2761 (N_2761,N_2563,N_2542);
nor U2762 (N_2762,N_2669,N_2585);
nor U2763 (N_2763,N_2553,N_2633);
nand U2764 (N_2764,N_2660,N_2664);
nor U2765 (N_2765,N_2521,N_2577);
and U2766 (N_2766,N_2534,N_2650);
nor U2767 (N_2767,N_2706,N_2529);
or U2768 (N_2768,N_2519,N_2598);
nor U2769 (N_2769,N_2522,N_2557);
nand U2770 (N_2770,N_2560,N_2574);
nor U2771 (N_2771,N_2501,N_2628);
nand U2772 (N_2772,N_2746,N_2535);
or U2773 (N_2773,N_2644,N_2552);
nand U2774 (N_2774,N_2566,N_2742);
or U2775 (N_2775,N_2596,N_2599);
nor U2776 (N_2776,N_2690,N_2556);
nand U2777 (N_2777,N_2718,N_2672);
nor U2778 (N_2778,N_2502,N_2508);
or U2779 (N_2779,N_2667,N_2643);
nand U2780 (N_2780,N_2589,N_2748);
or U2781 (N_2781,N_2680,N_2564);
and U2782 (N_2782,N_2580,N_2550);
and U2783 (N_2783,N_2554,N_2514);
and U2784 (N_2784,N_2532,N_2693);
nand U2785 (N_2785,N_2523,N_2601);
nand U2786 (N_2786,N_2517,N_2568);
nor U2787 (N_2787,N_2597,N_2716);
nor U2788 (N_2788,N_2578,N_2732);
nand U2789 (N_2789,N_2608,N_2604);
nor U2790 (N_2790,N_2695,N_2715);
and U2791 (N_2791,N_2636,N_2576);
nor U2792 (N_2792,N_2707,N_2668);
nand U2793 (N_2793,N_2545,N_2562);
nor U2794 (N_2794,N_2717,N_2737);
nor U2795 (N_2795,N_2651,N_2586);
nand U2796 (N_2796,N_2593,N_2561);
and U2797 (N_2797,N_2739,N_2687);
and U2798 (N_2798,N_2677,N_2731);
nand U2799 (N_2799,N_2620,N_2654);
nor U2800 (N_2800,N_2705,N_2642);
nand U2801 (N_2801,N_2536,N_2684);
or U2802 (N_2802,N_2740,N_2671);
and U2803 (N_2803,N_2656,N_2624);
or U2804 (N_2804,N_2530,N_2675);
or U2805 (N_2805,N_2551,N_2623);
or U2806 (N_2806,N_2531,N_2697);
and U2807 (N_2807,N_2520,N_2524);
nor U2808 (N_2808,N_2629,N_2526);
and U2809 (N_2809,N_2594,N_2509);
and U2810 (N_2810,N_2634,N_2541);
or U2811 (N_2811,N_2692,N_2658);
nor U2812 (N_2812,N_2600,N_2728);
and U2813 (N_2813,N_2506,N_2688);
nor U2814 (N_2814,N_2708,N_2749);
nor U2815 (N_2815,N_2673,N_2714);
and U2816 (N_2816,N_2632,N_2670);
nand U2817 (N_2817,N_2539,N_2648);
and U2818 (N_2818,N_2741,N_2546);
and U2819 (N_2819,N_2582,N_2666);
nand U2820 (N_2820,N_2736,N_2543);
nand U2821 (N_2821,N_2745,N_2518);
nor U2822 (N_2822,N_2579,N_2612);
nand U2823 (N_2823,N_2711,N_2699);
or U2824 (N_2824,N_2538,N_2515);
nand U2825 (N_2825,N_2730,N_2725);
nand U2826 (N_2826,N_2558,N_2681);
nand U2827 (N_2827,N_2694,N_2572);
nor U2828 (N_2828,N_2662,N_2565);
nor U2829 (N_2829,N_2595,N_2721);
nand U2830 (N_2830,N_2641,N_2647);
nand U2831 (N_2831,N_2587,N_2544);
nor U2832 (N_2832,N_2592,N_2617);
and U2833 (N_2833,N_2510,N_2645);
or U2834 (N_2834,N_2723,N_2630);
nand U2835 (N_2835,N_2685,N_2591);
and U2836 (N_2836,N_2663,N_2625);
and U2837 (N_2837,N_2609,N_2655);
and U2838 (N_2838,N_2719,N_2665);
nor U2839 (N_2839,N_2603,N_2689);
nand U2840 (N_2840,N_2686,N_2744);
nor U2841 (N_2841,N_2584,N_2638);
and U2842 (N_2842,N_2573,N_2607);
and U2843 (N_2843,N_2621,N_2555);
nor U2844 (N_2844,N_2627,N_2505);
nand U2845 (N_2845,N_2500,N_2703);
nand U2846 (N_2846,N_2674,N_2734);
and U2847 (N_2847,N_2513,N_2702);
xnor U2848 (N_2848,N_2652,N_2512);
and U2849 (N_2849,N_2507,N_2639);
or U2850 (N_2850,N_2569,N_2583);
and U2851 (N_2851,N_2709,N_2712);
nor U2852 (N_2852,N_2602,N_2571);
and U2853 (N_2853,N_2611,N_2649);
and U2854 (N_2854,N_2615,N_2678);
nor U2855 (N_2855,N_2722,N_2646);
and U2856 (N_2856,N_2713,N_2726);
and U2857 (N_2857,N_2503,N_2575);
nor U2858 (N_2858,N_2606,N_2605);
nand U2859 (N_2859,N_2588,N_2548);
or U2860 (N_2860,N_2525,N_2511);
and U2861 (N_2861,N_2724,N_2540);
and U2862 (N_2862,N_2735,N_2743);
or U2863 (N_2863,N_2618,N_2679);
nor U2864 (N_2864,N_2528,N_2701);
and U2865 (N_2865,N_2504,N_2747);
and U2866 (N_2866,N_2729,N_2653);
nor U2867 (N_2867,N_2547,N_2626);
or U2868 (N_2868,N_2691,N_2533);
or U2869 (N_2869,N_2698,N_2610);
or U2870 (N_2870,N_2537,N_2696);
nor U2871 (N_2871,N_2727,N_2631);
nor U2872 (N_2872,N_2661,N_2640);
nor U2873 (N_2873,N_2527,N_2570);
or U2874 (N_2874,N_2683,N_2676);
or U2875 (N_2875,N_2649,N_2703);
nand U2876 (N_2876,N_2559,N_2663);
and U2877 (N_2877,N_2708,N_2601);
or U2878 (N_2878,N_2504,N_2708);
and U2879 (N_2879,N_2685,N_2728);
and U2880 (N_2880,N_2577,N_2594);
nand U2881 (N_2881,N_2668,N_2609);
and U2882 (N_2882,N_2748,N_2600);
nor U2883 (N_2883,N_2561,N_2584);
nand U2884 (N_2884,N_2682,N_2597);
or U2885 (N_2885,N_2725,N_2693);
or U2886 (N_2886,N_2594,N_2525);
and U2887 (N_2887,N_2508,N_2668);
nand U2888 (N_2888,N_2612,N_2697);
and U2889 (N_2889,N_2635,N_2717);
and U2890 (N_2890,N_2649,N_2559);
or U2891 (N_2891,N_2626,N_2532);
nor U2892 (N_2892,N_2609,N_2645);
xnor U2893 (N_2893,N_2710,N_2572);
nand U2894 (N_2894,N_2732,N_2646);
and U2895 (N_2895,N_2563,N_2547);
nand U2896 (N_2896,N_2516,N_2738);
nand U2897 (N_2897,N_2666,N_2538);
or U2898 (N_2898,N_2746,N_2662);
xnor U2899 (N_2899,N_2532,N_2657);
nand U2900 (N_2900,N_2541,N_2676);
or U2901 (N_2901,N_2644,N_2526);
nor U2902 (N_2902,N_2637,N_2629);
or U2903 (N_2903,N_2664,N_2550);
or U2904 (N_2904,N_2730,N_2658);
xor U2905 (N_2905,N_2648,N_2684);
nand U2906 (N_2906,N_2528,N_2620);
nor U2907 (N_2907,N_2510,N_2648);
nor U2908 (N_2908,N_2628,N_2729);
nor U2909 (N_2909,N_2623,N_2574);
nand U2910 (N_2910,N_2665,N_2720);
or U2911 (N_2911,N_2705,N_2522);
or U2912 (N_2912,N_2688,N_2666);
or U2913 (N_2913,N_2575,N_2692);
or U2914 (N_2914,N_2700,N_2733);
nand U2915 (N_2915,N_2593,N_2733);
and U2916 (N_2916,N_2629,N_2573);
or U2917 (N_2917,N_2697,N_2593);
or U2918 (N_2918,N_2749,N_2540);
nor U2919 (N_2919,N_2583,N_2681);
nand U2920 (N_2920,N_2501,N_2706);
and U2921 (N_2921,N_2617,N_2565);
and U2922 (N_2922,N_2549,N_2523);
and U2923 (N_2923,N_2679,N_2717);
and U2924 (N_2924,N_2626,N_2546);
or U2925 (N_2925,N_2609,N_2546);
nand U2926 (N_2926,N_2585,N_2572);
nor U2927 (N_2927,N_2517,N_2681);
and U2928 (N_2928,N_2686,N_2677);
nor U2929 (N_2929,N_2653,N_2587);
nor U2930 (N_2930,N_2728,N_2629);
and U2931 (N_2931,N_2500,N_2648);
nand U2932 (N_2932,N_2552,N_2520);
or U2933 (N_2933,N_2591,N_2713);
nor U2934 (N_2934,N_2586,N_2659);
nand U2935 (N_2935,N_2573,N_2723);
nor U2936 (N_2936,N_2719,N_2600);
nor U2937 (N_2937,N_2527,N_2684);
nor U2938 (N_2938,N_2672,N_2562);
and U2939 (N_2939,N_2593,N_2724);
and U2940 (N_2940,N_2514,N_2629);
or U2941 (N_2941,N_2683,N_2713);
nand U2942 (N_2942,N_2515,N_2599);
and U2943 (N_2943,N_2648,N_2593);
nand U2944 (N_2944,N_2557,N_2620);
and U2945 (N_2945,N_2645,N_2541);
xnor U2946 (N_2946,N_2684,N_2729);
or U2947 (N_2947,N_2587,N_2633);
or U2948 (N_2948,N_2524,N_2661);
or U2949 (N_2949,N_2670,N_2668);
nand U2950 (N_2950,N_2636,N_2695);
or U2951 (N_2951,N_2592,N_2633);
nand U2952 (N_2952,N_2557,N_2595);
nor U2953 (N_2953,N_2595,N_2671);
or U2954 (N_2954,N_2643,N_2620);
and U2955 (N_2955,N_2559,N_2701);
or U2956 (N_2956,N_2551,N_2502);
and U2957 (N_2957,N_2620,N_2721);
nand U2958 (N_2958,N_2507,N_2714);
and U2959 (N_2959,N_2708,N_2736);
nor U2960 (N_2960,N_2725,N_2549);
nand U2961 (N_2961,N_2630,N_2717);
nand U2962 (N_2962,N_2636,N_2550);
and U2963 (N_2963,N_2608,N_2586);
or U2964 (N_2964,N_2629,N_2570);
nor U2965 (N_2965,N_2664,N_2529);
or U2966 (N_2966,N_2669,N_2541);
nand U2967 (N_2967,N_2511,N_2746);
and U2968 (N_2968,N_2739,N_2588);
and U2969 (N_2969,N_2520,N_2713);
nand U2970 (N_2970,N_2651,N_2666);
xor U2971 (N_2971,N_2659,N_2508);
nand U2972 (N_2972,N_2655,N_2652);
nor U2973 (N_2973,N_2689,N_2540);
nor U2974 (N_2974,N_2596,N_2654);
or U2975 (N_2975,N_2606,N_2718);
nor U2976 (N_2976,N_2624,N_2593);
or U2977 (N_2977,N_2729,N_2608);
and U2978 (N_2978,N_2519,N_2655);
nand U2979 (N_2979,N_2717,N_2659);
and U2980 (N_2980,N_2534,N_2590);
nand U2981 (N_2981,N_2531,N_2615);
nor U2982 (N_2982,N_2545,N_2599);
nor U2983 (N_2983,N_2562,N_2658);
nand U2984 (N_2984,N_2693,N_2664);
xor U2985 (N_2985,N_2650,N_2616);
or U2986 (N_2986,N_2601,N_2551);
and U2987 (N_2987,N_2614,N_2571);
and U2988 (N_2988,N_2703,N_2590);
nand U2989 (N_2989,N_2663,N_2512);
and U2990 (N_2990,N_2732,N_2659);
or U2991 (N_2991,N_2643,N_2571);
or U2992 (N_2992,N_2538,N_2727);
or U2993 (N_2993,N_2747,N_2598);
nor U2994 (N_2994,N_2615,N_2742);
nand U2995 (N_2995,N_2500,N_2730);
and U2996 (N_2996,N_2684,N_2740);
nand U2997 (N_2997,N_2647,N_2673);
and U2998 (N_2998,N_2678,N_2528);
or U2999 (N_2999,N_2658,N_2724);
and U3000 (N_3000,N_2917,N_2910);
or U3001 (N_3001,N_2802,N_2789);
and U3002 (N_3002,N_2860,N_2896);
nand U3003 (N_3003,N_2969,N_2766);
nand U3004 (N_3004,N_2924,N_2768);
nor U3005 (N_3005,N_2893,N_2778);
and U3006 (N_3006,N_2817,N_2866);
or U3007 (N_3007,N_2812,N_2947);
or U3008 (N_3008,N_2929,N_2763);
nand U3009 (N_3009,N_2788,N_2964);
or U3010 (N_3010,N_2993,N_2750);
and U3011 (N_3011,N_2983,N_2875);
or U3012 (N_3012,N_2940,N_2858);
nand U3013 (N_3013,N_2878,N_2882);
and U3014 (N_3014,N_2939,N_2867);
nor U3015 (N_3015,N_2876,N_2977);
nor U3016 (N_3016,N_2765,N_2863);
nor U3017 (N_3017,N_2805,N_2982);
or U3018 (N_3018,N_2755,N_2989);
and U3019 (N_3019,N_2773,N_2770);
or U3020 (N_3020,N_2962,N_2928);
nor U3021 (N_3021,N_2997,N_2897);
nand U3022 (N_3022,N_2963,N_2854);
nor U3023 (N_3023,N_2849,N_2790);
nand U3024 (N_3024,N_2829,N_2791);
xnor U3025 (N_3025,N_2864,N_2957);
nand U3026 (N_3026,N_2811,N_2974);
nand U3027 (N_3027,N_2880,N_2925);
nand U3028 (N_3028,N_2984,N_2921);
or U3029 (N_3029,N_2818,N_2938);
nor U3030 (N_3030,N_2777,N_2948);
and U3031 (N_3031,N_2869,N_2764);
nand U3032 (N_3032,N_2988,N_2753);
and U3033 (N_3033,N_2810,N_2760);
and U3034 (N_3034,N_2954,N_2841);
nand U3035 (N_3035,N_2752,N_2877);
nor U3036 (N_3036,N_2754,N_2949);
nor U3037 (N_3037,N_2767,N_2815);
nand U3038 (N_3038,N_2937,N_2952);
nor U3039 (N_3039,N_2950,N_2992);
or U3040 (N_3040,N_2907,N_2757);
nor U3041 (N_3041,N_2990,N_2853);
or U3042 (N_3042,N_2779,N_2965);
nor U3043 (N_3043,N_2881,N_2855);
and U3044 (N_3044,N_2851,N_2759);
and U3045 (N_3045,N_2830,N_2834);
nor U3046 (N_3046,N_2831,N_2865);
or U3047 (N_3047,N_2976,N_2933);
or U3048 (N_3048,N_2825,N_2839);
and U3049 (N_3049,N_2906,N_2919);
and U3050 (N_3050,N_2926,N_2951);
nand U3051 (N_3051,N_2874,N_2905);
nor U3052 (N_3052,N_2944,N_2783);
and U3053 (N_3053,N_2932,N_2889);
nor U3054 (N_3054,N_2769,N_2991);
nor U3055 (N_3055,N_2883,N_2935);
nor U3056 (N_3056,N_2968,N_2959);
or U3057 (N_3057,N_2895,N_2967);
nand U3058 (N_3058,N_2842,N_2918);
and U3059 (N_3059,N_2902,N_2973);
and U3060 (N_3060,N_2985,N_2971);
and U3061 (N_3061,N_2793,N_2823);
and U3062 (N_3062,N_2941,N_2972);
and U3063 (N_3063,N_2843,N_2814);
or U3064 (N_3064,N_2978,N_2792);
nand U3065 (N_3065,N_2872,N_2886);
or U3066 (N_3066,N_2786,N_2885);
or U3067 (N_3067,N_2821,N_2870);
nor U3068 (N_3068,N_2958,N_2794);
and U3069 (N_3069,N_2879,N_2931);
nand U3070 (N_3070,N_2837,N_2994);
or U3071 (N_3071,N_2943,N_2761);
nand U3072 (N_3072,N_2888,N_2975);
and U3073 (N_3073,N_2832,N_2887);
nor U3074 (N_3074,N_2912,N_2801);
or U3075 (N_3075,N_2809,N_2966);
nor U3076 (N_3076,N_2936,N_2771);
and U3077 (N_3077,N_2900,N_2840);
nor U3078 (N_3078,N_2822,N_2780);
and U3079 (N_3079,N_2758,N_2857);
and U3080 (N_3080,N_2844,N_2915);
and U3081 (N_3081,N_2946,N_2953);
and U3082 (N_3082,N_2942,N_2903);
nor U3083 (N_3083,N_2873,N_2826);
and U3084 (N_3084,N_2799,N_2806);
or U3085 (N_3085,N_2833,N_2894);
or U3086 (N_3086,N_2913,N_2803);
xnor U3087 (N_3087,N_2804,N_2784);
and U3088 (N_3088,N_2961,N_2927);
and U3089 (N_3089,N_2816,N_2782);
or U3090 (N_3090,N_2911,N_2787);
or U3091 (N_3091,N_2861,N_2772);
xnor U3092 (N_3092,N_2890,N_2960);
or U3093 (N_3093,N_2916,N_2797);
or U3094 (N_3094,N_2922,N_2774);
nor U3095 (N_3095,N_2891,N_2901);
nor U3096 (N_3096,N_2838,N_2798);
and U3097 (N_3097,N_2914,N_2996);
and U3098 (N_3098,N_2945,N_2835);
and U3099 (N_3099,N_2796,N_2956);
and U3100 (N_3100,N_2813,N_2923);
or U3101 (N_3101,N_2819,N_2751);
nand U3102 (N_3102,N_2859,N_2981);
or U3103 (N_3103,N_2785,N_2762);
and U3104 (N_3104,N_2756,N_2868);
nand U3105 (N_3105,N_2904,N_2970);
nor U3106 (N_3106,N_2980,N_2871);
and U3107 (N_3107,N_2808,N_2986);
or U3108 (N_3108,N_2934,N_2979);
and U3109 (N_3109,N_2827,N_2862);
nor U3110 (N_3110,N_2998,N_2892);
or U3111 (N_3111,N_2775,N_2848);
nand U3112 (N_3112,N_2987,N_2820);
nor U3113 (N_3113,N_2898,N_2836);
nor U3114 (N_3114,N_2899,N_2795);
or U3115 (N_3115,N_2828,N_2846);
and U3116 (N_3116,N_2824,N_2847);
nor U3117 (N_3117,N_2999,N_2955);
and U3118 (N_3118,N_2909,N_2850);
or U3119 (N_3119,N_2884,N_2852);
nand U3120 (N_3120,N_2856,N_2800);
or U3121 (N_3121,N_2908,N_2930);
nor U3122 (N_3122,N_2781,N_2920);
xor U3123 (N_3123,N_2845,N_2995);
and U3124 (N_3124,N_2776,N_2807);
nor U3125 (N_3125,N_2890,N_2845);
and U3126 (N_3126,N_2863,N_2790);
nand U3127 (N_3127,N_2941,N_2774);
nor U3128 (N_3128,N_2820,N_2910);
and U3129 (N_3129,N_2788,N_2817);
and U3130 (N_3130,N_2824,N_2870);
or U3131 (N_3131,N_2805,N_2937);
nor U3132 (N_3132,N_2776,N_2966);
nor U3133 (N_3133,N_2914,N_2757);
nor U3134 (N_3134,N_2927,N_2758);
nor U3135 (N_3135,N_2766,N_2757);
nor U3136 (N_3136,N_2759,N_2875);
nor U3137 (N_3137,N_2849,N_2969);
nand U3138 (N_3138,N_2844,N_2984);
nand U3139 (N_3139,N_2850,N_2863);
nor U3140 (N_3140,N_2953,N_2916);
and U3141 (N_3141,N_2783,N_2957);
and U3142 (N_3142,N_2900,N_2889);
or U3143 (N_3143,N_2792,N_2906);
nor U3144 (N_3144,N_2761,N_2974);
and U3145 (N_3145,N_2944,N_2871);
nor U3146 (N_3146,N_2918,N_2900);
nor U3147 (N_3147,N_2859,N_2924);
nor U3148 (N_3148,N_2795,N_2912);
nand U3149 (N_3149,N_2847,N_2849);
and U3150 (N_3150,N_2808,N_2867);
nand U3151 (N_3151,N_2852,N_2804);
or U3152 (N_3152,N_2880,N_2785);
xnor U3153 (N_3153,N_2948,N_2800);
and U3154 (N_3154,N_2946,N_2760);
and U3155 (N_3155,N_2936,N_2783);
nor U3156 (N_3156,N_2843,N_2800);
and U3157 (N_3157,N_2883,N_2961);
nand U3158 (N_3158,N_2801,N_2900);
or U3159 (N_3159,N_2799,N_2928);
nor U3160 (N_3160,N_2970,N_2924);
or U3161 (N_3161,N_2814,N_2859);
and U3162 (N_3162,N_2855,N_2937);
nor U3163 (N_3163,N_2953,N_2816);
and U3164 (N_3164,N_2767,N_2949);
and U3165 (N_3165,N_2885,N_2816);
nand U3166 (N_3166,N_2770,N_2832);
and U3167 (N_3167,N_2893,N_2986);
or U3168 (N_3168,N_2992,N_2897);
nand U3169 (N_3169,N_2809,N_2753);
or U3170 (N_3170,N_2963,N_2759);
or U3171 (N_3171,N_2794,N_2936);
or U3172 (N_3172,N_2766,N_2970);
xnor U3173 (N_3173,N_2783,N_2982);
nor U3174 (N_3174,N_2903,N_2946);
and U3175 (N_3175,N_2981,N_2769);
nand U3176 (N_3176,N_2807,N_2960);
nor U3177 (N_3177,N_2829,N_2809);
nand U3178 (N_3178,N_2940,N_2790);
or U3179 (N_3179,N_2967,N_2818);
and U3180 (N_3180,N_2889,N_2987);
and U3181 (N_3181,N_2990,N_2994);
and U3182 (N_3182,N_2874,N_2891);
or U3183 (N_3183,N_2970,N_2958);
nor U3184 (N_3184,N_2982,N_2784);
nand U3185 (N_3185,N_2919,N_2853);
nor U3186 (N_3186,N_2785,N_2844);
and U3187 (N_3187,N_2925,N_2936);
and U3188 (N_3188,N_2858,N_2785);
or U3189 (N_3189,N_2787,N_2945);
nand U3190 (N_3190,N_2752,N_2787);
and U3191 (N_3191,N_2964,N_2849);
and U3192 (N_3192,N_2921,N_2773);
nor U3193 (N_3193,N_2751,N_2851);
nand U3194 (N_3194,N_2758,N_2958);
and U3195 (N_3195,N_2798,N_2808);
nand U3196 (N_3196,N_2942,N_2827);
xnor U3197 (N_3197,N_2995,N_2930);
nor U3198 (N_3198,N_2838,N_2845);
or U3199 (N_3199,N_2789,N_2884);
and U3200 (N_3200,N_2793,N_2835);
and U3201 (N_3201,N_2995,N_2993);
nor U3202 (N_3202,N_2881,N_2945);
and U3203 (N_3203,N_2901,N_2988);
or U3204 (N_3204,N_2810,N_2889);
or U3205 (N_3205,N_2902,N_2888);
or U3206 (N_3206,N_2948,N_2993);
and U3207 (N_3207,N_2999,N_2848);
nor U3208 (N_3208,N_2883,N_2956);
or U3209 (N_3209,N_2917,N_2915);
or U3210 (N_3210,N_2873,N_2819);
nor U3211 (N_3211,N_2867,N_2909);
nand U3212 (N_3212,N_2830,N_2905);
or U3213 (N_3213,N_2822,N_2757);
nor U3214 (N_3214,N_2825,N_2877);
nor U3215 (N_3215,N_2865,N_2976);
or U3216 (N_3216,N_2874,N_2780);
and U3217 (N_3217,N_2852,N_2930);
nand U3218 (N_3218,N_2838,N_2981);
nor U3219 (N_3219,N_2865,N_2781);
nand U3220 (N_3220,N_2806,N_2773);
or U3221 (N_3221,N_2950,N_2819);
and U3222 (N_3222,N_2971,N_2957);
and U3223 (N_3223,N_2950,N_2772);
or U3224 (N_3224,N_2885,N_2848);
nor U3225 (N_3225,N_2940,N_2919);
nand U3226 (N_3226,N_2960,N_2985);
nor U3227 (N_3227,N_2776,N_2836);
xnor U3228 (N_3228,N_2973,N_2757);
and U3229 (N_3229,N_2785,N_2923);
nor U3230 (N_3230,N_2876,N_2969);
nor U3231 (N_3231,N_2917,N_2801);
nor U3232 (N_3232,N_2805,N_2778);
xnor U3233 (N_3233,N_2965,N_2791);
nand U3234 (N_3234,N_2975,N_2875);
xor U3235 (N_3235,N_2846,N_2965);
or U3236 (N_3236,N_2812,N_2869);
nor U3237 (N_3237,N_2799,N_2892);
or U3238 (N_3238,N_2782,N_2808);
nand U3239 (N_3239,N_2836,N_2770);
or U3240 (N_3240,N_2895,N_2863);
nand U3241 (N_3241,N_2806,N_2840);
and U3242 (N_3242,N_2836,N_2854);
or U3243 (N_3243,N_2754,N_2995);
or U3244 (N_3244,N_2873,N_2895);
or U3245 (N_3245,N_2940,N_2995);
or U3246 (N_3246,N_2986,N_2960);
nand U3247 (N_3247,N_2940,N_2854);
or U3248 (N_3248,N_2786,N_2904);
nand U3249 (N_3249,N_2993,N_2941);
and U3250 (N_3250,N_3043,N_3130);
nand U3251 (N_3251,N_3092,N_3086);
nand U3252 (N_3252,N_3041,N_3024);
and U3253 (N_3253,N_3172,N_3085);
or U3254 (N_3254,N_3112,N_3010);
nand U3255 (N_3255,N_3117,N_3033);
nand U3256 (N_3256,N_3109,N_3134);
and U3257 (N_3257,N_3071,N_3114);
and U3258 (N_3258,N_3019,N_3018);
nor U3259 (N_3259,N_3188,N_3240);
or U3260 (N_3260,N_3243,N_3137);
and U3261 (N_3261,N_3249,N_3177);
nor U3262 (N_3262,N_3124,N_3186);
or U3263 (N_3263,N_3003,N_3081);
nand U3264 (N_3264,N_3235,N_3139);
and U3265 (N_3265,N_3073,N_3210);
nand U3266 (N_3266,N_3074,N_3170);
nor U3267 (N_3267,N_3077,N_3103);
nor U3268 (N_3268,N_3217,N_3054);
and U3269 (N_3269,N_3023,N_3002);
or U3270 (N_3270,N_3095,N_3191);
nand U3271 (N_3271,N_3102,N_3029);
nor U3272 (N_3272,N_3146,N_3202);
nand U3273 (N_3273,N_3223,N_3218);
nor U3274 (N_3274,N_3066,N_3052);
or U3275 (N_3275,N_3208,N_3006);
and U3276 (N_3276,N_3214,N_3072);
nor U3277 (N_3277,N_3111,N_3198);
nand U3278 (N_3278,N_3174,N_3021);
and U3279 (N_3279,N_3084,N_3205);
and U3280 (N_3280,N_3050,N_3147);
or U3281 (N_3281,N_3157,N_3207);
nand U3282 (N_3282,N_3047,N_3094);
nand U3283 (N_3283,N_3036,N_3068);
nand U3284 (N_3284,N_3244,N_3197);
nor U3285 (N_3285,N_3220,N_3231);
xor U3286 (N_3286,N_3101,N_3224);
nor U3287 (N_3287,N_3125,N_3025);
nor U3288 (N_3288,N_3195,N_3184);
or U3289 (N_3289,N_3027,N_3219);
and U3290 (N_3290,N_3132,N_3065);
and U3291 (N_3291,N_3088,N_3087);
or U3292 (N_3292,N_3190,N_3135);
and U3293 (N_3293,N_3166,N_3230);
or U3294 (N_3294,N_3062,N_3100);
or U3295 (N_3295,N_3180,N_3129);
and U3296 (N_3296,N_3140,N_3200);
or U3297 (N_3297,N_3193,N_3007);
or U3298 (N_3298,N_3000,N_3121);
or U3299 (N_3299,N_3076,N_3167);
or U3300 (N_3300,N_3004,N_3143);
nor U3301 (N_3301,N_3211,N_3136);
nand U3302 (N_3302,N_3171,N_3032);
or U3303 (N_3303,N_3159,N_3001);
nor U3304 (N_3304,N_3040,N_3016);
nand U3305 (N_3305,N_3215,N_3096);
and U3306 (N_3306,N_3082,N_3141);
nor U3307 (N_3307,N_3097,N_3115);
or U3308 (N_3308,N_3080,N_3017);
nand U3309 (N_3309,N_3038,N_3067);
nor U3310 (N_3310,N_3221,N_3022);
nor U3311 (N_3311,N_3090,N_3175);
nor U3312 (N_3312,N_3131,N_3044);
and U3313 (N_3313,N_3160,N_3245);
and U3314 (N_3314,N_3222,N_3206);
nand U3315 (N_3315,N_3151,N_3042);
nor U3316 (N_3316,N_3083,N_3105);
nor U3317 (N_3317,N_3031,N_3149);
nor U3318 (N_3318,N_3216,N_3128);
nand U3319 (N_3319,N_3229,N_3045);
nor U3320 (N_3320,N_3236,N_3113);
nand U3321 (N_3321,N_3213,N_3011);
nand U3322 (N_3322,N_3093,N_3049);
nand U3323 (N_3323,N_3199,N_3148);
and U3324 (N_3324,N_3126,N_3212);
nor U3325 (N_3325,N_3106,N_3058);
nand U3326 (N_3326,N_3056,N_3069);
or U3327 (N_3327,N_3192,N_3183);
and U3328 (N_3328,N_3154,N_3242);
nand U3329 (N_3329,N_3122,N_3150);
nand U3330 (N_3330,N_3178,N_3107);
and U3331 (N_3331,N_3123,N_3039);
and U3332 (N_3332,N_3079,N_3165);
nand U3333 (N_3333,N_3098,N_3089);
nand U3334 (N_3334,N_3187,N_3037);
and U3335 (N_3335,N_3108,N_3034);
or U3336 (N_3336,N_3142,N_3005);
nor U3337 (N_3337,N_3026,N_3013);
and U3338 (N_3338,N_3110,N_3048);
nand U3339 (N_3339,N_3232,N_3008);
nand U3340 (N_3340,N_3091,N_3185);
nand U3341 (N_3341,N_3155,N_3168);
and U3342 (N_3342,N_3133,N_3203);
and U3343 (N_3343,N_3226,N_3099);
and U3344 (N_3344,N_3164,N_3169);
or U3345 (N_3345,N_3173,N_3209);
nor U3346 (N_3346,N_3120,N_3204);
and U3347 (N_3347,N_3233,N_3234);
or U3348 (N_3348,N_3063,N_3248);
nor U3349 (N_3349,N_3035,N_3070);
or U3350 (N_3350,N_3156,N_3162);
nand U3351 (N_3351,N_3051,N_3078);
and U3352 (N_3352,N_3020,N_3158);
xor U3353 (N_3353,N_3237,N_3189);
or U3354 (N_3354,N_3053,N_3012);
and U3355 (N_3355,N_3138,N_3104);
or U3356 (N_3356,N_3241,N_3163);
nor U3357 (N_3357,N_3227,N_3247);
nor U3358 (N_3358,N_3145,N_3118);
nand U3359 (N_3359,N_3060,N_3046);
and U3360 (N_3360,N_3064,N_3055);
xnor U3361 (N_3361,N_3194,N_3119);
and U3362 (N_3362,N_3228,N_3179);
and U3363 (N_3363,N_3061,N_3196);
and U3364 (N_3364,N_3127,N_3161);
and U3365 (N_3365,N_3182,N_3246);
and U3366 (N_3366,N_3009,N_3144);
nand U3367 (N_3367,N_3201,N_3181);
or U3368 (N_3368,N_3028,N_3239);
or U3369 (N_3369,N_3059,N_3176);
nand U3370 (N_3370,N_3030,N_3015);
nand U3371 (N_3371,N_3152,N_3116);
and U3372 (N_3372,N_3238,N_3075);
and U3373 (N_3373,N_3153,N_3225);
and U3374 (N_3374,N_3014,N_3057);
or U3375 (N_3375,N_3181,N_3208);
xnor U3376 (N_3376,N_3132,N_3162);
nor U3377 (N_3377,N_3025,N_3092);
xor U3378 (N_3378,N_3235,N_3067);
or U3379 (N_3379,N_3199,N_3126);
or U3380 (N_3380,N_3020,N_3096);
nor U3381 (N_3381,N_3006,N_3226);
or U3382 (N_3382,N_3012,N_3224);
nor U3383 (N_3383,N_3085,N_3235);
nand U3384 (N_3384,N_3150,N_3083);
nand U3385 (N_3385,N_3039,N_3083);
or U3386 (N_3386,N_3070,N_3132);
and U3387 (N_3387,N_3030,N_3231);
nand U3388 (N_3388,N_3022,N_3045);
and U3389 (N_3389,N_3069,N_3231);
nand U3390 (N_3390,N_3069,N_3052);
nor U3391 (N_3391,N_3162,N_3157);
or U3392 (N_3392,N_3093,N_3153);
nor U3393 (N_3393,N_3147,N_3008);
or U3394 (N_3394,N_3200,N_3234);
and U3395 (N_3395,N_3057,N_3021);
nor U3396 (N_3396,N_3022,N_3142);
nor U3397 (N_3397,N_3033,N_3240);
nor U3398 (N_3398,N_3147,N_3165);
nor U3399 (N_3399,N_3131,N_3099);
nand U3400 (N_3400,N_3105,N_3039);
nand U3401 (N_3401,N_3150,N_3135);
nor U3402 (N_3402,N_3247,N_3114);
or U3403 (N_3403,N_3117,N_3060);
nand U3404 (N_3404,N_3142,N_3163);
or U3405 (N_3405,N_3152,N_3177);
nand U3406 (N_3406,N_3074,N_3041);
nand U3407 (N_3407,N_3003,N_3138);
and U3408 (N_3408,N_3024,N_3028);
or U3409 (N_3409,N_3245,N_3005);
nand U3410 (N_3410,N_3003,N_3012);
and U3411 (N_3411,N_3071,N_3009);
or U3412 (N_3412,N_3117,N_3121);
nor U3413 (N_3413,N_3144,N_3057);
or U3414 (N_3414,N_3239,N_3108);
nor U3415 (N_3415,N_3089,N_3148);
and U3416 (N_3416,N_3080,N_3012);
or U3417 (N_3417,N_3233,N_3049);
nand U3418 (N_3418,N_3032,N_3057);
or U3419 (N_3419,N_3134,N_3249);
nor U3420 (N_3420,N_3245,N_3156);
nand U3421 (N_3421,N_3157,N_3210);
or U3422 (N_3422,N_3059,N_3026);
and U3423 (N_3423,N_3209,N_3178);
nor U3424 (N_3424,N_3209,N_3198);
nand U3425 (N_3425,N_3207,N_3076);
nor U3426 (N_3426,N_3052,N_3005);
or U3427 (N_3427,N_3107,N_3041);
or U3428 (N_3428,N_3131,N_3009);
xor U3429 (N_3429,N_3057,N_3031);
nand U3430 (N_3430,N_3120,N_3119);
and U3431 (N_3431,N_3105,N_3220);
nand U3432 (N_3432,N_3238,N_3112);
and U3433 (N_3433,N_3057,N_3240);
nor U3434 (N_3434,N_3070,N_3228);
and U3435 (N_3435,N_3022,N_3135);
nor U3436 (N_3436,N_3008,N_3033);
nor U3437 (N_3437,N_3034,N_3027);
nor U3438 (N_3438,N_3191,N_3131);
xnor U3439 (N_3439,N_3060,N_3137);
nor U3440 (N_3440,N_3056,N_3123);
or U3441 (N_3441,N_3165,N_3248);
nand U3442 (N_3442,N_3051,N_3010);
nor U3443 (N_3443,N_3082,N_3135);
xor U3444 (N_3444,N_3161,N_3060);
and U3445 (N_3445,N_3040,N_3083);
xor U3446 (N_3446,N_3224,N_3172);
nand U3447 (N_3447,N_3071,N_3175);
and U3448 (N_3448,N_3248,N_3071);
nand U3449 (N_3449,N_3114,N_3099);
nand U3450 (N_3450,N_3173,N_3075);
nand U3451 (N_3451,N_3179,N_3098);
and U3452 (N_3452,N_3063,N_3166);
nand U3453 (N_3453,N_3076,N_3018);
nor U3454 (N_3454,N_3162,N_3239);
and U3455 (N_3455,N_3112,N_3246);
nor U3456 (N_3456,N_3156,N_3136);
nor U3457 (N_3457,N_3146,N_3007);
and U3458 (N_3458,N_3150,N_3004);
or U3459 (N_3459,N_3244,N_3246);
or U3460 (N_3460,N_3049,N_3084);
nand U3461 (N_3461,N_3114,N_3187);
nor U3462 (N_3462,N_3049,N_3173);
nand U3463 (N_3463,N_3113,N_3222);
nor U3464 (N_3464,N_3048,N_3072);
or U3465 (N_3465,N_3139,N_3031);
or U3466 (N_3466,N_3134,N_3086);
or U3467 (N_3467,N_3088,N_3137);
nand U3468 (N_3468,N_3233,N_3030);
or U3469 (N_3469,N_3171,N_3003);
nor U3470 (N_3470,N_3025,N_3224);
and U3471 (N_3471,N_3026,N_3152);
nor U3472 (N_3472,N_3151,N_3103);
and U3473 (N_3473,N_3180,N_3220);
nor U3474 (N_3474,N_3004,N_3081);
nor U3475 (N_3475,N_3211,N_3099);
nor U3476 (N_3476,N_3083,N_3187);
and U3477 (N_3477,N_3042,N_3137);
nand U3478 (N_3478,N_3060,N_3032);
or U3479 (N_3479,N_3138,N_3026);
nor U3480 (N_3480,N_3232,N_3195);
nand U3481 (N_3481,N_3155,N_3002);
or U3482 (N_3482,N_3022,N_3069);
nand U3483 (N_3483,N_3117,N_3091);
nand U3484 (N_3484,N_3063,N_3050);
and U3485 (N_3485,N_3177,N_3104);
nand U3486 (N_3486,N_3042,N_3044);
nand U3487 (N_3487,N_3126,N_3167);
nand U3488 (N_3488,N_3151,N_3143);
and U3489 (N_3489,N_3053,N_3120);
and U3490 (N_3490,N_3005,N_3025);
or U3491 (N_3491,N_3102,N_3197);
or U3492 (N_3492,N_3133,N_3058);
and U3493 (N_3493,N_3091,N_3060);
nor U3494 (N_3494,N_3116,N_3189);
and U3495 (N_3495,N_3228,N_3037);
and U3496 (N_3496,N_3141,N_3207);
nand U3497 (N_3497,N_3208,N_3097);
or U3498 (N_3498,N_3080,N_3112);
and U3499 (N_3499,N_3095,N_3087);
and U3500 (N_3500,N_3335,N_3261);
nor U3501 (N_3501,N_3284,N_3357);
or U3502 (N_3502,N_3394,N_3437);
nand U3503 (N_3503,N_3493,N_3392);
or U3504 (N_3504,N_3298,N_3419);
or U3505 (N_3505,N_3269,N_3359);
or U3506 (N_3506,N_3280,N_3306);
xor U3507 (N_3507,N_3389,N_3473);
nor U3508 (N_3508,N_3301,N_3383);
and U3509 (N_3509,N_3267,N_3339);
nor U3510 (N_3510,N_3421,N_3498);
or U3511 (N_3511,N_3326,N_3397);
and U3512 (N_3512,N_3330,N_3379);
and U3513 (N_3513,N_3313,N_3453);
and U3514 (N_3514,N_3270,N_3444);
nor U3515 (N_3515,N_3406,N_3302);
nor U3516 (N_3516,N_3414,N_3290);
nand U3517 (N_3517,N_3430,N_3368);
nand U3518 (N_3518,N_3338,N_3289);
nand U3519 (N_3519,N_3426,N_3499);
or U3520 (N_3520,N_3467,N_3276);
nor U3521 (N_3521,N_3288,N_3366);
or U3522 (N_3522,N_3360,N_3463);
nand U3523 (N_3523,N_3398,N_3415);
and U3524 (N_3524,N_3312,N_3310);
nor U3525 (N_3525,N_3420,N_3395);
and U3526 (N_3526,N_3412,N_3402);
nor U3527 (N_3527,N_3293,N_3390);
and U3528 (N_3528,N_3454,N_3271);
and U3529 (N_3529,N_3345,N_3303);
and U3530 (N_3530,N_3381,N_3294);
nor U3531 (N_3531,N_3393,N_3364);
and U3532 (N_3532,N_3457,N_3468);
and U3533 (N_3533,N_3332,N_3484);
and U3534 (N_3534,N_3262,N_3275);
or U3535 (N_3535,N_3496,N_3340);
nor U3536 (N_3536,N_3328,N_3418);
or U3537 (N_3537,N_3342,N_3466);
and U3538 (N_3538,N_3321,N_3322);
nand U3539 (N_3539,N_3304,N_3341);
or U3540 (N_3540,N_3449,N_3474);
nor U3541 (N_3541,N_3378,N_3327);
xnor U3542 (N_3542,N_3403,N_3264);
nor U3543 (N_3543,N_3380,N_3459);
or U3544 (N_3544,N_3325,N_3350);
or U3545 (N_3545,N_3282,N_3472);
or U3546 (N_3546,N_3363,N_3433);
and U3547 (N_3547,N_3324,N_3291);
or U3548 (N_3548,N_3361,N_3452);
or U3549 (N_3549,N_3358,N_3408);
or U3550 (N_3550,N_3423,N_3251);
nor U3551 (N_3551,N_3354,N_3385);
nor U3552 (N_3552,N_3460,N_3254);
nand U3553 (N_3553,N_3456,N_3417);
and U3554 (N_3554,N_3431,N_3265);
nor U3555 (N_3555,N_3425,N_3268);
and U3556 (N_3556,N_3266,N_3349);
xnor U3557 (N_3557,N_3300,N_3318);
or U3558 (N_3558,N_3283,N_3387);
and U3559 (N_3559,N_3494,N_3388);
or U3560 (N_3560,N_3477,N_3478);
nand U3561 (N_3561,N_3427,N_3308);
nand U3562 (N_3562,N_3448,N_3292);
nand U3563 (N_3563,N_3485,N_3488);
and U3564 (N_3564,N_3407,N_3458);
and U3565 (N_3565,N_3272,N_3455);
or U3566 (N_3566,N_3344,N_3491);
and U3567 (N_3567,N_3329,N_3447);
nand U3568 (N_3568,N_3495,N_3476);
nand U3569 (N_3569,N_3483,N_3487);
and U3570 (N_3570,N_3400,N_3465);
or U3571 (N_3571,N_3347,N_3497);
and U3572 (N_3572,N_3299,N_3479);
or U3573 (N_3573,N_3286,N_3428);
and U3574 (N_3574,N_3445,N_3295);
and U3575 (N_3575,N_3320,N_3323);
nor U3576 (N_3576,N_3316,N_3376);
and U3577 (N_3577,N_3297,N_3355);
nor U3578 (N_3578,N_3352,N_3274);
nand U3579 (N_3579,N_3482,N_3377);
nand U3580 (N_3580,N_3409,N_3371);
nand U3581 (N_3581,N_3471,N_3351);
and U3582 (N_3582,N_3369,N_3461);
or U3583 (N_3583,N_3470,N_3353);
nor U3584 (N_3584,N_3372,N_3391);
or U3585 (N_3585,N_3384,N_3481);
or U3586 (N_3586,N_3439,N_3416);
nor U3587 (N_3587,N_3442,N_3252);
nor U3588 (N_3588,N_3255,N_3336);
and U3589 (N_3589,N_3489,N_3446);
or U3590 (N_3590,N_3256,N_3260);
nand U3591 (N_3591,N_3438,N_3362);
nor U3592 (N_3592,N_3365,N_3396);
and U3593 (N_3593,N_3374,N_3405);
or U3594 (N_3594,N_3287,N_3404);
and U3595 (N_3595,N_3399,N_3486);
nand U3596 (N_3596,N_3462,N_3337);
or U3597 (N_3597,N_3401,N_3424);
or U3598 (N_3598,N_3434,N_3314);
nor U3599 (N_3599,N_3348,N_3253);
nand U3600 (N_3600,N_3319,N_3281);
nor U3601 (N_3601,N_3250,N_3279);
and U3602 (N_3602,N_3490,N_3305);
or U3603 (N_3603,N_3413,N_3480);
nor U3604 (N_3604,N_3343,N_3296);
nor U3605 (N_3605,N_3333,N_3382);
nand U3606 (N_3606,N_3475,N_3432);
or U3607 (N_3607,N_3307,N_3315);
and U3608 (N_3608,N_3311,N_3410);
and U3609 (N_3609,N_3435,N_3469);
or U3610 (N_3610,N_3492,N_3440);
nor U3611 (N_3611,N_3464,N_3370);
or U3612 (N_3612,N_3429,N_3367);
or U3613 (N_3613,N_3263,N_3277);
nor U3614 (N_3614,N_3373,N_3422);
nand U3615 (N_3615,N_3443,N_3285);
nand U3616 (N_3616,N_3334,N_3411);
or U3617 (N_3617,N_3273,N_3258);
nand U3618 (N_3618,N_3257,N_3451);
or U3619 (N_3619,N_3278,N_3375);
and U3620 (N_3620,N_3386,N_3259);
nor U3621 (N_3621,N_3441,N_3436);
or U3622 (N_3622,N_3317,N_3346);
and U3623 (N_3623,N_3450,N_3331);
or U3624 (N_3624,N_3309,N_3356);
or U3625 (N_3625,N_3322,N_3303);
or U3626 (N_3626,N_3404,N_3441);
nor U3627 (N_3627,N_3439,N_3386);
nor U3628 (N_3628,N_3251,N_3300);
and U3629 (N_3629,N_3276,N_3274);
and U3630 (N_3630,N_3448,N_3424);
nor U3631 (N_3631,N_3443,N_3250);
or U3632 (N_3632,N_3272,N_3454);
nor U3633 (N_3633,N_3475,N_3256);
and U3634 (N_3634,N_3407,N_3499);
or U3635 (N_3635,N_3415,N_3481);
nand U3636 (N_3636,N_3371,N_3378);
and U3637 (N_3637,N_3405,N_3463);
nor U3638 (N_3638,N_3433,N_3396);
xnor U3639 (N_3639,N_3325,N_3431);
and U3640 (N_3640,N_3328,N_3305);
nand U3641 (N_3641,N_3379,N_3443);
and U3642 (N_3642,N_3452,N_3499);
and U3643 (N_3643,N_3398,N_3498);
nor U3644 (N_3644,N_3328,N_3327);
and U3645 (N_3645,N_3326,N_3472);
and U3646 (N_3646,N_3440,N_3344);
or U3647 (N_3647,N_3390,N_3338);
nor U3648 (N_3648,N_3493,N_3354);
nor U3649 (N_3649,N_3449,N_3358);
nand U3650 (N_3650,N_3386,N_3377);
and U3651 (N_3651,N_3404,N_3366);
or U3652 (N_3652,N_3337,N_3376);
nand U3653 (N_3653,N_3452,N_3441);
nor U3654 (N_3654,N_3476,N_3266);
nand U3655 (N_3655,N_3484,N_3317);
or U3656 (N_3656,N_3289,N_3367);
and U3657 (N_3657,N_3270,N_3492);
and U3658 (N_3658,N_3416,N_3322);
nand U3659 (N_3659,N_3463,N_3363);
nor U3660 (N_3660,N_3447,N_3324);
and U3661 (N_3661,N_3446,N_3456);
and U3662 (N_3662,N_3272,N_3452);
and U3663 (N_3663,N_3446,N_3481);
and U3664 (N_3664,N_3398,N_3253);
and U3665 (N_3665,N_3294,N_3458);
and U3666 (N_3666,N_3361,N_3324);
or U3667 (N_3667,N_3278,N_3338);
nor U3668 (N_3668,N_3467,N_3277);
nor U3669 (N_3669,N_3305,N_3326);
nor U3670 (N_3670,N_3416,N_3422);
and U3671 (N_3671,N_3283,N_3299);
or U3672 (N_3672,N_3293,N_3325);
and U3673 (N_3673,N_3397,N_3317);
or U3674 (N_3674,N_3309,N_3445);
or U3675 (N_3675,N_3300,N_3485);
or U3676 (N_3676,N_3425,N_3267);
and U3677 (N_3677,N_3339,N_3357);
nor U3678 (N_3678,N_3359,N_3363);
nand U3679 (N_3679,N_3379,N_3407);
and U3680 (N_3680,N_3319,N_3347);
and U3681 (N_3681,N_3393,N_3437);
nor U3682 (N_3682,N_3366,N_3317);
and U3683 (N_3683,N_3372,N_3272);
nand U3684 (N_3684,N_3267,N_3316);
nor U3685 (N_3685,N_3367,N_3279);
or U3686 (N_3686,N_3377,N_3411);
nor U3687 (N_3687,N_3313,N_3465);
nor U3688 (N_3688,N_3272,N_3426);
or U3689 (N_3689,N_3404,N_3391);
nor U3690 (N_3690,N_3483,N_3321);
or U3691 (N_3691,N_3397,N_3322);
and U3692 (N_3692,N_3451,N_3274);
and U3693 (N_3693,N_3319,N_3289);
nor U3694 (N_3694,N_3429,N_3415);
and U3695 (N_3695,N_3395,N_3306);
or U3696 (N_3696,N_3254,N_3383);
nor U3697 (N_3697,N_3402,N_3420);
nor U3698 (N_3698,N_3429,N_3460);
nor U3699 (N_3699,N_3459,N_3262);
nand U3700 (N_3700,N_3456,N_3309);
and U3701 (N_3701,N_3344,N_3494);
nor U3702 (N_3702,N_3286,N_3451);
nor U3703 (N_3703,N_3455,N_3270);
and U3704 (N_3704,N_3275,N_3424);
nand U3705 (N_3705,N_3317,N_3333);
and U3706 (N_3706,N_3425,N_3470);
nand U3707 (N_3707,N_3497,N_3323);
and U3708 (N_3708,N_3452,N_3268);
nor U3709 (N_3709,N_3293,N_3412);
nand U3710 (N_3710,N_3477,N_3423);
nand U3711 (N_3711,N_3406,N_3288);
nand U3712 (N_3712,N_3334,N_3369);
or U3713 (N_3713,N_3422,N_3465);
nand U3714 (N_3714,N_3425,N_3320);
or U3715 (N_3715,N_3396,N_3264);
nand U3716 (N_3716,N_3302,N_3310);
nand U3717 (N_3717,N_3481,N_3356);
and U3718 (N_3718,N_3463,N_3408);
nand U3719 (N_3719,N_3306,N_3391);
nor U3720 (N_3720,N_3493,N_3328);
nand U3721 (N_3721,N_3322,N_3405);
or U3722 (N_3722,N_3313,N_3309);
and U3723 (N_3723,N_3329,N_3303);
nand U3724 (N_3724,N_3347,N_3458);
or U3725 (N_3725,N_3279,N_3420);
or U3726 (N_3726,N_3451,N_3498);
xnor U3727 (N_3727,N_3447,N_3344);
nor U3728 (N_3728,N_3490,N_3356);
nand U3729 (N_3729,N_3454,N_3262);
nand U3730 (N_3730,N_3326,N_3417);
nor U3731 (N_3731,N_3274,N_3418);
nor U3732 (N_3732,N_3431,N_3440);
or U3733 (N_3733,N_3390,N_3355);
or U3734 (N_3734,N_3282,N_3385);
nand U3735 (N_3735,N_3386,N_3436);
nand U3736 (N_3736,N_3364,N_3422);
nor U3737 (N_3737,N_3405,N_3473);
and U3738 (N_3738,N_3322,N_3341);
nand U3739 (N_3739,N_3496,N_3459);
nand U3740 (N_3740,N_3301,N_3490);
nand U3741 (N_3741,N_3370,N_3413);
and U3742 (N_3742,N_3366,N_3367);
or U3743 (N_3743,N_3390,N_3445);
nand U3744 (N_3744,N_3284,N_3461);
or U3745 (N_3745,N_3465,N_3271);
or U3746 (N_3746,N_3277,N_3426);
or U3747 (N_3747,N_3496,N_3341);
xnor U3748 (N_3748,N_3482,N_3479);
xor U3749 (N_3749,N_3493,N_3443);
nor U3750 (N_3750,N_3676,N_3665);
nand U3751 (N_3751,N_3728,N_3715);
and U3752 (N_3752,N_3587,N_3515);
and U3753 (N_3753,N_3637,N_3577);
and U3754 (N_3754,N_3694,N_3718);
nand U3755 (N_3755,N_3734,N_3615);
and U3756 (N_3756,N_3574,N_3569);
nor U3757 (N_3757,N_3592,N_3525);
nand U3758 (N_3758,N_3705,N_3541);
nor U3759 (N_3759,N_3596,N_3651);
and U3760 (N_3760,N_3554,N_3548);
and U3761 (N_3761,N_3578,N_3723);
nor U3762 (N_3762,N_3649,N_3602);
nand U3763 (N_3763,N_3608,N_3538);
nor U3764 (N_3764,N_3560,N_3601);
or U3765 (N_3765,N_3725,N_3518);
nand U3766 (N_3766,N_3652,N_3612);
nand U3767 (N_3767,N_3675,N_3598);
and U3768 (N_3768,N_3663,N_3542);
nand U3769 (N_3769,N_3567,N_3724);
nor U3770 (N_3770,N_3590,N_3650);
and U3771 (N_3771,N_3661,N_3540);
nand U3772 (N_3772,N_3636,N_3623);
nor U3773 (N_3773,N_3660,N_3735);
xor U3774 (N_3774,N_3581,N_3579);
nor U3775 (N_3775,N_3528,N_3511);
nand U3776 (N_3776,N_3668,N_3603);
nor U3777 (N_3777,N_3563,N_3575);
nor U3778 (N_3778,N_3604,N_3642);
and U3779 (N_3779,N_3533,N_3729);
or U3780 (N_3780,N_3654,N_3509);
or U3781 (N_3781,N_3619,N_3513);
nor U3782 (N_3782,N_3613,N_3512);
nor U3783 (N_3783,N_3564,N_3736);
nand U3784 (N_3784,N_3698,N_3720);
and U3785 (N_3785,N_3672,N_3625);
nand U3786 (N_3786,N_3614,N_3670);
nor U3787 (N_3787,N_3693,N_3529);
nand U3788 (N_3788,N_3551,N_3706);
and U3789 (N_3789,N_3722,N_3659);
or U3790 (N_3790,N_3745,N_3633);
nor U3791 (N_3791,N_3562,N_3582);
or U3792 (N_3792,N_3657,N_3617);
nor U3793 (N_3793,N_3552,N_3621);
nor U3794 (N_3794,N_3643,N_3641);
and U3795 (N_3795,N_3702,N_3710);
nor U3796 (N_3796,N_3532,N_3656);
and U3797 (N_3797,N_3543,N_3520);
or U3798 (N_3798,N_3704,N_3635);
xnor U3799 (N_3799,N_3684,N_3519);
and U3800 (N_3800,N_3558,N_3576);
and U3801 (N_3801,N_3742,N_3658);
nor U3802 (N_3802,N_3687,N_3536);
and U3803 (N_3803,N_3727,N_3610);
and U3804 (N_3804,N_3624,N_3547);
nor U3805 (N_3805,N_3737,N_3546);
xor U3806 (N_3806,N_3644,N_3732);
and U3807 (N_3807,N_3686,N_3648);
nand U3808 (N_3808,N_3726,N_3580);
or U3809 (N_3809,N_3550,N_3516);
and U3810 (N_3810,N_3571,N_3632);
or U3811 (N_3811,N_3561,N_3739);
xnor U3812 (N_3812,N_3688,N_3628);
or U3813 (N_3813,N_3589,N_3749);
or U3814 (N_3814,N_3714,N_3646);
nand U3815 (N_3815,N_3530,N_3701);
and U3816 (N_3816,N_3593,N_3741);
nand U3817 (N_3817,N_3600,N_3647);
nand U3818 (N_3818,N_3591,N_3709);
nand U3819 (N_3819,N_3539,N_3618);
and U3820 (N_3820,N_3692,N_3506);
nand U3821 (N_3821,N_3640,N_3507);
and U3822 (N_3822,N_3522,N_3622);
or U3823 (N_3823,N_3616,N_3504);
and U3824 (N_3824,N_3746,N_3607);
or U3825 (N_3825,N_3743,N_3740);
or U3826 (N_3826,N_3620,N_3671);
nand U3827 (N_3827,N_3664,N_3708);
nor U3828 (N_3828,N_3586,N_3630);
or U3829 (N_3829,N_3677,N_3697);
and U3830 (N_3830,N_3549,N_3583);
and U3831 (N_3831,N_3711,N_3502);
and U3832 (N_3832,N_3700,N_3597);
or U3833 (N_3833,N_3594,N_3611);
or U3834 (N_3834,N_3559,N_3748);
nor U3835 (N_3835,N_3527,N_3713);
nor U3836 (N_3836,N_3521,N_3662);
or U3837 (N_3837,N_3517,N_3501);
and U3838 (N_3838,N_3689,N_3556);
nand U3839 (N_3839,N_3505,N_3629);
nor U3840 (N_3840,N_3712,N_3655);
nor U3841 (N_3841,N_3634,N_3573);
nor U3842 (N_3842,N_3747,N_3609);
or U3843 (N_3843,N_3699,N_3627);
or U3844 (N_3844,N_3557,N_3570);
nor U3845 (N_3845,N_3500,N_3738);
nand U3846 (N_3846,N_3626,N_3673);
and U3847 (N_3847,N_3514,N_3695);
or U3848 (N_3848,N_3669,N_3510);
and U3849 (N_3849,N_3553,N_3674);
nand U3850 (N_3850,N_3680,N_3572);
nor U3851 (N_3851,N_3683,N_3685);
and U3852 (N_3852,N_3719,N_3744);
nand U3853 (N_3853,N_3588,N_3595);
or U3854 (N_3854,N_3733,N_3645);
or U3855 (N_3855,N_3523,N_3696);
and U3856 (N_3856,N_3638,N_3524);
and U3857 (N_3857,N_3566,N_3703);
nor U3858 (N_3858,N_3678,N_3526);
and U3859 (N_3859,N_3605,N_3679);
and U3860 (N_3860,N_3537,N_3717);
or U3861 (N_3861,N_3653,N_3565);
or U3862 (N_3862,N_3730,N_3682);
nor U3863 (N_3863,N_3503,N_3508);
and U3864 (N_3864,N_3534,N_3585);
nor U3865 (N_3865,N_3599,N_3681);
nand U3866 (N_3866,N_3606,N_3631);
nor U3867 (N_3867,N_3544,N_3731);
nor U3868 (N_3868,N_3535,N_3545);
and U3869 (N_3869,N_3690,N_3555);
nand U3870 (N_3870,N_3568,N_3691);
and U3871 (N_3871,N_3531,N_3584);
nand U3872 (N_3872,N_3639,N_3721);
and U3873 (N_3873,N_3667,N_3666);
nand U3874 (N_3874,N_3716,N_3707);
or U3875 (N_3875,N_3582,N_3560);
or U3876 (N_3876,N_3731,N_3617);
or U3877 (N_3877,N_3737,N_3553);
and U3878 (N_3878,N_3705,N_3573);
nor U3879 (N_3879,N_3567,N_3569);
xnor U3880 (N_3880,N_3511,N_3690);
and U3881 (N_3881,N_3552,N_3630);
nor U3882 (N_3882,N_3706,N_3564);
or U3883 (N_3883,N_3687,N_3508);
nor U3884 (N_3884,N_3613,N_3567);
or U3885 (N_3885,N_3541,N_3712);
nand U3886 (N_3886,N_3692,N_3543);
or U3887 (N_3887,N_3674,N_3561);
and U3888 (N_3888,N_3635,N_3686);
nand U3889 (N_3889,N_3589,N_3565);
nor U3890 (N_3890,N_3637,N_3556);
nand U3891 (N_3891,N_3739,N_3686);
xnor U3892 (N_3892,N_3578,N_3645);
nor U3893 (N_3893,N_3532,N_3673);
nor U3894 (N_3894,N_3518,N_3658);
nand U3895 (N_3895,N_3597,N_3650);
nand U3896 (N_3896,N_3528,N_3747);
and U3897 (N_3897,N_3669,N_3529);
nand U3898 (N_3898,N_3701,N_3671);
nor U3899 (N_3899,N_3737,N_3662);
xor U3900 (N_3900,N_3749,N_3534);
nand U3901 (N_3901,N_3728,N_3506);
nand U3902 (N_3902,N_3548,N_3523);
xnor U3903 (N_3903,N_3544,N_3569);
or U3904 (N_3904,N_3527,N_3738);
nand U3905 (N_3905,N_3668,N_3607);
nand U3906 (N_3906,N_3636,N_3549);
and U3907 (N_3907,N_3531,N_3585);
nor U3908 (N_3908,N_3699,N_3530);
and U3909 (N_3909,N_3585,N_3620);
and U3910 (N_3910,N_3640,N_3678);
nand U3911 (N_3911,N_3618,N_3672);
and U3912 (N_3912,N_3587,N_3731);
and U3913 (N_3913,N_3573,N_3597);
and U3914 (N_3914,N_3690,N_3663);
or U3915 (N_3915,N_3609,N_3527);
nor U3916 (N_3916,N_3687,N_3562);
and U3917 (N_3917,N_3712,N_3705);
xnor U3918 (N_3918,N_3562,N_3540);
nor U3919 (N_3919,N_3665,N_3708);
nor U3920 (N_3920,N_3666,N_3525);
nor U3921 (N_3921,N_3524,N_3674);
or U3922 (N_3922,N_3690,N_3660);
xnor U3923 (N_3923,N_3689,N_3522);
nand U3924 (N_3924,N_3611,N_3632);
and U3925 (N_3925,N_3671,N_3583);
or U3926 (N_3926,N_3720,N_3723);
and U3927 (N_3927,N_3501,N_3644);
nor U3928 (N_3928,N_3506,N_3600);
nand U3929 (N_3929,N_3702,N_3704);
and U3930 (N_3930,N_3543,N_3630);
or U3931 (N_3931,N_3579,N_3594);
nand U3932 (N_3932,N_3659,N_3692);
and U3933 (N_3933,N_3637,N_3668);
nor U3934 (N_3934,N_3681,N_3678);
nor U3935 (N_3935,N_3631,N_3700);
and U3936 (N_3936,N_3622,N_3543);
or U3937 (N_3937,N_3544,N_3638);
and U3938 (N_3938,N_3604,N_3510);
xor U3939 (N_3939,N_3520,N_3715);
nor U3940 (N_3940,N_3626,N_3678);
nor U3941 (N_3941,N_3532,N_3516);
nor U3942 (N_3942,N_3614,N_3506);
and U3943 (N_3943,N_3570,N_3549);
or U3944 (N_3944,N_3629,N_3544);
nor U3945 (N_3945,N_3641,N_3506);
and U3946 (N_3946,N_3604,N_3732);
and U3947 (N_3947,N_3543,N_3689);
and U3948 (N_3948,N_3734,N_3521);
and U3949 (N_3949,N_3607,N_3636);
or U3950 (N_3950,N_3627,N_3717);
and U3951 (N_3951,N_3561,N_3732);
nand U3952 (N_3952,N_3691,N_3581);
nor U3953 (N_3953,N_3728,N_3555);
nand U3954 (N_3954,N_3546,N_3610);
and U3955 (N_3955,N_3565,N_3642);
or U3956 (N_3956,N_3516,N_3657);
nand U3957 (N_3957,N_3735,N_3546);
and U3958 (N_3958,N_3502,N_3683);
nor U3959 (N_3959,N_3702,N_3664);
and U3960 (N_3960,N_3510,N_3656);
nand U3961 (N_3961,N_3560,N_3747);
nor U3962 (N_3962,N_3522,N_3697);
and U3963 (N_3963,N_3504,N_3661);
nand U3964 (N_3964,N_3633,N_3677);
nand U3965 (N_3965,N_3637,N_3703);
or U3966 (N_3966,N_3573,N_3666);
or U3967 (N_3967,N_3624,N_3573);
or U3968 (N_3968,N_3728,N_3558);
xnor U3969 (N_3969,N_3549,N_3643);
and U3970 (N_3970,N_3583,N_3521);
nor U3971 (N_3971,N_3536,N_3633);
nand U3972 (N_3972,N_3610,N_3682);
or U3973 (N_3973,N_3655,N_3534);
and U3974 (N_3974,N_3544,N_3652);
or U3975 (N_3975,N_3594,N_3739);
nor U3976 (N_3976,N_3708,N_3631);
and U3977 (N_3977,N_3589,N_3739);
nand U3978 (N_3978,N_3501,N_3679);
nor U3979 (N_3979,N_3679,N_3570);
nor U3980 (N_3980,N_3665,N_3501);
or U3981 (N_3981,N_3625,N_3501);
nand U3982 (N_3982,N_3570,N_3701);
nor U3983 (N_3983,N_3540,N_3665);
nor U3984 (N_3984,N_3747,N_3737);
nor U3985 (N_3985,N_3652,N_3572);
nand U3986 (N_3986,N_3552,N_3745);
nand U3987 (N_3987,N_3508,N_3555);
nand U3988 (N_3988,N_3748,N_3690);
nand U3989 (N_3989,N_3600,N_3574);
and U3990 (N_3990,N_3609,N_3543);
nand U3991 (N_3991,N_3678,N_3550);
and U3992 (N_3992,N_3606,N_3736);
nand U3993 (N_3993,N_3578,N_3673);
nor U3994 (N_3994,N_3579,N_3604);
or U3995 (N_3995,N_3653,N_3729);
or U3996 (N_3996,N_3603,N_3635);
and U3997 (N_3997,N_3531,N_3638);
and U3998 (N_3998,N_3674,N_3527);
nor U3999 (N_3999,N_3657,N_3599);
or U4000 (N_4000,N_3852,N_3867);
nand U4001 (N_4001,N_3836,N_3967);
nor U4002 (N_4002,N_3813,N_3959);
nor U4003 (N_4003,N_3884,N_3982);
and U4004 (N_4004,N_3767,N_3935);
nor U4005 (N_4005,N_3898,N_3974);
nand U4006 (N_4006,N_3986,N_3896);
nand U4007 (N_4007,N_3886,N_3955);
or U4008 (N_4008,N_3766,N_3837);
or U4009 (N_4009,N_3754,N_3811);
nand U4010 (N_4010,N_3944,N_3812);
and U4011 (N_4011,N_3956,N_3933);
nor U4012 (N_4012,N_3819,N_3804);
nor U4013 (N_4013,N_3822,N_3755);
or U4014 (N_4014,N_3885,N_3774);
and U4015 (N_4015,N_3783,N_3840);
nand U4016 (N_4016,N_3798,N_3921);
nand U4017 (N_4017,N_3868,N_3865);
and U4018 (N_4018,N_3940,N_3937);
and U4019 (N_4019,N_3838,N_3781);
and U4020 (N_4020,N_3958,N_3832);
and U4021 (N_4021,N_3963,N_3862);
and U4022 (N_4022,N_3787,N_3759);
nand U4023 (N_4023,N_3768,N_3792);
nand U4024 (N_4024,N_3820,N_3960);
and U4025 (N_4025,N_3823,N_3797);
nand U4026 (N_4026,N_3914,N_3976);
xnor U4027 (N_4027,N_3917,N_3827);
or U4028 (N_4028,N_3999,N_3948);
xor U4029 (N_4029,N_3764,N_3830);
xnor U4030 (N_4030,N_3772,N_3786);
and U4031 (N_4031,N_3841,N_3907);
xor U4032 (N_4032,N_3848,N_3775);
nor U4033 (N_4033,N_3779,N_3995);
or U4034 (N_4034,N_3845,N_3828);
nand U4035 (N_4035,N_3780,N_3784);
nor U4036 (N_4036,N_3824,N_3923);
or U4037 (N_4037,N_3864,N_3901);
or U4038 (N_4038,N_3990,N_3961);
or U4039 (N_4039,N_3928,N_3926);
nand U4040 (N_4040,N_3790,N_3782);
and U4041 (N_4041,N_3954,N_3910);
nor U4042 (N_4042,N_3763,N_3972);
or U4043 (N_4043,N_3752,N_3850);
and U4044 (N_4044,N_3808,N_3874);
nand U4045 (N_4045,N_3984,N_3858);
or U4046 (N_4046,N_3908,N_3891);
nor U4047 (N_4047,N_3873,N_3916);
and U4048 (N_4048,N_3939,N_3849);
or U4049 (N_4049,N_3801,N_3789);
and U4050 (N_4050,N_3796,N_3882);
or U4051 (N_4051,N_3860,N_3800);
nor U4052 (N_4052,N_3943,N_3810);
and U4053 (N_4053,N_3970,N_3969);
nand U4054 (N_4054,N_3871,N_3977);
and U4055 (N_4055,N_3883,N_3994);
nand U4056 (N_4056,N_3757,N_3981);
and U4057 (N_4057,N_3842,N_3900);
nor U4058 (N_4058,N_3869,N_3919);
and U4059 (N_4059,N_3904,N_3911);
nor U4060 (N_4060,N_3794,N_3834);
nand U4061 (N_4061,N_3889,N_3776);
and U4062 (N_4062,N_3906,N_3750);
and U4063 (N_4063,N_3978,N_3816);
or U4064 (N_4064,N_3931,N_3851);
nor U4065 (N_4065,N_3949,N_3902);
or U4066 (N_4066,N_3847,N_3903);
nand U4067 (N_4067,N_3866,N_3778);
nor U4068 (N_4068,N_3785,N_3802);
nand U4069 (N_4069,N_3947,N_3991);
and U4070 (N_4070,N_3980,N_3887);
nor U4071 (N_4071,N_3894,N_3912);
nor U4072 (N_4072,N_3892,N_3859);
or U4073 (N_4073,N_3951,N_3975);
nor U4074 (N_4074,N_3998,N_3756);
or U4075 (N_4075,N_3825,N_3992);
and U4076 (N_4076,N_3761,N_3833);
nand U4077 (N_4077,N_3880,N_3915);
or U4078 (N_4078,N_3815,N_3795);
nand U4079 (N_4079,N_3973,N_3979);
or U4080 (N_4080,N_3888,N_3769);
nand U4081 (N_4081,N_3964,N_3922);
nor U4082 (N_4082,N_3881,N_3762);
nor U4083 (N_4083,N_3872,N_3773);
nor U4084 (N_4084,N_3936,N_3829);
nand U4085 (N_4085,N_3770,N_3993);
or U4086 (N_4086,N_3853,N_3855);
nand U4087 (N_4087,N_3817,N_3826);
and U4088 (N_4088,N_3909,N_3895);
nand U4089 (N_4089,N_3927,N_3953);
or U4090 (N_4090,N_3989,N_3988);
xnor U4091 (N_4091,N_3918,N_3839);
and U4092 (N_4092,N_3925,N_3863);
and U4093 (N_4093,N_3791,N_3777);
or U4094 (N_4094,N_3932,N_3965);
nor U4095 (N_4095,N_3878,N_3983);
xnor U4096 (N_4096,N_3875,N_3805);
nor U4097 (N_4097,N_3893,N_3771);
and U4098 (N_4098,N_3877,N_3843);
and U4099 (N_4099,N_3929,N_3854);
nor U4100 (N_4100,N_3890,N_3920);
or U4101 (N_4101,N_3856,N_3799);
nand U4102 (N_4102,N_3788,N_3861);
nor U4103 (N_4103,N_3818,N_3942);
nor U4104 (N_4104,N_3985,N_3962);
nor U4105 (N_4105,N_3831,N_3879);
nand U4106 (N_4106,N_3941,N_3751);
and U4107 (N_4107,N_3996,N_3803);
nand U4108 (N_4108,N_3899,N_3946);
nor U4109 (N_4109,N_3938,N_3987);
nand U4110 (N_4110,N_3870,N_3930);
nand U4111 (N_4111,N_3876,N_3760);
and U4112 (N_4112,N_3809,N_3758);
nand U4113 (N_4113,N_3934,N_3966);
and U4114 (N_4114,N_3765,N_3950);
or U4115 (N_4115,N_3924,N_3793);
or U4116 (N_4116,N_3945,N_3957);
and U4117 (N_4117,N_3968,N_3807);
nor U4118 (N_4118,N_3971,N_3952);
or U4119 (N_4119,N_3814,N_3997);
or U4120 (N_4120,N_3857,N_3897);
xnor U4121 (N_4121,N_3913,N_3846);
and U4122 (N_4122,N_3806,N_3753);
nand U4123 (N_4123,N_3844,N_3905);
nor U4124 (N_4124,N_3835,N_3821);
nand U4125 (N_4125,N_3912,N_3793);
nand U4126 (N_4126,N_3801,N_3862);
nor U4127 (N_4127,N_3941,N_3784);
nor U4128 (N_4128,N_3793,N_3867);
nor U4129 (N_4129,N_3951,N_3800);
or U4130 (N_4130,N_3852,N_3910);
and U4131 (N_4131,N_3802,N_3979);
nand U4132 (N_4132,N_3831,N_3974);
or U4133 (N_4133,N_3854,N_3799);
and U4134 (N_4134,N_3926,N_3783);
and U4135 (N_4135,N_3922,N_3982);
nand U4136 (N_4136,N_3999,N_3986);
or U4137 (N_4137,N_3850,N_3948);
nor U4138 (N_4138,N_3854,N_3893);
nor U4139 (N_4139,N_3841,N_3903);
nor U4140 (N_4140,N_3840,N_3771);
nor U4141 (N_4141,N_3977,N_3769);
or U4142 (N_4142,N_3839,N_3844);
nand U4143 (N_4143,N_3912,N_3952);
nand U4144 (N_4144,N_3817,N_3782);
nor U4145 (N_4145,N_3820,N_3957);
and U4146 (N_4146,N_3929,N_3806);
and U4147 (N_4147,N_3851,N_3808);
and U4148 (N_4148,N_3895,N_3844);
or U4149 (N_4149,N_3822,N_3900);
nand U4150 (N_4150,N_3871,N_3774);
nor U4151 (N_4151,N_3767,N_3969);
and U4152 (N_4152,N_3991,N_3772);
or U4153 (N_4153,N_3897,N_3780);
nand U4154 (N_4154,N_3892,N_3817);
nor U4155 (N_4155,N_3985,N_3778);
and U4156 (N_4156,N_3899,N_3951);
nand U4157 (N_4157,N_3967,N_3997);
nor U4158 (N_4158,N_3771,N_3978);
nor U4159 (N_4159,N_3877,N_3995);
or U4160 (N_4160,N_3853,N_3844);
and U4161 (N_4161,N_3934,N_3858);
nand U4162 (N_4162,N_3870,N_3938);
or U4163 (N_4163,N_3826,N_3990);
nor U4164 (N_4164,N_3758,N_3904);
and U4165 (N_4165,N_3796,N_3856);
nand U4166 (N_4166,N_3885,N_3876);
nand U4167 (N_4167,N_3782,N_3975);
and U4168 (N_4168,N_3985,N_3909);
nor U4169 (N_4169,N_3875,N_3780);
nor U4170 (N_4170,N_3826,N_3769);
or U4171 (N_4171,N_3934,N_3971);
or U4172 (N_4172,N_3885,N_3952);
xnor U4173 (N_4173,N_3809,N_3820);
or U4174 (N_4174,N_3957,N_3876);
or U4175 (N_4175,N_3952,N_3945);
and U4176 (N_4176,N_3884,N_3986);
nand U4177 (N_4177,N_3825,N_3852);
nor U4178 (N_4178,N_3827,N_3923);
or U4179 (N_4179,N_3784,N_3837);
nor U4180 (N_4180,N_3771,N_3838);
and U4181 (N_4181,N_3912,N_3996);
nand U4182 (N_4182,N_3926,N_3801);
and U4183 (N_4183,N_3939,N_3883);
or U4184 (N_4184,N_3863,N_3983);
nand U4185 (N_4185,N_3899,N_3956);
and U4186 (N_4186,N_3981,N_3921);
nand U4187 (N_4187,N_3926,N_3915);
and U4188 (N_4188,N_3812,N_3972);
and U4189 (N_4189,N_3866,N_3823);
or U4190 (N_4190,N_3929,N_3753);
or U4191 (N_4191,N_3769,N_3770);
and U4192 (N_4192,N_3973,N_3897);
or U4193 (N_4193,N_3997,N_3821);
or U4194 (N_4194,N_3960,N_3941);
and U4195 (N_4195,N_3846,N_3939);
nand U4196 (N_4196,N_3858,N_3961);
nor U4197 (N_4197,N_3799,N_3803);
or U4198 (N_4198,N_3883,N_3820);
and U4199 (N_4199,N_3819,N_3769);
nand U4200 (N_4200,N_3992,N_3894);
or U4201 (N_4201,N_3971,N_3861);
or U4202 (N_4202,N_3931,N_3971);
nand U4203 (N_4203,N_3801,N_3886);
nor U4204 (N_4204,N_3963,N_3902);
and U4205 (N_4205,N_3836,N_3959);
nor U4206 (N_4206,N_3854,N_3875);
and U4207 (N_4207,N_3881,N_3908);
and U4208 (N_4208,N_3803,N_3842);
and U4209 (N_4209,N_3959,N_3789);
and U4210 (N_4210,N_3915,N_3948);
or U4211 (N_4211,N_3984,N_3959);
nand U4212 (N_4212,N_3992,N_3827);
and U4213 (N_4213,N_3943,N_3993);
or U4214 (N_4214,N_3803,N_3773);
nand U4215 (N_4215,N_3997,N_3785);
or U4216 (N_4216,N_3799,N_3996);
or U4217 (N_4217,N_3786,N_3970);
or U4218 (N_4218,N_3761,N_3774);
nand U4219 (N_4219,N_3984,N_3854);
nand U4220 (N_4220,N_3928,N_3921);
nor U4221 (N_4221,N_3994,N_3829);
and U4222 (N_4222,N_3918,N_3795);
or U4223 (N_4223,N_3838,N_3958);
nand U4224 (N_4224,N_3773,N_3774);
or U4225 (N_4225,N_3925,N_3932);
and U4226 (N_4226,N_3950,N_3919);
nor U4227 (N_4227,N_3987,N_3862);
nor U4228 (N_4228,N_3837,N_3986);
nand U4229 (N_4229,N_3860,N_3981);
nand U4230 (N_4230,N_3879,N_3810);
nor U4231 (N_4231,N_3880,N_3800);
nor U4232 (N_4232,N_3751,N_3861);
nand U4233 (N_4233,N_3964,N_3893);
or U4234 (N_4234,N_3835,N_3804);
xor U4235 (N_4235,N_3951,N_3890);
nor U4236 (N_4236,N_3916,N_3871);
and U4237 (N_4237,N_3926,N_3978);
and U4238 (N_4238,N_3861,N_3940);
nor U4239 (N_4239,N_3849,N_3870);
and U4240 (N_4240,N_3960,N_3881);
xor U4241 (N_4241,N_3883,N_3905);
and U4242 (N_4242,N_3751,N_3884);
nand U4243 (N_4243,N_3937,N_3904);
nand U4244 (N_4244,N_3769,N_3911);
and U4245 (N_4245,N_3767,N_3925);
and U4246 (N_4246,N_3858,N_3926);
nor U4247 (N_4247,N_3914,N_3861);
nor U4248 (N_4248,N_3964,N_3783);
nand U4249 (N_4249,N_3895,N_3918);
and U4250 (N_4250,N_4018,N_4130);
nor U4251 (N_4251,N_4029,N_4120);
nor U4252 (N_4252,N_4003,N_4000);
and U4253 (N_4253,N_4241,N_4210);
nor U4254 (N_4254,N_4221,N_4036);
and U4255 (N_4255,N_4246,N_4046);
nand U4256 (N_4256,N_4009,N_4235);
nor U4257 (N_4257,N_4019,N_4111);
nor U4258 (N_4258,N_4214,N_4158);
or U4259 (N_4259,N_4169,N_4022);
or U4260 (N_4260,N_4094,N_4107);
nand U4261 (N_4261,N_4030,N_4016);
or U4262 (N_4262,N_4198,N_4223);
nand U4263 (N_4263,N_4162,N_4099);
nand U4264 (N_4264,N_4207,N_4227);
and U4265 (N_4265,N_4248,N_4050);
or U4266 (N_4266,N_4134,N_4177);
nand U4267 (N_4267,N_4201,N_4231);
nor U4268 (N_4268,N_4102,N_4163);
and U4269 (N_4269,N_4108,N_4017);
nor U4270 (N_4270,N_4185,N_4088);
or U4271 (N_4271,N_4047,N_4125);
nor U4272 (N_4272,N_4247,N_4178);
nor U4273 (N_4273,N_4195,N_4048);
nand U4274 (N_4274,N_4085,N_4187);
nor U4275 (N_4275,N_4174,N_4095);
nor U4276 (N_4276,N_4043,N_4073);
nand U4277 (N_4277,N_4066,N_4014);
nand U4278 (N_4278,N_4194,N_4217);
nand U4279 (N_4279,N_4062,N_4059);
nor U4280 (N_4280,N_4069,N_4166);
and U4281 (N_4281,N_4209,N_4119);
nor U4282 (N_4282,N_4113,N_4087);
and U4283 (N_4283,N_4037,N_4196);
nor U4284 (N_4284,N_4152,N_4151);
nor U4285 (N_4285,N_4086,N_4243);
and U4286 (N_4286,N_4096,N_4123);
nand U4287 (N_4287,N_4191,N_4068);
and U4288 (N_4288,N_4025,N_4127);
nor U4289 (N_4289,N_4135,N_4071);
nor U4290 (N_4290,N_4168,N_4006);
nand U4291 (N_4291,N_4224,N_4184);
and U4292 (N_4292,N_4153,N_4133);
nor U4293 (N_4293,N_4027,N_4218);
nand U4294 (N_4294,N_4203,N_4122);
nand U4295 (N_4295,N_4226,N_4052);
or U4296 (N_4296,N_4034,N_4023);
or U4297 (N_4297,N_4090,N_4117);
and U4298 (N_4298,N_4060,N_4129);
nand U4299 (N_4299,N_4079,N_4212);
and U4300 (N_4300,N_4072,N_4081);
and U4301 (N_4301,N_4232,N_4200);
nor U4302 (N_4302,N_4115,N_4156);
or U4303 (N_4303,N_4026,N_4020);
nor U4304 (N_4304,N_4054,N_4067);
or U4305 (N_4305,N_4197,N_4057);
or U4306 (N_4306,N_4128,N_4244);
or U4307 (N_4307,N_4164,N_4161);
nand U4308 (N_4308,N_4055,N_4121);
or U4309 (N_4309,N_4202,N_4249);
nand U4310 (N_4310,N_4045,N_4171);
nand U4311 (N_4311,N_4091,N_4189);
or U4312 (N_4312,N_4101,N_4175);
and U4313 (N_4313,N_4064,N_4065);
and U4314 (N_4314,N_4206,N_4109);
nand U4315 (N_4315,N_4167,N_4076);
and U4316 (N_4316,N_4005,N_4082);
nor U4317 (N_4317,N_4242,N_4222);
or U4318 (N_4318,N_4116,N_4042);
and U4319 (N_4319,N_4155,N_4228);
nand U4320 (N_4320,N_4002,N_4110);
and U4321 (N_4321,N_4051,N_4040);
nor U4322 (N_4322,N_4233,N_4032);
nor U4323 (N_4323,N_4035,N_4229);
and U4324 (N_4324,N_4139,N_4031);
or U4325 (N_4325,N_4058,N_4092);
and U4326 (N_4326,N_4104,N_4093);
or U4327 (N_4327,N_4188,N_4216);
xnor U4328 (N_4328,N_4183,N_4103);
or U4329 (N_4329,N_4186,N_4080);
and U4330 (N_4330,N_4049,N_4159);
nand U4331 (N_4331,N_4170,N_4001);
and U4332 (N_4332,N_4074,N_4213);
or U4333 (N_4333,N_4225,N_4124);
and U4334 (N_4334,N_4230,N_4148);
nor U4335 (N_4335,N_4220,N_4179);
nor U4336 (N_4336,N_4078,N_4041);
nor U4337 (N_4337,N_4118,N_4089);
nor U4338 (N_4338,N_4144,N_4245);
or U4339 (N_4339,N_4138,N_4160);
nor U4340 (N_4340,N_4021,N_4176);
nor U4341 (N_4341,N_4199,N_4114);
nor U4342 (N_4342,N_4204,N_4173);
nor U4343 (N_4343,N_4208,N_4237);
nand U4344 (N_4344,N_4236,N_4147);
and U4345 (N_4345,N_4182,N_4097);
and U4346 (N_4346,N_4075,N_4239);
and U4347 (N_4347,N_4011,N_4146);
nand U4348 (N_4348,N_4140,N_4149);
nand U4349 (N_4349,N_4083,N_4056);
or U4350 (N_4350,N_4131,N_4157);
nor U4351 (N_4351,N_4033,N_4077);
or U4352 (N_4352,N_4063,N_4126);
nand U4353 (N_4353,N_4215,N_4013);
and U4354 (N_4354,N_4007,N_4172);
xor U4355 (N_4355,N_4238,N_4098);
and U4356 (N_4356,N_4240,N_4137);
and U4357 (N_4357,N_4105,N_4061);
and U4358 (N_4358,N_4136,N_4015);
nor U4359 (N_4359,N_4004,N_4012);
or U4360 (N_4360,N_4154,N_4044);
and U4361 (N_4361,N_4180,N_4010);
or U4362 (N_4362,N_4211,N_4028);
nand U4363 (N_4363,N_4132,N_4234);
or U4364 (N_4364,N_4150,N_4143);
nand U4365 (N_4365,N_4084,N_4145);
or U4366 (N_4366,N_4039,N_4100);
and U4367 (N_4367,N_4219,N_4142);
or U4368 (N_4368,N_4070,N_4181);
and U4369 (N_4369,N_4112,N_4008);
or U4370 (N_4370,N_4141,N_4038);
nor U4371 (N_4371,N_4205,N_4106);
nor U4372 (N_4372,N_4024,N_4165);
or U4373 (N_4373,N_4193,N_4190);
nor U4374 (N_4374,N_4192,N_4053);
nor U4375 (N_4375,N_4060,N_4210);
nor U4376 (N_4376,N_4193,N_4002);
or U4377 (N_4377,N_4230,N_4005);
nand U4378 (N_4378,N_4113,N_4111);
or U4379 (N_4379,N_4072,N_4164);
and U4380 (N_4380,N_4070,N_4101);
or U4381 (N_4381,N_4216,N_4206);
nor U4382 (N_4382,N_4196,N_4053);
or U4383 (N_4383,N_4127,N_4140);
xor U4384 (N_4384,N_4249,N_4036);
or U4385 (N_4385,N_4161,N_4029);
and U4386 (N_4386,N_4191,N_4224);
or U4387 (N_4387,N_4198,N_4029);
and U4388 (N_4388,N_4179,N_4180);
nand U4389 (N_4389,N_4091,N_4000);
nor U4390 (N_4390,N_4215,N_4202);
nor U4391 (N_4391,N_4226,N_4100);
or U4392 (N_4392,N_4185,N_4122);
and U4393 (N_4393,N_4195,N_4161);
xnor U4394 (N_4394,N_4027,N_4185);
or U4395 (N_4395,N_4151,N_4127);
nor U4396 (N_4396,N_4196,N_4135);
nor U4397 (N_4397,N_4106,N_4068);
nand U4398 (N_4398,N_4089,N_4005);
and U4399 (N_4399,N_4099,N_4038);
nor U4400 (N_4400,N_4143,N_4205);
and U4401 (N_4401,N_4218,N_4052);
xor U4402 (N_4402,N_4003,N_4085);
or U4403 (N_4403,N_4128,N_4042);
nor U4404 (N_4404,N_4108,N_4112);
or U4405 (N_4405,N_4045,N_4000);
nand U4406 (N_4406,N_4096,N_4074);
nor U4407 (N_4407,N_4043,N_4107);
xor U4408 (N_4408,N_4243,N_4209);
or U4409 (N_4409,N_4162,N_4072);
nand U4410 (N_4410,N_4144,N_4042);
nor U4411 (N_4411,N_4090,N_4213);
or U4412 (N_4412,N_4064,N_4234);
nand U4413 (N_4413,N_4238,N_4207);
nor U4414 (N_4414,N_4012,N_4048);
or U4415 (N_4415,N_4120,N_4181);
and U4416 (N_4416,N_4204,N_4162);
nand U4417 (N_4417,N_4163,N_4143);
nand U4418 (N_4418,N_4200,N_4149);
nand U4419 (N_4419,N_4027,N_4235);
or U4420 (N_4420,N_4146,N_4202);
nand U4421 (N_4421,N_4068,N_4110);
or U4422 (N_4422,N_4245,N_4090);
nand U4423 (N_4423,N_4047,N_4121);
nor U4424 (N_4424,N_4000,N_4050);
or U4425 (N_4425,N_4185,N_4061);
nand U4426 (N_4426,N_4243,N_4239);
and U4427 (N_4427,N_4106,N_4098);
nor U4428 (N_4428,N_4027,N_4070);
or U4429 (N_4429,N_4243,N_4025);
and U4430 (N_4430,N_4164,N_4079);
and U4431 (N_4431,N_4130,N_4001);
and U4432 (N_4432,N_4229,N_4093);
or U4433 (N_4433,N_4078,N_4114);
nor U4434 (N_4434,N_4218,N_4091);
nor U4435 (N_4435,N_4145,N_4130);
or U4436 (N_4436,N_4051,N_4125);
or U4437 (N_4437,N_4073,N_4150);
nand U4438 (N_4438,N_4043,N_4103);
nor U4439 (N_4439,N_4144,N_4208);
nand U4440 (N_4440,N_4074,N_4056);
and U4441 (N_4441,N_4119,N_4221);
nor U4442 (N_4442,N_4205,N_4021);
or U4443 (N_4443,N_4125,N_4142);
or U4444 (N_4444,N_4157,N_4217);
nand U4445 (N_4445,N_4159,N_4154);
and U4446 (N_4446,N_4120,N_4040);
or U4447 (N_4447,N_4083,N_4066);
and U4448 (N_4448,N_4094,N_4057);
and U4449 (N_4449,N_4079,N_4066);
or U4450 (N_4450,N_4047,N_4040);
nor U4451 (N_4451,N_4130,N_4135);
nand U4452 (N_4452,N_4109,N_4026);
or U4453 (N_4453,N_4239,N_4100);
or U4454 (N_4454,N_4110,N_4209);
or U4455 (N_4455,N_4116,N_4124);
or U4456 (N_4456,N_4227,N_4033);
nor U4457 (N_4457,N_4207,N_4193);
nand U4458 (N_4458,N_4063,N_4093);
nor U4459 (N_4459,N_4201,N_4230);
nand U4460 (N_4460,N_4209,N_4039);
or U4461 (N_4461,N_4098,N_4012);
and U4462 (N_4462,N_4189,N_4007);
nor U4463 (N_4463,N_4132,N_4201);
or U4464 (N_4464,N_4085,N_4102);
or U4465 (N_4465,N_4171,N_4215);
nand U4466 (N_4466,N_4238,N_4239);
nand U4467 (N_4467,N_4175,N_4119);
nor U4468 (N_4468,N_4186,N_4015);
nand U4469 (N_4469,N_4130,N_4050);
or U4470 (N_4470,N_4245,N_4009);
and U4471 (N_4471,N_4003,N_4228);
and U4472 (N_4472,N_4000,N_4196);
or U4473 (N_4473,N_4095,N_4144);
and U4474 (N_4474,N_4190,N_4161);
nand U4475 (N_4475,N_4197,N_4021);
nand U4476 (N_4476,N_4182,N_4158);
and U4477 (N_4477,N_4036,N_4147);
and U4478 (N_4478,N_4130,N_4141);
and U4479 (N_4479,N_4212,N_4056);
nor U4480 (N_4480,N_4112,N_4229);
nand U4481 (N_4481,N_4211,N_4128);
and U4482 (N_4482,N_4176,N_4108);
nor U4483 (N_4483,N_4243,N_4249);
nor U4484 (N_4484,N_4052,N_4205);
or U4485 (N_4485,N_4136,N_4028);
nand U4486 (N_4486,N_4169,N_4184);
nand U4487 (N_4487,N_4070,N_4151);
and U4488 (N_4488,N_4249,N_4205);
xnor U4489 (N_4489,N_4007,N_4195);
nor U4490 (N_4490,N_4173,N_4044);
nor U4491 (N_4491,N_4181,N_4199);
or U4492 (N_4492,N_4004,N_4220);
nor U4493 (N_4493,N_4162,N_4226);
or U4494 (N_4494,N_4027,N_4097);
or U4495 (N_4495,N_4084,N_4130);
nor U4496 (N_4496,N_4233,N_4101);
nor U4497 (N_4497,N_4249,N_4143);
nand U4498 (N_4498,N_4075,N_4110);
or U4499 (N_4499,N_4025,N_4092);
or U4500 (N_4500,N_4267,N_4388);
or U4501 (N_4501,N_4392,N_4461);
or U4502 (N_4502,N_4362,N_4473);
nor U4503 (N_4503,N_4291,N_4372);
and U4504 (N_4504,N_4403,N_4444);
and U4505 (N_4505,N_4465,N_4307);
nand U4506 (N_4506,N_4463,N_4471);
nor U4507 (N_4507,N_4357,N_4278);
nor U4508 (N_4508,N_4319,N_4289);
or U4509 (N_4509,N_4412,N_4353);
or U4510 (N_4510,N_4356,N_4429);
or U4511 (N_4511,N_4468,N_4343);
or U4512 (N_4512,N_4269,N_4454);
nand U4513 (N_4513,N_4433,N_4294);
nand U4514 (N_4514,N_4358,N_4474);
nand U4515 (N_4515,N_4333,N_4484);
nor U4516 (N_4516,N_4308,N_4446);
and U4517 (N_4517,N_4327,N_4389);
and U4518 (N_4518,N_4469,N_4300);
nor U4519 (N_4519,N_4281,N_4260);
nand U4520 (N_4520,N_4415,N_4424);
or U4521 (N_4521,N_4251,N_4445);
nor U4522 (N_4522,N_4489,N_4328);
nand U4523 (N_4523,N_4317,N_4293);
and U4524 (N_4524,N_4441,N_4414);
nand U4525 (N_4525,N_4304,N_4273);
and U4526 (N_4526,N_4338,N_4364);
nand U4527 (N_4527,N_4398,N_4282);
or U4528 (N_4528,N_4418,N_4452);
and U4529 (N_4529,N_4383,N_4368);
and U4530 (N_4530,N_4386,N_4494);
and U4531 (N_4531,N_4331,N_4453);
and U4532 (N_4532,N_4262,N_4394);
xor U4533 (N_4533,N_4421,N_4384);
and U4534 (N_4534,N_4395,N_4376);
or U4535 (N_4535,N_4400,N_4408);
or U4536 (N_4536,N_4464,N_4451);
nand U4537 (N_4537,N_4252,N_4296);
nand U4538 (N_4538,N_4265,N_4298);
nand U4539 (N_4539,N_4332,N_4431);
or U4540 (N_4540,N_4275,N_4306);
nor U4541 (N_4541,N_4344,N_4315);
nand U4542 (N_4542,N_4261,N_4342);
or U4543 (N_4543,N_4310,N_4277);
and U4544 (N_4544,N_4409,N_4425);
or U4545 (N_4545,N_4360,N_4348);
or U4546 (N_4546,N_4435,N_4434);
and U4547 (N_4547,N_4486,N_4416);
and U4548 (N_4548,N_4462,N_4438);
or U4549 (N_4549,N_4391,N_4426);
nor U4550 (N_4550,N_4407,N_4318);
xor U4551 (N_4551,N_4349,N_4259);
nand U4552 (N_4552,N_4363,N_4255);
and U4553 (N_4553,N_4288,N_4498);
nand U4554 (N_4554,N_4427,N_4459);
or U4555 (N_4555,N_4345,N_4487);
nand U4556 (N_4556,N_4413,N_4351);
nor U4557 (N_4557,N_4377,N_4287);
or U4558 (N_4558,N_4271,N_4479);
or U4559 (N_4559,N_4258,N_4477);
nand U4560 (N_4560,N_4305,N_4417);
or U4561 (N_4561,N_4430,N_4390);
and U4562 (N_4562,N_4264,N_4483);
nand U4563 (N_4563,N_4490,N_4420);
nor U4564 (N_4564,N_4436,N_4457);
nand U4565 (N_4565,N_4257,N_4485);
and U4566 (N_4566,N_4268,N_4439);
nand U4567 (N_4567,N_4361,N_4374);
and U4568 (N_4568,N_4292,N_4455);
nand U4569 (N_4569,N_4385,N_4402);
xor U4570 (N_4570,N_4456,N_4303);
nand U4571 (N_4571,N_4380,N_4330);
nand U4572 (N_4572,N_4411,N_4309);
and U4573 (N_4573,N_4340,N_4316);
or U4574 (N_4574,N_4354,N_4443);
or U4575 (N_4575,N_4382,N_4397);
nor U4576 (N_4576,N_4285,N_4396);
or U4577 (N_4577,N_4495,N_4335);
nand U4578 (N_4578,N_4336,N_4373);
nand U4579 (N_4579,N_4410,N_4447);
nor U4580 (N_4580,N_4312,N_4337);
nand U4581 (N_4581,N_4476,N_4405);
nor U4582 (N_4582,N_4379,N_4286);
nor U4583 (N_4583,N_4346,N_4284);
nand U4584 (N_4584,N_4470,N_4324);
xnor U4585 (N_4585,N_4279,N_4272);
or U4586 (N_4586,N_4266,N_4321);
nand U4587 (N_4587,N_4352,N_4491);
nand U4588 (N_4588,N_4320,N_4263);
and U4589 (N_4589,N_4442,N_4322);
or U4590 (N_4590,N_4297,N_4256);
nor U4591 (N_4591,N_4460,N_4314);
or U4592 (N_4592,N_4499,N_4301);
and U4593 (N_4593,N_4428,N_4365);
nand U4594 (N_4594,N_4448,N_4437);
or U4595 (N_4595,N_4270,N_4472);
and U4596 (N_4596,N_4381,N_4422);
nor U4597 (N_4597,N_4493,N_4401);
and U4598 (N_4598,N_4299,N_4488);
xnor U4599 (N_4599,N_4481,N_4480);
or U4600 (N_4600,N_4478,N_4404);
or U4601 (N_4601,N_4355,N_4334);
or U4602 (N_4602,N_4250,N_4496);
nand U4603 (N_4603,N_4466,N_4366);
or U4604 (N_4604,N_4450,N_4311);
and U4605 (N_4605,N_4387,N_4283);
nand U4606 (N_4606,N_4406,N_4329);
or U4607 (N_4607,N_4325,N_4370);
nand U4608 (N_4608,N_4313,N_4359);
or U4609 (N_4609,N_4399,N_4339);
xor U4610 (N_4610,N_4253,N_4378);
nor U4611 (N_4611,N_4393,N_4280);
nand U4612 (N_4612,N_4449,N_4350);
nor U4613 (N_4613,N_4467,N_4367);
or U4614 (N_4614,N_4347,N_4274);
or U4615 (N_4615,N_4369,N_4276);
and U4616 (N_4616,N_4432,N_4290);
and U4617 (N_4617,N_4371,N_4492);
nor U4618 (N_4618,N_4475,N_4323);
and U4619 (N_4619,N_4302,N_4458);
nor U4620 (N_4620,N_4326,N_4423);
and U4621 (N_4621,N_4482,N_4295);
and U4622 (N_4622,N_4254,N_4497);
nor U4623 (N_4623,N_4375,N_4419);
or U4624 (N_4624,N_4341,N_4440);
nand U4625 (N_4625,N_4301,N_4252);
nor U4626 (N_4626,N_4467,N_4426);
nand U4627 (N_4627,N_4395,N_4444);
nor U4628 (N_4628,N_4262,N_4327);
nand U4629 (N_4629,N_4303,N_4250);
and U4630 (N_4630,N_4431,N_4256);
nand U4631 (N_4631,N_4432,N_4433);
nand U4632 (N_4632,N_4321,N_4416);
and U4633 (N_4633,N_4478,N_4451);
nor U4634 (N_4634,N_4252,N_4255);
nor U4635 (N_4635,N_4278,N_4258);
or U4636 (N_4636,N_4487,N_4335);
and U4637 (N_4637,N_4375,N_4355);
nand U4638 (N_4638,N_4253,N_4267);
or U4639 (N_4639,N_4455,N_4268);
nor U4640 (N_4640,N_4465,N_4254);
nand U4641 (N_4641,N_4365,N_4484);
nand U4642 (N_4642,N_4401,N_4442);
and U4643 (N_4643,N_4268,N_4491);
nand U4644 (N_4644,N_4341,N_4337);
and U4645 (N_4645,N_4384,N_4396);
nand U4646 (N_4646,N_4390,N_4358);
or U4647 (N_4647,N_4333,N_4401);
nand U4648 (N_4648,N_4252,N_4433);
nand U4649 (N_4649,N_4389,N_4363);
or U4650 (N_4650,N_4367,N_4327);
or U4651 (N_4651,N_4279,N_4474);
nand U4652 (N_4652,N_4365,N_4444);
nand U4653 (N_4653,N_4373,N_4460);
or U4654 (N_4654,N_4363,N_4485);
nand U4655 (N_4655,N_4285,N_4474);
or U4656 (N_4656,N_4276,N_4273);
nand U4657 (N_4657,N_4411,N_4393);
or U4658 (N_4658,N_4468,N_4480);
nand U4659 (N_4659,N_4255,N_4250);
nand U4660 (N_4660,N_4453,N_4444);
nand U4661 (N_4661,N_4497,N_4345);
nor U4662 (N_4662,N_4259,N_4384);
and U4663 (N_4663,N_4406,N_4398);
and U4664 (N_4664,N_4280,N_4344);
and U4665 (N_4665,N_4487,N_4492);
nand U4666 (N_4666,N_4440,N_4321);
nor U4667 (N_4667,N_4408,N_4495);
or U4668 (N_4668,N_4330,N_4468);
or U4669 (N_4669,N_4316,N_4480);
nand U4670 (N_4670,N_4315,N_4350);
and U4671 (N_4671,N_4444,N_4410);
nand U4672 (N_4672,N_4378,N_4368);
or U4673 (N_4673,N_4271,N_4270);
nand U4674 (N_4674,N_4465,N_4287);
or U4675 (N_4675,N_4318,N_4452);
nor U4676 (N_4676,N_4394,N_4407);
and U4677 (N_4677,N_4264,N_4468);
or U4678 (N_4678,N_4491,N_4478);
and U4679 (N_4679,N_4383,N_4492);
nand U4680 (N_4680,N_4462,N_4307);
nand U4681 (N_4681,N_4405,N_4338);
nor U4682 (N_4682,N_4395,N_4272);
or U4683 (N_4683,N_4326,N_4340);
or U4684 (N_4684,N_4444,N_4303);
nor U4685 (N_4685,N_4316,N_4464);
and U4686 (N_4686,N_4451,N_4421);
or U4687 (N_4687,N_4320,N_4492);
nor U4688 (N_4688,N_4408,N_4284);
or U4689 (N_4689,N_4328,N_4432);
nand U4690 (N_4690,N_4284,N_4470);
and U4691 (N_4691,N_4278,N_4337);
and U4692 (N_4692,N_4284,N_4388);
nor U4693 (N_4693,N_4283,N_4498);
or U4694 (N_4694,N_4365,N_4269);
or U4695 (N_4695,N_4468,N_4440);
and U4696 (N_4696,N_4331,N_4462);
or U4697 (N_4697,N_4434,N_4471);
or U4698 (N_4698,N_4290,N_4435);
and U4699 (N_4699,N_4382,N_4417);
nor U4700 (N_4700,N_4258,N_4471);
nand U4701 (N_4701,N_4499,N_4496);
or U4702 (N_4702,N_4361,N_4426);
or U4703 (N_4703,N_4369,N_4368);
and U4704 (N_4704,N_4439,N_4259);
nor U4705 (N_4705,N_4409,N_4450);
or U4706 (N_4706,N_4399,N_4431);
or U4707 (N_4707,N_4398,N_4474);
and U4708 (N_4708,N_4496,N_4467);
nand U4709 (N_4709,N_4448,N_4257);
and U4710 (N_4710,N_4313,N_4413);
and U4711 (N_4711,N_4433,N_4347);
nor U4712 (N_4712,N_4486,N_4488);
and U4713 (N_4713,N_4431,N_4261);
nor U4714 (N_4714,N_4358,N_4298);
nand U4715 (N_4715,N_4320,N_4479);
nand U4716 (N_4716,N_4368,N_4275);
and U4717 (N_4717,N_4359,N_4411);
nor U4718 (N_4718,N_4436,N_4412);
nand U4719 (N_4719,N_4467,N_4292);
or U4720 (N_4720,N_4448,N_4254);
nor U4721 (N_4721,N_4256,N_4266);
and U4722 (N_4722,N_4414,N_4346);
nor U4723 (N_4723,N_4490,N_4397);
xor U4724 (N_4724,N_4393,N_4406);
nand U4725 (N_4725,N_4288,N_4343);
nor U4726 (N_4726,N_4479,N_4420);
or U4727 (N_4727,N_4338,N_4377);
or U4728 (N_4728,N_4362,N_4352);
and U4729 (N_4729,N_4344,N_4329);
and U4730 (N_4730,N_4327,N_4282);
or U4731 (N_4731,N_4310,N_4498);
nand U4732 (N_4732,N_4265,N_4438);
nor U4733 (N_4733,N_4270,N_4498);
nor U4734 (N_4734,N_4483,N_4419);
and U4735 (N_4735,N_4333,N_4399);
and U4736 (N_4736,N_4282,N_4311);
nor U4737 (N_4737,N_4480,N_4428);
or U4738 (N_4738,N_4484,N_4274);
xor U4739 (N_4739,N_4264,N_4497);
or U4740 (N_4740,N_4337,N_4457);
and U4741 (N_4741,N_4476,N_4251);
nand U4742 (N_4742,N_4469,N_4449);
or U4743 (N_4743,N_4404,N_4455);
or U4744 (N_4744,N_4420,N_4473);
or U4745 (N_4745,N_4489,N_4322);
nor U4746 (N_4746,N_4414,N_4324);
nand U4747 (N_4747,N_4265,N_4397);
nor U4748 (N_4748,N_4302,N_4326);
or U4749 (N_4749,N_4346,N_4366);
or U4750 (N_4750,N_4700,N_4540);
nor U4751 (N_4751,N_4592,N_4695);
nor U4752 (N_4752,N_4690,N_4623);
nor U4753 (N_4753,N_4671,N_4645);
and U4754 (N_4754,N_4585,N_4688);
nor U4755 (N_4755,N_4720,N_4500);
xnor U4756 (N_4756,N_4638,N_4524);
or U4757 (N_4757,N_4625,N_4566);
or U4758 (N_4758,N_4632,N_4675);
and U4759 (N_4759,N_4655,N_4532);
nor U4760 (N_4760,N_4610,N_4571);
and U4761 (N_4761,N_4712,N_4670);
nand U4762 (N_4762,N_4740,N_4711);
and U4763 (N_4763,N_4698,N_4515);
nand U4764 (N_4764,N_4564,N_4741);
nand U4765 (N_4765,N_4531,N_4680);
nand U4766 (N_4766,N_4665,N_4516);
nor U4767 (N_4767,N_4646,N_4501);
and U4768 (N_4768,N_4683,N_4565);
nand U4769 (N_4769,N_4710,N_4613);
and U4770 (N_4770,N_4668,N_4512);
or U4771 (N_4771,N_4550,N_4744);
nand U4772 (N_4772,N_4560,N_4651);
xor U4773 (N_4773,N_4616,N_4597);
or U4774 (N_4774,N_4731,N_4563);
nor U4775 (N_4775,N_4621,N_4510);
or U4776 (N_4776,N_4725,N_4647);
and U4777 (N_4777,N_4745,N_4611);
nand U4778 (N_4778,N_4533,N_4549);
or U4779 (N_4779,N_4539,N_4528);
or U4780 (N_4780,N_4547,N_4506);
or U4781 (N_4781,N_4575,N_4691);
nand U4782 (N_4782,N_4584,N_4591);
nand U4783 (N_4783,N_4618,N_4535);
nand U4784 (N_4784,N_4583,N_4617);
nand U4785 (N_4785,N_4749,N_4570);
or U4786 (N_4786,N_4538,N_4518);
and U4787 (N_4787,N_4542,N_4608);
and U4788 (N_4788,N_4743,N_4713);
nand U4789 (N_4789,N_4662,N_4544);
or U4790 (N_4790,N_4703,N_4656);
and U4791 (N_4791,N_4652,N_4529);
or U4792 (N_4792,N_4619,N_4735);
or U4793 (N_4793,N_4513,N_4622);
and U4794 (N_4794,N_4676,N_4636);
or U4795 (N_4795,N_4525,N_4577);
or U4796 (N_4796,N_4555,N_4620);
nor U4797 (N_4797,N_4567,N_4643);
and U4798 (N_4798,N_4686,N_4728);
or U4799 (N_4799,N_4558,N_4521);
or U4800 (N_4800,N_4705,N_4747);
nand U4801 (N_4801,N_4586,N_4718);
nor U4802 (N_4802,N_4504,N_4677);
nor U4803 (N_4803,N_4574,N_4708);
and U4804 (N_4804,N_4669,N_4733);
nand U4805 (N_4805,N_4674,N_4508);
nor U4806 (N_4806,N_4736,N_4590);
or U4807 (N_4807,N_4634,N_4603);
nor U4808 (N_4808,N_4694,N_4534);
or U4809 (N_4809,N_4522,N_4629);
or U4810 (N_4810,N_4523,N_4598);
nand U4811 (N_4811,N_4648,N_4687);
and U4812 (N_4812,N_4554,N_4546);
and U4813 (N_4813,N_4738,N_4601);
and U4814 (N_4814,N_4511,N_4660);
and U4815 (N_4815,N_4596,N_4692);
and U4816 (N_4816,N_4702,N_4509);
or U4817 (N_4817,N_4579,N_4721);
and U4818 (N_4818,N_4657,N_4658);
or U4819 (N_4819,N_4639,N_4595);
and U4820 (N_4820,N_4576,N_4562);
nor U4821 (N_4821,N_4704,N_4607);
or U4822 (N_4822,N_4707,N_4605);
and U4823 (N_4823,N_4719,N_4734);
nand U4824 (N_4824,N_4682,N_4678);
or U4825 (N_4825,N_4673,N_4502);
nand U4826 (N_4826,N_4653,N_4514);
or U4827 (N_4827,N_4701,N_4724);
nor U4828 (N_4828,N_4589,N_4527);
nand U4829 (N_4829,N_4545,N_4536);
or U4830 (N_4830,N_4697,N_4530);
and U4831 (N_4831,N_4650,N_4582);
xnor U4832 (N_4832,N_4594,N_4602);
nand U4833 (N_4833,N_4635,N_4681);
and U4834 (N_4834,N_4716,N_4730);
and U4835 (N_4835,N_4526,N_4722);
and U4836 (N_4836,N_4631,N_4726);
or U4837 (N_4837,N_4679,N_4553);
xor U4838 (N_4838,N_4599,N_4559);
nor U4839 (N_4839,N_4715,N_4664);
and U4840 (N_4840,N_4606,N_4604);
nand U4841 (N_4841,N_4537,N_4737);
nor U4842 (N_4842,N_4551,N_4661);
and U4843 (N_4843,N_4615,N_4569);
nor U4844 (N_4844,N_4552,N_4609);
or U4845 (N_4845,N_4746,N_4580);
nor U4846 (N_4846,N_4709,N_4503);
and U4847 (N_4847,N_4748,N_4654);
and U4848 (N_4848,N_4519,N_4543);
and U4849 (N_4849,N_4742,N_4572);
nor U4850 (N_4850,N_4696,N_4627);
nand U4851 (N_4851,N_4717,N_4689);
nand U4852 (N_4852,N_4568,N_4706);
or U4853 (N_4853,N_4723,N_4633);
or U4854 (N_4854,N_4699,N_4541);
nor U4855 (N_4855,N_4663,N_4626);
or U4856 (N_4856,N_4628,N_4581);
nand U4857 (N_4857,N_4693,N_4573);
and U4858 (N_4858,N_4659,N_4644);
or U4859 (N_4859,N_4624,N_4729);
or U4860 (N_4860,N_4556,N_4587);
and U4861 (N_4861,N_4641,N_4642);
nor U4862 (N_4862,N_4684,N_4714);
nand U4863 (N_4863,N_4630,N_4666);
or U4864 (N_4864,N_4640,N_4600);
nand U4865 (N_4865,N_4739,N_4520);
nand U4866 (N_4866,N_4507,N_4517);
nand U4867 (N_4867,N_4505,N_4727);
or U4868 (N_4868,N_4548,N_4649);
nor U4869 (N_4869,N_4667,N_4578);
and U4870 (N_4870,N_4685,N_4561);
or U4871 (N_4871,N_4672,N_4557);
and U4872 (N_4872,N_4588,N_4612);
nor U4873 (N_4873,N_4732,N_4637);
nor U4874 (N_4874,N_4614,N_4593);
or U4875 (N_4875,N_4715,N_4735);
nand U4876 (N_4876,N_4664,N_4551);
or U4877 (N_4877,N_4664,N_4602);
nand U4878 (N_4878,N_4506,N_4503);
and U4879 (N_4879,N_4668,N_4714);
nand U4880 (N_4880,N_4519,N_4579);
xor U4881 (N_4881,N_4630,N_4662);
nor U4882 (N_4882,N_4507,N_4738);
nor U4883 (N_4883,N_4642,N_4513);
nor U4884 (N_4884,N_4616,N_4531);
or U4885 (N_4885,N_4579,N_4689);
nor U4886 (N_4886,N_4616,N_4686);
nand U4887 (N_4887,N_4686,N_4673);
nand U4888 (N_4888,N_4665,N_4538);
nand U4889 (N_4889,N_4565,N_4686);
and U4890 (N_4890,N_4701,N_4524);
nand U4891 (N_4891,N_4725,N_4612);
or U4892 (N_4892,N_4654,N_4644);
and U4893 (N_4893,N_4574,N_4649);
and U4894 (N_4894,N_4668,N_4653);
and U4895 (N_4895,N_4710,N_4589);
or U4896 (N_4896,N_4555,N_4708);
and U4897 (N_4897,N_4738,N_4510);
nand U4898 (N_4898,N_4711,N_4680);
and U4899 (N_4899,N_4714,N_4509);
nor U4900 (N_4900,N_4726,N_4724);
nor U4901 (N_4901,N_4719,N_4662);
and U4902 (N_4902,N_4728,N_4515);
and U4903 (N_4903,N_4617,N_4520);
nor U4904 (N_4904,N_4653,N_4695);
and U4905 (N_4905,N_4732,N_4606);
nand U4906 (N_4906,N_4556,N_4710);
nand U4907 (N_4907,N_4736,N_4554);
nand U4908 (N_4908,N_4743,N_4690);
or U4909 (N_4909,N_4724,N_4645);
nor U4910 (N_4910,N_4692,N_4658);
and U4911 (N_4911,N_4745,N_4525);
and U4912 (N_4912,N_4627,N_4660);
and U4913 (N_4913,N_4714,N_4533);
and U4914 (N_4914,N_4687,N_4707);
or U4915 (N_4915,N_4734,N_4619);
or U4916 (N_4916,N_4549,N_4576);
or U4917 (N_4917,N_4622,N_4540);
and U4918 (N_4918,N_4582,N_4675);
or U4919 (N_4919,N_4538,N_4723);
or U4920 (N_4920,N_4664,N_4734);
or U4921 (N_4921,N_4691,N_4505);
or U4922 (N_4922,N_4569,N_4563);
nor U4923 (N_4923,N_4714,N_4516);
and U4924 (N_4924,N_4696,N_4599);
nand U4925 (N_4925,N_4501,N_4500);
nor U4926 (N_4926,N_4743,N_4641);
and U4927 (N_4927,N_4695,N_4698);
or U4928 (N_4928,N_4525,N_4705);
nand U4929 (N_4929,N_4596,N_4627);
and U4930 (N_4930,N_4639,N_4600);
or U4931 (N_4931,N_4579,N_4725);
nor U4932 (N_4932,N_4705,N_4628);
nor U4933 (N_4933,N_4602,N_4587);
nor U4934 (N_4934,N_4504,N_4638);
or U4935 (N_4935,N_4612,N_4690);
or U4936 (N_4936,N_4509,N_4624);
and U4937 (N_4937,N_4555,N_4618);
or U4938 (N_4938,N_4691,N_4528);
and U4939 (N_4939,N_4615,N_4697);
and U4940 (N_4940,N_4590,N_4656);
or U4941 (N_4941,N_4530,N_4648);
or U4942 (N_4942,N_4571,N_4565);
or U4943 (N_4943,N_4514,N_4561);
and U4944 (N_4944,N_4504,N_4532);
and U4945 (N_4945,N_4592,N_4618);
nor U4946 (N_4946,N_4645,N_4684);
nor U4947 (N_4947,N_4563,N_4501);
and U4948 (N_4948,N_4511,N_4662);
and U4949 (N_4949,N_4562,N_4639);
nand U4950 (N_4950,N_4604,N_4585);
nand U4951 (N_4951,N_4747,N_4703);
or U4952 (N_4952,N_4649,N_4640);
and U4953 (N_4953,N_4564,N_4605);
or U4954 (N_4954,N_4645,N_4727);
or U4955 (N_4955,N_4716,N_4529);
nand U4956 (N_4956,N_4612,N_4746);
and U4957 (N_4957,N_4720,N_4574);
nor U4958 (N_4958,N_4605,N_4681);
nor U4959 (N_4959,N_4701,N_4573);
or U4960 (N_4960,N_4611,N_4672);
and U4961 (N_4961,N_4600,N_4721);
nor U4962 (N_4962,N_4541,N_4617);
nand U4963 (N_4963,N_4591,N_4567);
nor U4964 (N_4964,N_4642,N_4530);
or U4965 (N_4965,N_4553,N_4521);
nand U4966 (N_4966,N_4638,N_4521);
nand U4967 (N_4967,N_4633,N_4721);
nor U4968 (N_4968,N_4723,N_4582);
or U4969 (N_4969,N_4522,N_4741);
nand U4970 (N_4970,N_4740,N_4664);
or U4971 (N_4971,N_4744,N_4709);
nand U4972 (N_4972,N_4742,N_4532);
nor U4973 (N_4973,N_4731,N_4504);
or U4974 (N_4974,N_4631,N_4604);
nor U4975 (N_4975,N_4660,N_4735);
and U4976 (N_4976,N_4646,N_4667);
and U4977 (N_4977,N_4503,N_4542);
nand U4978 (N_4978,N_4698,N_4630);
and U4979 (N_4979,N_4526,N_4694);
and U4980 (N_4980,N_4650,N_4501);
nand U4981 (N_4981,N_4719,N_4710);
nor U4982 (N_4982,N_4658,N_4694);
xnor U4983 (N_4983,N_4722,N_4647);
xnor U4984 (N_4984,N_4718,N_4699);
or U4985 (N_4985,N_4564,N_4747);
and U4986 (N_4986,N_4668,N_4605);
xnor U4987 (N_4987,N_4724,N_4520);
nand U4988 (N_4988,N_4509,N_4586);
xnor U4989 (N_4989,N_4603,N_4723);
or U4990 (N_4990,N_4747,N_4522);
or U4991 (N_4991,N_4625,N_4658);
and U4992 (N_4992,N_4527,N_4607);
or U4993 (N_4993,N_4614,N_4676);
and U4994 (N_4994,N_4665,N_4666);
or U4995 (N_4995,N_4663,N_4566);
and U4996 (N_4996,N_4502,N_4569);
nor U4997 (N_4997,N_4628,N_4515);
nand U4998 (N_4998,N_4644,N_4619);
nand U4999 (N_4999,N_4656,N_4748);
or U5000 (N_5000,N_4766,N_4953);
and U5001 (N_5001,N_4773,N_4963);
nand U5002 (N_5002,N_4911,N_4800);
and U5003 (N_5003,N_4883,N_4961);
or U5004 (N_5004,N_4970,N_4787);
or U5005 (N_5005,N_4808,N_4954);
nor U5006 (N_5006,N_4930,N_4843);
or U5007 (N_5007,N_4905,N_4979);
nor U5008 (N_5008,N_4775,N_4925);
nor U5009 (N_5009,N_4794,N_4856);
nor U5010 (N_5010,N_4875,N_4886);
and U5011 (N_5011,N_4922,N_4982);
nor U5012 (N_5012,N_4806,N_4943);
and U5013 (N_5013,N_4802,N_4910);
nor U5014 (N_5014,N_4816,N_4926);
nor U5015 (N_5015,N_4940,N_4769);
and U5016 (N_5016,N_4859,N_4965);
or U5017 (N_5017,N_4903,N_4960);
or U5018 (N_5018,N_4871,N_4818);
nor U5019 (N_5019,N_4945,N_4861);
nand U5020 (N_5020,N_4869,N_4784);
or U5021 (N_5021,N_4948,N_4919);
nand U5022 (N_5022,N_4901,N_4882);
and U5023 (N_5023,N_4830,N_4900);
nand U5024 (N_5024,N_4754,N_4924);
nand U5025 (N_5025,N_4967,N_4796);
or U5026 (N_5026,N_4938,N_4975);
or U5027 (N_5027,N_4892,N_4837);
nor U5028 (N_5028,N_4986,N_4931);
nor U5029 (N_5029,N_4854,N_4973);
nor U5030 (N_5030,N_4848,N_4791);
nor U5031 (N_5031,N_4913,N_4809);
nor U5032 (N_5032,N_4998,N_4864);
nand U5033 (N_5033,N_4904,N_4958);
and U5034 (N_5034,N_4857,N_4815);
and U5035 (N_5035,N_4813,N_4946);
nand U5036 (N_5036,N_4881,N_4836);
nor U5037 (N_5037,N_4990,N_4797);
nor U5038 (N_5038,N_4758,N_4751);
and U5039 (N_5039,N_4974,N_4752);
and U5040 (N_5040,N_4980,N_4778);
nor U5041 (N_5041,N_4834,N_4753);
and U5042 (N_5042,N_4803,N_4937);
nand U5043 (N_5043,N_4914,N_4842);
nand U5044 (N_5044,N_4876,N_4829);
and U5045 (N_5045,N_4865,N_4933);
nand U5046 (N_5046,N_4821,N_4838);
or U5047 (N_5047,N_4855,N_4862);
and U5048 (N_5048,N_4971,N_4899);
and U5049 (N_5049,N_4868,N_4777);
and U5050 (N_5050,N_4764,N_4920);
nand U5051 (N_5051,N_4983,N_4955);
nand U5052 (N_5052,N_4906,N_4957);
nand U5053 (N_5053,N_4844,N_4894);
or U5054 (N_5054,N_4944,N_4879);
and U5055 (N_5055,N_4941,N_4968);
nand U5056 (N_5056,N_4959,N_4759);
nand U5057 (N_5057,N_4755,N_4782);
nand U5058 (N_5058,N_4962,N_4846);
nand U5059 (N_5059,N_4994,N_4776);
nand U5060 (N_5060,N_4780,N_4811);
nand U5061 (N_5061,N_4935,N_4912);
nor U5062 (N_5062,N_4889,N_4793);
nand U5063 (N_5063,N_4972,N_4887);
nor U5064 (N_5064,N_4828,N_4898);
and U5065 (N_5065,N_4795,N_4885);
nand U5066 (N_5066,N_4772,N_4849);
and U5067 (N_5067,N_4798,N_4841);
nor U5068 (N_5068,N_4950,N_4774);
nor U5069 (N_5069,N_4907,N_4872);
nor U5070 (N_5070,N_4999,N_4890);
nor U5071 (N_5071,N_4987,N_4978);
and U5072 (N_5072,N_4845,N_4863);
or U5073 (N_5073,N_4750,N_4989);
and U5074 (N_5074,N_4847,N_4824);
or U5075 (N_5075,N_4783,N_4820);
nor U5076 (N_5076,N_4947,N_4895);
nor U5077 (N_5077,N_4840,N_4921);
and U5078 (N_5078,N_4915,N_4814);
nand U5079 (N_5079,N_4851,N_4992);
and U5080 (N_5080,N_4917,N_4833);
or U5081 (N_5081,N_4767,N_4810);
or U5082 (N_5082,N_4760,N_4853);
nor U5083 (N_5083,N_4936,N_4880);
and U5084 (N_5084,N_4969,N_4805);
or U5085 (N_5085,N_4785,N_4991);
and U5086 (N_5086,N_4981,N_4779);
and U5087 (N_5087,N_4888,N_4762);
nand U5088 (N_5088,N_4790,N_4984);
or U5089 (N_5089,N_4812,N_4819);
nand U5090 (N_5090,N_4822,N_4909);
or U5091 (N_5091,N_4770,N_4934);
xnor U5092 (N_5092,N_4939,N_4825);
and U5093 (N_5093,N_4878,N_4817);
nand U5094 (N_5094,N_4757,N_4789);
nor U5095 (N_5095,N_4923,N_4952);
or U5096 (N_5096,N_4964,N_4997);
nor U5097 (N_5097,N_4756,N_4977);
or U5098 (N_5098,N_4891,N_4765);
and U5099 (N_5099,N_4799,N_4877);
and U5100 (N_5100,N_4839,N_4942);
nor U5101 (N_5101,N_4761,N_4993);
nand U5102 (N_5102,N_4771,N_4932);
nor U5103 (N_5103,N_4976,N_4788);
nor U5104 (N_5104,N_4781,N_4902);
nor U5105 (N_5105,N_4832,N_4858);
or U5106 (N_5106,N_4928,N_4786);
or U5107 (N_5107,N_4823,N_4867);
and U5108 (N_5108,N_4792,N_4897);
and U5109 (N_5109,N_4927,N_4966);
or U5110 (N_5110,N_4804,N_4831);
or U5111 (N_5111,N_4852,N_4860);
nand U5112 (N_5112,N_4866,N_4929);
and U5113 (N_5113,N_4996,N_4995);
nor U5114 (N_5114,N_4850,N_4988);
nand U5115 (N_5115,N_4951,N_4949);
or U5116 (N_5116,N_4916,N_4893);
and U5117 (N_5117,N_4956,N_4827);
or U5118 (N_5118,N_4835,N_4896);
or U5119 (N_5119,N_4870,N_4908);
and U5120 (N_5120,N_4918,N_4807);
or U5121 (N_5121,N_4801,N_4884);
and U5122 (N_5122,N_4874,N_4763);
nor U5123 (N_5123,N_4768,N_4985);
or U5124 (N_5124,N_4873,N_4826);
and U5125 (N_5125,N_4825,N_4769);
or U5126 (N_5126,N_4841,N_4971);
nor U5127 (N_5127,N_4781,N_4770);
nor U5128 (N_5128,N_4833,N_4924);
nor U5129 (N_5129,N_4864,N_4759);
xnor U5130 (N_5130,N_4880,N_4860);
and U5131 (N_5131,N_4805,N_4981);
nand U5132 (N_5132,N_4863,N_4894);
nand U5133 (N_5133,N_4765,N_4903);
nand U5134 (N_5134,N_4774,N_4996);
nand U5135 (N_5135,N_4990,N_4759);
or U5136 (N_5136,N_4977,N_4929);
nand U5137 (N_5137,N_4977,N_4782);
nand U5138 (N_5138,N_4888,N_4991);
or U5139 (N_5139,N_4915,N_4772);
nor U5140 (N_5140,N_4820,N_4789);
and U5141 (N_5141,N_4767,N_4871);
nor U5142 (N_5142,N_4884,N_4984);
nor U5143 (N_5143,N_4943,N_4989);
or U5144 (N_5144,N_4871,N_4814);
or U5145 (N_5145,N_4818,N_4896);
nand U5146 (N_5146,N_4907,N_4848);
and U5147 (N_5147,N_4871,N_4884);
or U5148 (N_5148,N_4973,N_4796);
or U5149 (N_5149,N_4858,N_4947);
and U5150 (N_5150,N_4817,N_4797);
nand U5151 (N_5151,N_4897,N_4912);
or U5152 (N_5152,N_4835,N_4901);
or U5153 (N_5153,N_4751,N_4845);
nor U5154 (N_5154,N_4947,N_4859);
or U5155 (N_5155,N_4927,N_4839);
nor U5156 (N_5156,N_4836,N_4813);
or U5157 (N_5157,N_4805,N_4874);
nand U5158 (N_5158,N_4976,N_4996);
nand U5159 (N_5159,N_4910,N_4751);
and U5160 (N_5160,N_4965,N_4768);
nand U5161 (N_5161,N_4767,N_4885);
or U5162 (N_5162,N_4930,N_4968);
nor U5163 (N_5163,N_4846,N_4986);
nor U5164 (N_5164,N_4984,N_4802);
nor U5165 (N_5165,N_4909,N_4939);
nand U5166 (N_5166,N_4927,N_4945);
and U5167 (N_5167,N_4836,N_4915);
and U5168 (N_5168,N_4993,N_4904);
nor U5169 (N_5169,N_4881,N_4834);
or U5170 (N_5170,N_4825,N_4927);
nor U5171 (N_5171,N_4773,N_4900);
nor U5172 (N_5172,N_4839,N_4786);
and U5173 (N_5173,N_4987,N_4762);
nand U5174 (N_5174,N_4888,N_4957);
or U5175 (N_5175,N_4781,N_4766);
or U5176 (N_5176,N_4828,N_4840);
nand U5177 (N_5177,N_4847,N_4777);
or U5178 (N_5178,N_4766,N_4938);
or U5179 (N_5179,N_4870,N_4768);
or U5180 (N_5180,N_4761,N_4937);
nor U5181 (N_5181,N_4861,N_4930);
or U5182 (N_5182,N_4939,N_4873);
or U5183 (N_5183,N_4876,N_4755);
and U5184 (N_5184,N_4836,N_4848);
or U5185 (N_5185,N_4972,N_4982);
nor U5186 (N_5186,N_4907,N_4974);
nand U5187 (N_5187,N_4855,N_4879);
nor U5188 (N_5188,N_4945,N_4942);
and U5189 (N_5189,N_4782,N_4919);
nor U5190 (N_5190,N_4922,N_4800);
and U5191 (N_5191,N_4772,N_4833);
or U5192 (N_5192,N_4971,N_4755);
nor U5193 (N_5193,N_4992,N_4906);
or U5194 (N_5194,N_4900,N_4755);
nand U5195 (N_5195,N_4834,N_4814);
and U5196 (N_5196,N_4791,N_4846);
or U5197 (N_5197,N_4947,N_4844);
nor U5198 (N_5198,N_4944,N_4821);
nor U5199 (N_5199,N_4848,N_4853);
nor U5200 (N_5200,N_4913,N_4879);
and U5201 (N_5201,N_4973,N_4892);
nor U5202 (N_5202,N_4898,N_4761);
and U5203 (N_5203,N_4988,N_4986);
and U5204 (N_5204,N_4986,N_4767);
nand U5205 (N_5205,N_4907,N_4903);
nand U5206 (N_5206,N_4859,N_4930);
nand U5207 (N_5207,N_4814,N_4974);
or U5208 (N_5208,N_4895,N_4788);
nand U5209 (N_5209,N_4862,N_4772);
or U5210 (N_5210,N_4986,N_4800);
nor U5211 (N_5211,N_4905,N_4871);
xnor U5212 (N_5212,N_4981,N_4892);
nor U5213 (N_5213,N_4977,N_4792);
or U5214 (N_5214,N_4823,N_4873);
and U5215 (N_5215,N_4802,N_4800);
nand U5216 (N_5216,N_4946,N_4861);
nand U5217 (N_5217,N_4971,N_4973);
and U5218 (N_5218,N_4949,N_4878);
nor U5219 (N_5219,N_4805,N_4768);
and U5220 (N_5220,N_4905,N_4858);
or U5221 (N_5221,N_4997,N_4824);
nand U5222 (N_5222,N_4809,N_4905);
nor U5223 (N_5223,N_4950,N_4870);
or U5224 (N_5224,N_4777,N_4945);
nand U5225 (N_5225,N_4791,N_4875);
nor U5226 (N_5226,N_4761,N_4769);
nor U5227 (N_5227,N_4891,N_4780);
or U5228 (N_5228,N_4910,N_4927);
nand U5229 (N_5229,N_4904,N_4994);
nor U5230 (N_5230,N_4922,N_4763);
nor U5231 (N_5231,N_4782,N_4891);
nand U5232 (N_5232,N_4967,N_4775);
and U5233 (N_5233,N_4768,N_4964);
or U5234 (N_5234,N_4918,N_4869);
or U5235 (N_5235,N_4839,N_4986);
nor U5236 (N_5236,N_4899,N_4786);
nand U5237 (N_5237,N_4823,N_4875);
or U5238 (N_5238,N_4981,N_4975);
or U5239 (N_5239,N_4792,N_4906);
nand U5240 (N_5240,N_4804,N_4895);
or U5241 (N_5241,N_4928,N_4886);
or U5242 (N_5242,N_4975,N_4919);
nor U5243 (N_5243,N_4986,N_4989);
or U5244 (N_5244,N_4750,N_4758);
nand U5245 (N_5245,N_4882,N_4764);
nand U5246 (N_5246,N_4762,N_4944);
and U5247 (N_5247,N_4785,N_4919);
nor U5248 (N_5248,N_4776,N_4901);
nor U5249 (N_5249,N_4992,N_4804);
nand U5250 (N_5250,N_5164,N_5202);
or U5251 (N_5251,N_5126,N_5035);
or U5252 (N_5252,N_5226,N_5163);
nor U5253 (N_5253,N_5076,N_5200);
or U5254 (N_5254,N_5101,N_5123);
nor U5255 (N_5255,N_5143,N_5033);
or U5256 (N_5256,N_5026,N_5037);
or U5257 (N_5257,N_5241,N_5045);
and U5258 (N_5258,N_5144,N_5220);
and U5259 (N_5259,N_5223,N_5088);
nor U5260 (N_5260,N_5134,N_5083);
and U5261 (N_5261,N_5050,N_5116);
and U5262 (N_5262,N_5136,N_5153);
nor U5263 (N_5263,N_5063,N_5169);
nor U5264 (N_5264,N_5181,N_5117);
nor U5265 (N_5265,N_5173,N_5093);
nor U5266 (N_5266,N_5216,N_5174);
nand U5267 (N_5267,N_5219,N_5238);
or U5268 (N_5268,N_5006,N_5046);
xnor U5269 (N_5269,N_5055,N_5078);
nor U5270 (N_5270,N_5179,N_5073);
nor U5271 (N_5271,N_5043,N_5038);
nand U5272 (N_5272,N_5162,N_5007);
or U5273 (N_5273,N_5131,N_5068);
nand U5274 (N_5274,N_5044,N_5086);
and U5275 (N_5275,N_5079,N_5108);
nor U5276 (N_5276,N_5067,N_5036);
nor U5277 (N_5277,N_5170,N_5167);
or U5278 (N_5278,N_5203,N_5205);
xnor U5279 (N_5279,N_5127,N_5064);
nand U5280 (N_5280,N_5227,N_5014);
nand U5281 (N_5281,N_5018,N_5056);
and U5282 (N_5282,N_5146,N_5081);
nor U5283 (N_5283,N_5189,N_5102);
nand U5284 (N_5284,N_5210,N_5247);
or U5285 (N_5285,N_5011,N_5152);
and U5286 (N_5286,N_5154,N_5161);
nor U5287 (N_5287,N_5147,N_5091);
or U5288 (N_5288,N_5071,N_5157);
nand U5289 (N_5289,N_5158,N_5021);
nand U5290 (N_5290,N_5048,N_5185);
or U5291 (N_5291,N_5066,N_5115);
or U5292 (N_5292,N_5195,N_5032);
nor U5293 (N_5293,N_5053,N_5072);
or U5294 (N_5294,N_5142,N_5025);
nand U5295 (N_5295,N_5125,N_5233);
and U5296 (N_5296,N_5121,N_5224);
and U5297 (N_5297,N_5246,N_5201);
and U5298 (N_5298,N_5130,N_5028);
and U5299 (N_5299,N_5057,N_5094);
or U5300 (N_5300,N_5090,N_5074);
nor U5301 (N_5301,N_5128,N_5236);
nand U5302 (N_5302,N_5141,N_5119);
nor U5303 (N_5303,N_5022,N_5168);
and U5304 (N_5304,N_5193,N_5133);
or U5305 (N_5305,N_5058,N_5020);
and U5306 (N_5306,N_5062,N_5124);
xnor U5307 (N_5307,N_5249,N_5225);
nor U5308 (N_5308,N_5148,N_5176);
nor U5309 (N_5309,N_5013,N_5184);
or U5310 (N_5310,N_5190,N_5001);
or U5311 (N_5311,N_5120,N_5217);
and U5312 (N_5312,N_5109,N_5030);
or U5313 (N_5313,N_5106,N_5103);
or U5314 (N_5314,N_5230,N_5017);
nor U5315 (N_5315,N_5237,N_5034);
nand U5316 (N_5316,N_5098,N_5151);
nor U5317 (N_5317,N_5159,N_5183);
or U5318 (N_5318,N_5019,N_5080);
and U5319 (N_5319,N_5150,N_5077);
nand U5320 (N_5320,N_5009,N_5160);
nor U5321 (N_5321,N_5140,N_5051);
and U5322 (N_5322,N_5244,N_5047);
and U5323 (N_5323,N_5214,N_5084);
or U5324 (N_5324,N_5138,N_5222);
nor U5325 (N_5325,N_5110,N_5052);
nor U5326 (N_5326,N_5192,N_5187);
nor U5327 (N_5327,N_5008,N_5012);
and U5328 (N_5328,N_5029,N_5059);
or U5329 (N_5329,N_5186,N_5003);
or U5330 (N_5330,N_5129,N_5027);
and U5331 (N_5331,N_5218,N_5239);
and U5332 (N_5332,N_5092,N_5191);
nor U5333 (N_5333,N_5112,N_5175);
nand U5334 (N_5334,N_5070,N_5165);
or U5335 (N_5335,N_5105,N_5228);
nand U5336 (N_5336,N_5206,N_5075);
and U5337 (N_5337,N_5211,N_5061);
nor U5338 (N_5338,N_5135,N_5213);
or U5339 (N_5339,N_5229,N_5005);
nor U5340 (N_5340,N_5010,N_5221);
nand U5341 (N_5341,N_5235,N_5095);
xor U5342 (N_5342,N_5232,N_5039);
nand U5343 (N_5343,N_5215,N_5082);
nor U5344 (N_5344,N_5099,N_5182);
or U5345 (N_5345,N_5245,N_5100);
and U5346 (N_5346,N_5031,N_5197);
nand U5347 (N_5347,N_5137,N_5002);
nand U5348 (N_5348,N_5234,N_5188);
and U5349 (N_5349,N_5016,N_5097);
or U5350 (N_5350,N_5114,N_5107);
nor U5351 (N_5351,N_5004,N_5089);
and U5352 (N_5352,N_5209,N_5023);
and U5353 (N_5353,N_5207,N_5196);
or U5354 (N_5354,N_5118,N_5122);
or U5355 (N_5355,N_5149,N_5243);
nand U5356 (N_5356,N_5171,N_5156);
nand U5357 (N_5357,N_5240,N_5015);
or U5358 (N_5358,N_5212,N_5178);
or U5359 (N_5359,N_5177,N_5069);
and U5360 (N_5360,N_5054,N_5111);
or U5361 (N_5361,N_5049,N_5198);
and U5362 (N_5362,N_5113,N_5248);
or U5363 (N_5363,N_5208,N_5132);
and U5364 (N_5364,N_5060,N_5041);
and U5365 (N_5365,N_5096,N_5231);
nor U5366 (N_5366,N_5204,N_5085);
nor U5367 (N_5367,N_5194,N_5042);
nand U5368 (N_5368,N_5242,N_5145);
and U5369 (N_5369,N_5087,N_5139);
and U5370 (N_5370,N_5000,N_5180);
nor U5371 (N_5371,N_5024,N_5040);
nand U5372 (N_5372,N_5155,N_5104);
nand U5373 (N_5373,N_5199,N_5166);
or U5374 (N_5374,N_5172,N_5065);
nor U5375 (N_5375,N_5163,N_5188);
or U5376 (N_5376,N_5119,N_5062);
nor U5377 (N_5377,N_5017,N_5220);
nand U5378 (N_5378,N_5192,N_5199);
nor U5379 (N_5379,N_5094,N_5093);
nand U5380 (N_5380,N_5188,N_5105);
and U5381 (N_5381,N_5121,N_5041);
nor U5382 (N_5382,N_5222,N_5086);
or U5383 (N_5383,N_5194,N_5186);
and U5384 (N_5384,N_5068,N_5034);
and U5385 (N_5385,N_5025,N_5186);
nor U5386 (N_5386,N_5093,N_5210);
and U5387 (N_5387,N_5016,N_5163);
or U5388 (N_5388,N_5057,N_5208);
nor U5389 (N_5389,N_5238,N_5161);
xnor U5390 (N_5390,N_5081,N_5065);
or U5391 (N_5391,N_5063,N_5012);
nand U5392 (N_5392,N_5055,N_5026);
nor U5393 (N_5393,N_5081,N_5230);
or U5394 (N_5394,N_5137,N_5064);
and U5395 (N_5395,N_5036,N_5224);
or U5396 (N_5396,N_5023,N_5200);
and U5397 (N_5397,N_5005,N_5038);
and U5398 (N_5398,N_5041,N_5013);
nor U5399 (N_5399,N_5222,N_5103);
nand U5400 (N_5400,N_5066,N_5127);
and U5401 (N_5401,N_5227,N_5151);
nand U5402 (N_5402,N_5066,N_5197);
nor U5403 (N_5403,N_5189,N_5156);
nand U5404 (N_5404,N_5119,N_5035);
and U5405 (N_5405,N_5188,N_5025);
nor U5406 (N_5406,N_5142,N_5108);
or U5407 (N_5407,N_5032,N_5125);
nand U5408 (N_5408,N_5104,N_5182);
nor U5409 (N_5409,N_5040,N_5168);
and U5410 (N_5410,N_5143,N_5160);
nand U5411 (N_5411,N_5121,N_5099);
or U5412 (N_5412,N_5223,N_5181);
or U5413 (N_5413,N_5004,N_5024);
or U5414 (N_5414,N_5239,N_5067);
or U5415 (N_5415,N_5219,N_5173);
and U5416 (N_5416,N_5234,N_5016);
and U5417 (N_5417,N_5197,N_5006);
nor U5418 (N_5418,N_5100,N_5029);
nand U5419 (N_5419,N_5065,N_5210);
or U5420 (N_5420,N_5248,N_5030);
and U5421 (N_5421,N_5166,N_5101);
or U5422 (N_5422,N_5113,N_5164);
nand U5423 (N_5423,N_5199,N_5049);
nor U5424 (N_5424,N_5199,N_5185);
nor U5425 (N_5425,N_5200,N_5133);
or U5426 (N_5426,N_5239,N_5157);
nor U5427 (N_5427,N_5155,N_5024);
and U5428 (N_5428,N_5160,N_5208);
and U5429 (N_5429,N_5188,N_5231);
and U5430 (N_5430,N_5231,N_5243);
nor U5431 (N_5431,N_5167,N_5175);
nor U5432 (N_5432,N_5032,N_5176);
nor U5433 (N_5433,N_5160,N_5153);
nor U5434 (N_5434,N_5048,N_5145);
nand U5435 (N_5435,N_5069,N_5016);
nor U5436 (N_5436,N_5117,N_5030);
and U5437 (N_5437,N_5113,N_5173);
and U5438 (N_5438,N_5210,N_5226);
or U5439 (N_5439,N_5130,N_5240);
or U5440 (N_5440,N_5193,N_5205);
nand U5441 (N_5441,N_5171,N_5064);
nand U5442 (N_5442,N_5004,N_5099);
nor U5443 (N_5443,N_5162,N_5126);
nor U5444 (N_5444,N_5045,N_5046);
or U5445 (N_5445,N_5157,N_5191);
and U5446 (N_5446,N_5115,N_5203);
and U5447 (N_5447,N_5109,N_5071);
or U5448 (N_5448,N_5181,N_5086);
nor U5449 (N_5449,N_5026,N_5219);
nor U5450 (N_5450,N_5071,N_5014);
and U5451 (N_5451,N_5110,N_5103);
or U5452 (N_5452,N_5003,N_5045);
or U5453 (N_5453,N_5236,N_5057);
nor U5454 (N_5454,N_5114,N_5090);
nor U5455 (N_5455,N_5080,N_5168);
and U5456 (N_5456,N_5136,N_5174);
nand U5457 (N_5457,N_5019,N_5125);
or U5458 (N_5458,N_5172,N_5149);
nand U5459 (N_5459,N_5223,N_5025);
or U5460 (N_5460,N_5137,N_5009);
nand U5461 (N_5461,N_5196,N_5181);
nor U5462 (N_5462,N_5223,N_5006);
nor U5463 (N_5463,N_5077,N_5162);
nand U5464 (N_5464,N_5110,N_5011);
xor U5465 (N_5465,N_5079,N_5202);
or U5466 (N_5466,N_5063,N_5133);
and U5467 (N_5467,N_5184,N_5131);
nor U5468 (N_5468,N_5029,N_5114);
and U5469 (N_5469,N_5126,N_5086);
or U5470 (N_5470,N_5055,N_5228);
xor U5471 (N_5471,N_5240,N_5083);
nor U5472 (N_5472,N_5207,N_5137);
or U5473 (N_5473,N_5221,N_5050);
and U5474 (N_5474,N_5101,N_5238);
and U5475 (N_5475,N_5009,N_5034);
and U5476 (N_5476,N_5161,N_5019);
or U5477 (N_5477,N_5124,N_5086);
nand U5478 (N_5478,N_5039,N_5220);
nand U5479 (N_5479,N_5147,N_5099);
or U5480 (N_5480,N_5096,N_5016);
or U5481 (N_5481,N_5082,N_5005);
and U5482 (N_5482,N_5013,N_5093);
nand U5483 (N_5483,N_5032,N_5158);
or U5484 (N_5484,N_5192,N_5201);
nand U5485 (N_5485,N_5035,N_5175);
or U5486 (N_5486,N_5101,N_5041);
nor U5487 (N_5487,N_5048,N_5148);
or U5488 (N_5488,N_5061,N_5205);
and U5489 (N_5489,N_5153,N_5132);
or U5490 (N_5490,N_5067,N_5225);
or U5491 (N_5491,N_5011,N_5112);
nand U5492 (N_5492,N_5001,N_5053);
nor U5493 (N_5493,N_5215,N_5153);
or U5494 (N_5494,N_5197,N_5232);
nor U5495 (N_5495,N_5098,N_5161);
nand U5496 (N_5496,N_5229,N_5057);
or U5497 (N_5497,N_5069,N_5075);
nand U5498 (N_5498,N_5232,N_5087);
nand U5499 (N_5499,N_5140,N_5055);
xor U5500 (N_5500,N_5384,N_5393);
or U5501 (N_5501,N_5389,N_5490);
and U5502 (N_5502,N_5317,N_5252);
nor U5503 (N_5503,N_5479,N_5411);
nor U5504 (N_5504,N_5325,N_5355);
nor U5505 (N_5505,N_5354,N_5254);
nand U5506 (N_5506,N_5425,N_5265);
and U5507 (N_5507,N_5263,N_5272);
nand U5508 (N_5508,N_5438,N_5312);
nor U5509 (N_5509,N_5324,N_5498);
nand U5510 (N_5510,N_5337,N_5465);
and U5511 (N_5511,N_5435,N_5437);
nor U5512 (N_5512,N_5305,N_5304);
nand U5513 (N_5513,N_5471,N_5373);
nand U5514 (N_5514,N_5356,N_5366);
or U5515 (N_5515,N_5341,N_5378);
and U5516 (N_5516,N_5381,N_5274);
nor U5517 (N_5517,N_5408,N_5387);
nand U5518 (N_5518,N_5333,N_5376);
and U5519 (N_5519,N_5262,N_5415);
and U5520 (N_5520,N_5307,N_5273);
nor U5521 (N_5521,N_5461,N_5445);
nor U5522 (N_5522,N_5342,N_5475);
or U5523 (N_5523,N_5266,N_5357);
nand U5524 (N_5524,N_5386,N_5298);
nand U5525 (N_5525,N_5303,N_5410);
nand U5526 (N_5526,N_5493,N_5279);
and U5527 (N_5527,N_5494,N_5350);
or U5528 (N_5528,N_5396,N_5450);
nor U5529 (N_5529,N_5278,N_5383);
nor U5530 (N_5530,N_5469,N_5316);
or U5531 (N_5531,N_5453,N_5267);
or U5532 (N_5532,N_5491,N_5323);
nand U5533 (N_5533,N_5463,N_5289);
xor U5534 (N_5534,N_5483,N_5372);
nand U5535 (N_5535,N_5467,N_5306);
nor U5536 (N_5536,N_5433,N_5331);
nor U5537 (N_5537,N_5375,N_5299);
nor U5538 (N_5538,N_5477,N_5426);
nand U5539 (N_5539,N_5363,N_5311);
or U5540 (N_5540,N_5476,N_5414);
or U5541 (N_5541,N_5346,N_5286);
or U5542 (N_5542,N_5351,N_5416);
and U5543 (N_5543,N_5462,N_5485);
nand U5544 (N_5544,N_5321,N_5487);
nand U5545 (N_5545,N_5427,N_5436);
or U5546 (N_5546,N_5472,N_5420);
nor U5547 (N_5547,N_5345,N_5295);
xnor U5548 (N_5548,N_5318,N_5454);
nand U5549 (N_5549,N_5404,N_5353);
or U5550 (N_5550,N_5447,N_5407);
nand U5551 (N_5551,N_5256,N_5470);
or U5552 (N_5552,N_5313,N_5259);
or U5553 (N_5553,N_5429,N_5369);
nand U5554 (N_5554,N_5365,N_5294);
or U5555 (N_5555,N_5388,N_5255);
nor U5556 (N_5556,N_5330,N_5495);
or U5557 (N_5557,N_5394,N_5322);
nand U5558 (N_5558,N_5257,N_5301);
and U5559 (N_5559,N_5293,N_5338);
or U5560 (N_5560,N_5360,N_5328);
or U5561 (N_5561,N_5385,N_5452);
and U5562 (N_5562,N_5348,N_5401);
nor U5563 (N_5563,N_5290,N_5443);
nor U5564 (N_5564,N_5280,N_5309);
or U5565 (N_5565,N_5496,N_5268);
nor U5566 (N_5566,N_5468,N_5347);
or U5567 (N_5567,N_5340,N_5497);
nor U5568 (N_5568,N_5292,N_5466);
nor U5569 (N_5569,N_5269,N_5264);
or U5570 (N_5570,N_5329,N_5302);
nor U5571 (N_5571,N_5260,N_5282);
and U5572 (N_5572,N_5283,N_5349);
nand U5573 (N_5573,N_5288,N_5406);
and U5574 (N_5574,N_5380,N_5364);
nand U5575 (N_5575,N_5412,N_5423);
nand U5576 (N_5576,N_5276,N_5326);
and U5577 (N_5577,N_5335,N_5275);
and U5578 (N_5578,N_5344,N_5456);
and U5579 (N_5579,N_5474,N_5339);
or U5580 (N_5580,N_5382,N_5367);
nand U5581 (N_5581,N_5368,N_5319);
nor U5582 (N_5582,N_5361,N_5358);
nor U5583 (N_5583,N_5400,N_5419);
nand U5584 (N_5584,N_5359,N_5297);
and U5585 (N_5585,N_5455,N_5459);
or U5586 (N_5586,N_5362,N_5424);
and U5587 (N_5587,N_5308,N_5473);
nand U5588 (N_5588,N_5489,N_5417);
nand U5589 (N_5589,N_5391,N_5440);
and U5590 (N_5590,N_5374,N_5277);
nor U5591 (N_5591,N_5480,N_5392);
and U5592 (N_5592,N_5499,N_5336);
nor U5593 (N_5593,N_5315,N_5270);
nor U5594 (N_5594,N_5399,N_5352);
and U5595 (N_5595,N_5430,N_5250);
nand U5596 (N_5596,N_5261,N_5284);
and U5597 (N_5597,N_5464,N_5441);
nor U5598 (N_5598,N_5451,N_5409);
or U5599 (N_5599,N_5334,N_5332);
and U5600 (N_5600,N_5478,N_5442);
and U5601 (N_5601,N_5413,N_5291);
nor U5602 (N_5602,N_5398,N_5320);
nor U5603 (N_5603,N_5481,N_5484);
nand U5604 (N_5604,N_5296,N_5314);
nand U5605 (N_5605,N_5327,N_5251);
nor U5606 (N_5606,N_5418,N_5300);
nor U5607 (N_5607,N_5448,N_5253);
nor U5608 (N_5608,N_5281,N_5449);
nor U5609 (N_5609,N_5444,N_5379);
or U5610 (N_5610,N_5371,N_5258);
nor U5611 (N_5611,N_5432,N_5343);
nand U5612 (N_5612,N_5457,N_5285);
or U5613 (N_5613,N_5421,N_5460);
nor U5614 (N_5614,N_5422,N_5482);
nand U5615 (N_5615,N_5488,N_5434);
xnor U5616 (N_5616,N_5397,N_5405);
or U5617 (N_5617,N_5439,N_5428);
and U5618 (N_5618,N_5486,N_5446);
and U5619 (N_5619,N_5458,N_5492);
and U5620 (N_5620,N_5403,N_5431);
nand U5621 (N_5621,N_5271,N_5390);
nor U5622 (N_5622,N_5310,N_5370);
nor U5623 (N_5623,N_5402,N_5287);
nor U5624 (N_5624,N_5395,N_5377);
nor U5625 (N_5625,N_5427,N_5435);
or U5626 (N_5626,N_5389,N_5452);
nand U5627 (N_5627,N_5400,N_5413);
or U5628 (N_5628,N_5387,N_5306);
nand U5629 (N_5629,N_5280,N_5481);
or U5630 (N_5630,N_5467,N_5486);
and U5631 (N_5631,N_5343,N_5439);
or U5632 (N_5632,N_5449,N_5492);
nor U5633 (N_5633,N_5316,N_5434);
or U5634 (N_5634,N_5398,N_5401);
nor U5635 (N_5635,N_5496,N_5284);
nand U5636 (N_5636,N_5263,N_5435);
or U5637 (N_5637,N_5407,N_5380);
nand U5638 (N_5638,N_5309,N_5458);
xor U5639 (N_5639,N_5388,N_5398);
nor U5640 (N_5640,N_5277,N_5347);
or U5641 (N_5641,N_5423,N_5254);
or U5642 (N_5642,N_5407,N_5486);
nor U5643 (N_5643,N_5411,N_5335);
and U5644 (N_5644,N_5430,N_5478);
and U5645 (N_5645,N_5392,N_5325);
nand U5646 (N_5646,N_5446,N_5414);
and U5647 (N_5647,N_5477,N_5344);
and U5648 (N_5648,N_5311,N_5359);
nand U5649 (N_5649,N_5409,N_5381);
nor U5650 (N_5650,N_5295,N_5422);
nand U5651 (N_5651,N_5368,N_5281);
and U5652 (N_5652,N_5276,N_5471);
nand U5653 (N_5653,N_5271,N_5262);
and U5654 (N_5654,N_5400,N_5388);
nor U5655 (N_5655,N_5319,N_5385);
nand U5656 (N_5656,N_5293,N_5464);
nand U5657 (N_5657,N_5286,N_5416);
and U5658 (N_5658,N_5264,N_5488);
and U5659 (N_5659,N_5468,N_5318);
and U5660 (N_5660,N_5403,N_5300);
or U5661 (N_5661,N_5492,N_5267);
or U5662 (N_5662,N_5481,N_5400);
xnor U5663 (N_5663,N_5400,N_5476);
nor U5664 (N_5664,N_5468,N_5432);
nand U5665 (N_5665,N_5434,N_5294);
or U5666 (N_5666,N_5462,N_5277);
nor U5667 (N_5667,N_5445,N_5252);
nor U5668 (N_5668,N_5318,N_5438);
and U5669 (N_5669,N_5383,N_5297);
and U5670 (N_5670,N_5260,N_5256);
or U5671 (N_5671,N_5442,N_5449);
nand U5672 (N_5672,N_5267,N_5259);
and U5673 (N_5673,N_5282,N_5465);
and U5674 (N_5674,N_5309,N_5421);
nand U5675 (N_5675,N_5287,N_5378);
and U5676 (N_5676,N_5486,N_5272);
nor U5677 (N_5677,N_5320,N_5311);
nor U5678 (N_5678,N_5478,N_5331);
nor U5679 (N_5679,N_5298,N_5292);
nor U5680 (N_5680,N_5364,N_5446);
nor U5681 (N_5681,N_5480,N_5400);
nand U5682 (N_5682,N_5304,N_5405);
and U5683 (N_5683,N_5357,N_5335);
xnor U5684 (N_5684,N_5306,N_5361);
nor U5685 (N_5685,N_5309,N_5288);
or U5686 (N_5686,N_5261,N_5258);
nand U5687 (N_5687,N_5273,N_5275);
and U5688 (N_5688,N_5387,N_5350);
or U5689 (N_5689,N_5289,N_5365);
or U5690 (N_5690,N_5479,N_5353);
nor U5691 (N_5691,N_5252,N_5428);
or U5692 (N_5692,N_5383,N_5372);
nand U5693 (N_5693,N_5313,N_5466);
nand U5694 (N_5694,N_5323,N_5462);
and U5695 (N_5695,N_5490,N_5477);
and U5696 (N_5696,N_5287,N_5471);
xor U5697 (N_5697,N_5272,N_5386);
nor U5698 (N_5698,N_5257,N_5335);
or U5699 (N_5699,N_5346,N_5300);
nor U5700 (N_5700,N_5494,N_5323);
nor U5701 (N_5701,N_5338,N_5393);
and U5702 (N_5702,N_5464,N_5381);
and U5703 (N_5703,N_5267,N_5324);
nand U5704 (N_5704,N_5477,N_5340);
and U5705 (N_5705,N_5354,N_5308);
or U5706 (N_5706,N_5499,N_5378);
or U5707 (N_5707,N_5440,N_5493);
nand U5708 (N_5708,N_5272,N_5411);
nand U5709 (N_5709,N_5309,N_5429);
xnor U5710 (N_5710,N_5408,N_5388);
nand U5711 (N_5711,N_5463,N_5451);
nor U5712 (N_5712,N_5454,N_5260);
and U5713 (N_5713,N_5267,N_5454);
and U5714 (N_5714,N_5416,N_5320);
or U5715 (N_5715,N_5412,N_5312);
and U5716 (N_5716,N_5483,N_5368);
nor U5717 (N_5717,N_5477,N_5338);
and U5718 (N_5718,N_5407,N_5301);
or U5719 (N_5719,N_5435,N_5480);
xor U5720 (N_5720,N_5418,N_5445);
or U5721 (N_5721,N_5259,N_5353);
and U5722 (N_5722,N_5470,N_5299);
or U5723 (N_5723,N_5439,N_5409);
or U5724 (N_5724,N_5463,N_5361);
nand U5725 (N_5725,N_5410,N_5317);
xnor U5726 (N_5726,N_5424,N_5393);
nor U5727 (N_5727,N_5330,N_5378);
nand U5728 (N_5728,N_5326,N_5388);
nand U5729 (N_5729,N_5349,N_5414);
or U5730 (N_5730,N_5478,N_5340);
xor U5731 (N_5731,N_5306,N_5359);
nand U5732 (N_5732,N_5348,N_5444);
and U5733 (N_5733,N_5278,N_5282);
or U5734 (N_5734,N_5451,N_5268);
nor U5735 (N_5735,N_5305,N_5333);
nor U5736 (N_5736,N_5415,N_5360);
nor U5737 (N_5737,N_5320,N_5434);
nand U5738 (N_5738,N_5362,N_5361);
nand U5739 (N_5739,N_5269,N_5360);
or U5740 (N_5740,N_5459,N_5366);
or U5741 (N_5741,N_5410,N_5283);
or U5742 (N_5742,N_5366,N_5422);
nor U5743 (N_5743,N_5496,N_5419);
or U5744 (N_5744,N_5258,N_5439);
nand U5745 (N_5745,N_5472,N_5284);
or U5746 (N_5746,N_5405,N_5441);
or U5747 (N_5747,N_5364,N_5415);
nor U5748 (N_5748,N_5355,N_5497);
nand U5749 (N_5749,N_5482,N_5477);
nand U5750 (N_5750,N_5722,N_5683);
nand U5751 (N_5751,N_5573,N_5597);
or U5752 (N_5752,N_5625,N_5661);
and U5753 (N_5753,N_5679,N_5638);
nand U5754 (N_5754,N_5581,N_5596);
nor U5755 (N_5755,N_5739,N_5572);
nor U5756 (N_5756,N_5614,N_5673);
nor U5757 (N_5757,N_5512,N_5709);
xnor U5758 (N_5758,N_5632,N_5726);
nand U5759 (N_5759,N_5557,N_5667);
nor U5760 (N_5760,N_5730,N_5601);
or U5761 (N_5761,N_5708,N_5584);
nor U5762 (N_5762,N_5501,N_5513);
nand U5763 (N_5763,N_5594,N_5669);
nand U5764 (N_5764,N_5665,N_5509);
nor U5765 (N_5765,N_5619,N_5643);
and U5766 (N_5766,N_5518,N_5712);
nand U5767 (N_5767,N_5687,N_5651);
or U5768 (N_5768,N_5743,N_5727);
and U5769 (N_5769,N_5700,N_5617);
xor U5770 (N_5770,N_5503,N_5747);
nor U5771 (N_5771,N_5694,N_5566);
or U5772 (N_5772,N_5570,N_5689);
or U5773 (N_5773,N_5606,N_5721);
and U5774 (N_5774,N_5630,N_5642);
nand U5775 (N_5775,N_5541,N_5540);
nand U5776 (N_5776,N_5500,N_5682);
nor U5777 (N_5777,N_5582,N_5553);
nor U5778 (N_5778,N_5531,N_5530);
or U5779 (N_5779,N_5666,N_5748);
and U5780 (N_5780,N_5588,N_5529);
nor U5781 (N_5781,N_5519,N_5569);
nor U5782 (N_5782,N_5655,N_5567);
nand U5783 (N_5783,N_5662,N_5628);
or U5784 (N_5784,N_5670,N_5671);
or U5785 (N_5785,N_5631,N_5506);
nand U5786 (N_5786,N_5731,N_5647);
nor U5787 (N_5787,N_5608,N_5545);
nor U5788 (N_5788,N_5609,N_5741);
nand U5789 (N_5789,N_5677,N_5510);
nor U5790 (N_5790,N_5544,N_5734);
nor U5791 (N_5791,N_5688,N_5641);
nand U5792 (N_5792,N_5593,N_5524);
nor U5793 (N_5793,N_5615,N_5561);
or U5794 (N_5794,N_5652,N_5668);
and U5795 (N_5795,N_5595,N_5654);
nor U5796 (N_5796,N_5587,N_5728);
nor U5797 (N_5797,N_5681,N_5663);
and U5798 (N_5798,N_5556,N_5575);
or U5799 (N_5799,N_5613,N_5550);
and U5800 (N_5800,N_5563,N_5580);
or U5801 (N_5801,N_5622,N_5571);
nor U5802 (N_5802,N_5577,N_5644);
nand U5803 (N_5803,N_5589,N_5514);
nand U5804 (N_5804,N_5618,N_5583);
and U5805 (N_5805,N_5605,N_5505);
nand U5806 (N_5806,N_5711,N_5650);
nor U5807 (N_5807,N_5659,N_5626);
nand U5808 (N_5808,N_5685,N_5559);
nand U5809 (N_5809,N_5610,N_5525);
and U5810 (N_5810,N_5522,N_5627);
nor U5811 (N_5811,N_5736,N_5724);
and U5812 (N_5812,N_5542,N_5749);
and U5813 (N_5813,N_5612,N_5723);
and U5814 (N_5814,N_5735,N_5534);
nor U5815 (N_5815,N_5558,N_5701);
nor U5816 (N_5816,N_5546,N_5591);
and U5817 (N_5817,N_5664,N_5649);
or U5818 (N_5818,N_5656,N_5692);
and U5819 (N_5819,N_5674,N_5725);
nor U5820 (N_5820,N_5599,N_5699);
or U5821 (N_5821,N_5660,N_5547);
or U5822 (N_5822,N_5634,N_5537);
nand U5823 (N_5823,N_5719,N_5629);
and U5824 (N_5824,N_5675,N_5740);
or U5825 (N_5825,N_5718,N_5729);
nor U5826 (N_5826,N_5707,N_5502);
or U5827 (N_5827,N_5635,N_5691);
and U5828 (N_5828,N_5680,N_5744);
nor U5829 (N_5829,N_5678,N_5543);
and U5830 (N_5830,N_5578,N_5536);
and U5831 (N_5831,N_5602,N_5598);
nand U5832 (N_5832,N_5604,N_5693);
and U5833 (N_5833,N_5672,N_5697);
nand U5834 (N_5834,N_5703,N_5551);
nand U5835 (N_5835,N_5562,N_5516);
and U5836 (N_5836,N_5515,N_5676);
nor U5837 (N_5837,N_5716,N_5704);
nand U5838 (N_5838,N_5527,N_5538);
and U5839 (N_5839,N_5633,N_5742);
or U5840 (N_5840,N_5623,N_5560);
and U5841 (N_5841,N_5745,N_5520);
or U5842 (N_5842,N_5523,N_5713);
or U5843 (N_5843,N_5600,N_5717);
nor U5844 (N_5844,N_5698,N_5504);
and U5845 (N_5845,N_5620,N_5535);
or U5846 (N_5846,N_5646,N_5616);
or U5847 (N_5847,N_5579,N_5702);
and U5848 (N_5848,N_5548,N_5684);
nor U5849 (N_5849,N_5576,N_5732);
nor U5850 (N_5850,N_5710,N_5657);
nand U5851 (N_5851,N_5720,N_5621);
or U5852 (N_5852,N_5738,N_5554);
and U5853 (N_5853,N_5528,N_5636);
or U5854 (N_5854,N_5696,N_5586);
or U5855 (N_5855,N_5607,N_5549);
nor U5856 (N_5856,N_5508,N_5611);
or U5857 (N_5857,N_5564,N_5690);
nor U5858 (N_5858,N_5714,N_5658);
and U5859 (N_5859,N_5624,N_5695);
or U5860 (N_5860,N_5737,N_5590);
nand U5861 (N_5861,N_5592,N_5511);
nor U5862 (N_5862,N_5640,N_5648);
or U5863 (N_5863,N_5733,N_5565);
and U5864 (N_5864,N_5539,N_5532);
or U5865 (N_5865,N_5507,N_5706);
nor U5866 (N_5866,N_5603,N_5746);
nand U5867 (N_5867,N_5585,N_5555);
nor U5868 (N_5868,N_5526,N_5533);
and U5869 (N_5869,N_5568,N_5574);
xnor U5870 (N_5870,N_5521,N_5653);
or U5871 (N_5871,N_5705,N_5552);
or U5872 (N_5872,N_5637,N_5639);
nor U5873 (N_5873,N_5715,N_5686);
or U5874 (N_5874,N_5645,N_5517);
nand U5875 (N_5875,N_5688,N_5646);
or U5876 (N_5876,N_5550,N_5611);
or U5877 (N_5877,N_5594,N_5681);
or U5878 (N_5878,N_5628,N_5684);
nor U5879 (N_5879,N_5746,N_5513);
nor U5880 (N_5880,N_5741,N_5500);
nor U5881 (N_5881,N_5581,N_5636);
or U5882 (N_5882,N_5538,N_5555);
or U5883 (N_5883,N_5509,N_5519);
nor U5884 (N_5884,N_5728,N_5637);
nand U5885 (N_5885,N_5667,N_5716);
xnor U5886 (N_5886,N_5562,N_5549);
and U5887 (N_5887,N_5684,N_5691);
and U5888 (N_5888,N_5676,N_5690);
and U5889 (N_5889,N_5583,N_5670);
nor U5890 (N_5890,N_5618,N_5616);
or U5891 (N_5891,N_5627,N_5716);
nand U5892 (N_5892,N_5676,N_5662);
or U5893 (N_5893,N_5629,N_5526);
or U5894 (N_5894,N_5715,N_5548);
or U5895 (N_5895,N_5633,N_5638);
nand U5896 (N_5896,N_5507,N_5623);
and U5897 (N_5897,N_5525,N_5593);
nor U5898 (N_5898,N_5521,N_5593);
nand U5899 (N_5899,N_5645,N_5557);
nand U5900 (N_5900,N_5687,N_5705);
or U5901 (N_5901,N_5654,N_5569);
xnor U5902 (N_5902,N_5732,N_5598);
nor U5903 (N_5903,N_5571,N_5680);
nor U5904 (N_5904,N_5700,N_5542);
and U5905 (N_5905,N_5711,N_5661);
nor U5906 (N_5906,N_5528,N_5682);
nor U5907 (N_5907,N_5588,N_5591);
or U5908 (N_5908,N_5667,N_5738);
nor U5909 (N_5909,N_5526,N_5580);
nand U5910 (N_5910,N_5560,N_5739);
and U5911 (N_5911,N_5714,N_5746);
or U5912 (N_5912,N_5524,N_5692);
xnor U5913 (N_5913,N_5586,N_5610);
nor U5914 (N_5914,N_5518,N_5574);
nand U5915 (N_5915,N_5503,N_5712);
nand U5916 (N_5916,N_5655,N_5658);
nand U5917 (N_5917,N_5520,N_5514);
nand U5918 (N_5918,N_5732,N_5604);
or U5919 (N_5919,N_5558,N_5538);
nand U5920 (N_5920,N_5502,N_5666);
or U5921 (N_5921,N_5682,N_5573);
nand U5922 (N_5922,N_5617,N_5534);
nand U5923 (N_5923,N_5597,N_5696);
or U5924 (N_5924,N_5529,N_5700);
nand U5925 (N_5925,N_5542,N_5546);
or U5926 (N_5926,N_5551,N_5643);
and U5927 (N_5927,N_5685,N_5627);
and U5928 (N_5928,N_5653,N_5685);
nor U5929 (N_5929,N_5519,N_5506);
nor U5930 (N_5930,N_5597,N_5644);
and U5931 (N_5931,N_5546,N_5513);
or U5932 (N_5932,N_5610,N_5744);
nor U5933 (N_5933,N_5697,N_5688);
or U5934 (N_5934,N_5558,N_5678);
or U5935 (N_5935,N_5671,N_5673);
nor U5936 (N_5936,N_5659,N_5643);
xnor U5937 (N_5937,N_5608,N_5519);
nand U5938 (N_5938,N_5696,N_5562);
nand U5939 (N_5939,N_5595,N_5600);
and U5940 (N_5940,N_5629,N_5663);
nor U5941 (N_5941,N_5683,N_5521);
and U5942 (N_5942,N_5598,N_5518);
or U5943 (N_5943,N_5671,N_5550);
nor U5944 (N_5944,N_5529,N_5681);
or U5945 (N_5945,N_5650,N_5554);
nor U5946 (N_5946,N_5529,N_5713);
nor U5947 (N_5947,N_5520,N_5712);
or U5948 (N_5948,N_5532,N_5660);
nor U5949 (N_5949,N_5670,N_5504);
and U5950 (N_5950,N_5699,N_5638);
and U5951 (N_5951,N_5624,N_5544);
nand U5952 (N_5952,N_5511,N_5602);
nor U5953 (N_5953,N_5574,N_5519);
and U5954 (N_5954,N_5714,N_5560);
and U5955 (N_5955,N_5722,N_5567);
or U5956 (N_5956,N_5667,N_5563);
nand U5957 (N_5957,N_5652,N_5611);
or U5958 (N_5958,N_5502,N_5505);
nand U5959 (N_5959,N_5617,N_5631);
or U5960 (N_5960,N_5549,N_5610);
and U5961 (N_5961,N_5640,N_5711);
nor U5962 (N_5962,N_5711,N_5714);
nor U5963 (N_5963,N_5600,N_5700);
and U5964 (N_5964,N_5643,N_5662);
and U5965 (N_5965,N_5614,N_5583);
or U5966 (N_5966,N_5617,N_5648);
and U5967 (N_5967,N_5553,N_5665);
nor U5968 (N_5968,N_5593,N_5594);
nor U5969 (N_5969,N_5708,N_5611);
nor U5970 (N_5970,N_5571,N_5528);
nand U5971 (N_5971,N_5622,N_5573);
nor U5972 (N_5972,N_5663,N_5704);
and U5973 (N_5973,N_5527,N_5521);
or U5974 (N_5974,N_5540,N_5573);
nand U5975 (N_5975,N_5603,N_5744);
and U5976 (N_5976,N_5731,N_5561);
nor U5977 (N_5977,N_5719,N_5525);
or U5978 (N_5978,N_5671,N_5646);
and U5979 (N_5979,N_5718,N_5691);
nand U5980 (N_5980,N_5746,N_5699);
and U5981 (N_5981,N_5632,N_5714);
nor U5982 (N_5982,N_5554,N_5593);
and U5983 (N_5983,N_5733,N_5578);
nor U5984 (N_5984,N_5589,N_5515);
nand U5985 (N_5985,N_5745,N_5536);
xnor U5986 (N_5986,N_5561,N_5676);
and U5987 (N_5987,N_5724,N_5519);
nand U5988 (N_5988,N_5635,N_5682);
nor U5989 (N_5989,N_5581,N_5727);
or U5990 (N_5990,N_5745,N_5655);
and U5991 (N_5991,N_5746,N_5560);
or U5992 (N_5992,N_5697,N_5626);
nand U5993 (N_5993,N_5589,N_5575);
nand U5994 (N_5994,N_5700,N_5512);
and U5995 (N_5995,N_5676,N_5708);
nor U5996 (N_5996,N_5579,N_5713);
and U5997 (N_5997,N_5706,N_5665);
and U5998 (N_5998,N_5581,N_5512);
and U5999 (N_5999,N_5524,N_5520);
nor U6000 (N_6000,N_5783,N_5913);
or U6001 (N_6001,N_5983,N_5961);
or U6002 (N_6002,N_5832,N_5933);
nor U6003 (N_6003,N_5819,N_5801);
and U6004 (N_6004,N_5874,N_5849);
nand U6005 (N_6005,N_5804,N_5791);
and U6006 (N_6006,N_5784,N_5937);
nand U6007 (N_6007,N_5993,N_5864);
nor U6008 (N_6008,N_5788,N_5778);
and U6009 (N_6009,N_5988,N_5807);
and U6010 (N_6010,N_5960,N_5934);
nand U6011 (N_6011,N_5941,N_5894);
nor U6012 (N_6012,N_5827,N_5877);
nor U6013 (N_6013,N_5981,N_5906);
and U6014 (N_6014,N_5978,N_5859);
nand U6015 (N_6015,N_5964,N_5817);
and U6016 (N_6016,N_5890,N_5947);
nand U6017 (N_6017,N_5892,N_5997);
nand U6018 (N_6018,N_5850,N_5806);
or U6019 (N_6019,N_5863,N_5833);
and U6020 (N_6020,N_5875,N_5840);
or U6021 (N_6021,N_5949,N_5766);
and U6022 (N_6022,N_5810,N_5761);
or U6023 (N_6023,N_5758,N_5882);
or U6024 (N_6024,N_5835,N_5975);
or U6025 (N_6025,N_5816,N_5929);
and U6026 (N_6026,N_5914,N_5879);
nand U6027 (N_6027,N_5809,N_5823);
nand U6028 (N_6028,N_5812,N_5769);
nand U6029 (N_6029,N_5869,N_5985);
or U6030 (N_6030,N_5773,N_5899);
and U6031 (N_6031,N_5786,N_5854);
or U6032 (N_6032,N_5943,N_5918);
or U6033 (N_6033,N_5953,N_5866);
xor U6034 (N_6034,N_5963,N_5842);
or U6035 (N_6035,N_5768,N_5995);
and U6036 (N_6036,N_5930,N_5803);
nor U6037 (N_6037,N_5822,N_5886);
or U6038 (N_6038,N_5779,N_5767);
nand U6039 (N_6039,N_5878,N_5826);
and U6040 (N_6040,N_5919,N_5861);
nor U6041 (N_6041,N_5813,N_5972);
nor U6042 (N_6042,N_5772,N_5956);
or U6043 (N_6043,N_5920,N_5948);
nand U6044 (N_6044,N_5962,N_5828);
nand U6045 (N_6045,N_5935,N_5764);
nand U6046 (N_6046,N_5959,N_5876);
nor U6047 (N_6047,N_5977,N_5910);
nor U6048 (N_6048,N_5916,N_5844);
nor U6049 (N_6049,N_5846,N_5752);
and U6050 (N_6050,N_5946,N_5834);
and U6051 (N_6051,N_5904,N_5777);
nand U6052 (N_6052,N_5982,N_5903);
nor U6053 (N_6053,N_5802,N_5986);
nand U6054 (N_6054,N_5887,N_5763);
nor U6055 (N_6055,N_5818,N_5765);
or U6056 (N_6056,N_5987,N_5790);
or U6057 (N_6057,N_5808,N_5858);
nor U6058 (N_6058,N_5824,N_5780);
nand U6059 (N_6059,N_5900,N_5957);
or U6060 (N_6060,N_5944,N_5925);
nand U6061 (N_6061,N_5781,N_5831);
nor U6062 (N_6062,N_5966,N_5893);
or U6063 (N_6063,N_5760,N_5862);
nor U6064 (N_6064,N_5901,N_5774);
and U6065 (N_6065,N_5942,N_5787);
nor U6066 (N_6066,N_5751,N_5830);
or U6067 (N_6067,N_5821,N_5841);
and U6068 (N_6068,N_5902,N_5847);
xnor U6069 (N_6069,N_5915,N_5815);
or U6070 (N_6070,N_5825,N_5928);
nor U6071 (N_6071,N_5958,N_5990);
nand U6072 (N_6072,N_5836,N_5911);
or U6073 (N_6073,N_5852,N_5843);
or U6074 (N_6074,N_5857,N_5923);
or U6075 (N_6075,N_5955,N_5938);
nand U6076 (N_6076,N_5888,N_5873);
nand U6077 (N_6077,N_5771,N_5896);
nor U6078 (N_6078,N_5980,N_5907);
and U6079 (N_6079,N_5940,N_5932);
or U6080 (N_6080,N_5922,N_5994);
nand U6081 (N_6081,N_5754,N_5908);
nand U6082 (N_6082,N_5762,N_5883);
and U6083 (N_6083,N_5973,N_5820);
and U6084 (N_6084,N_5775,N_5970);
nor U6085 (N_6085,N_5889,N_5897);
nor U6086 (N_6086,N_5891,N_5884);
nand U6087 (N_6087,N_5931,N_5989);
or U6088 (N_6088,N_5998,N_5755);
or U6089 (N_6089,N_5976,N_5789);
and U6090 (N_6090,N_5881,N_5872);
or U6091 (N_6091,N_5839,N_5776);
nand U6092 (N_6092,N_5950,N_5793);
and U6093 (N_6093,N_5848,N_5871);
nor U6094 (N_6094,N_5856,N_5805);
nand U6095 (N_6095,N_5853,N_5792);
and U6096 (N_6096,N_5984,N_5860);
and U6097 (N_6097,N_5867,N_5814);
nor U6098 (N_6098,N_5799,N_5905);
nor U6099 (N_6099,N_5855,N_5979);
nor U6100 (N_6100,N_5895,N_5991);
nor U6101 (N_6101,N_5999,N_5927);
or U6102 (N_6102,N_5885,N_5909);
nand U6103 (N_6103,N_5796,N_5870);
and U6104 (N_6104,N_5936,N_5757);
and U6105 (N_6105,N_5912,N_5969);
nor U6106 (N_6106,N_5794,N_5880);
or U6107 (N_6107,N_5797,N_5945);
and U6108 (N_6108,N_5838,N_5750);
nand U6109 (N_6109,N_5954,N_5926);
nor U6110 (N_6110,N_5800,N_5837);
and U6111 (N_6111,N_5898,N_5756);
nand U6112 (N_6112,N_5996,N_5951);
and U6113 (N_6113,N_5939,N_5917);
nor U6114 (N_6114,N_5952,N_5753);
and U6115 (N_6115,N_5967,N_5924);
or U6116 (N_6116,N_5845,N_5851);
nand U6117 (N_6117,N_5770,N_5971);
nor U6118 (N_6118,N_5795,N_5868);
and U6119 (N_6119,N_5992,N_5974);
and U6120 (N_6120,N_5921,N_5785);
nand U6121 (N_6121,N_5965,N_5865);
or U6122 (N_6122,N_5759,N_5968);
or U6123 (N_6123,N_5798,N_5811);
nor U6124 (N_6124,N_5829,N_5782);
xor U6125 (N_6125,N_5867,N_5863);
or U6126 (N_6126,N_5935,N_5840);
or U6127 (N_6127,N_5983,N_5974);
xnor U6128 (N_6128,N_5938,N_5868);
nand U6129 (N_6129,N_5980,N_5874);
nor U6130 (N_6130,N_5918,N_5941);
nand U6131 (N_6131,N_5803,N_5883);
and U6132 (N_6132,N_5888,N_5810);
nor U6133 (N_6133,N_5859,N_5814);
or U6134 (N_6134,N_5772,N_5892);
and U6135 (N_6135,N_5864,N_5833);
nor U6136 (N_6136,N_5833,N_5781);
and U6137 (N_6137,N_5980,N_5900);
nor U6138 (N_6138,N_5752,N_5754);
or U6139 (N_6139,N_5757,N_5985);
nor U6140 (N_6140,N_5969,N_5944);
nand U6141 (N_6141,N_5770,N_5968);
nor U6142 (N_6142,N_5914,N_5934);
or U6143 (N_6143,N_5995,N_5799);
and U6144 (N_6144,N_5903,N_5937);
nand U6145 (N_6145,N_5978,N_5789);
nor U6146 (N_6146,N_5788,N_5777);
nand U6147 (N_6147,N_5759,N_5947);
nor U6148 (N_6148,N_5763,N_5878);
and U6149 (N_6149,N_5968,N_5863);
nor U6150 (N_6150,N_5955,N_5859);
nand U6151 (N_6151,N_5755,N_5786);
nor U6152 (N_6152,N_5902,N_5873);
nand U6153 (N_6153,N_5833,N_5912);
nand U6154 (N_6154,N_5996,N_5946);
or U6155 (N_6155,N_5985,N_5961);
nand U6156 (N_6156,N_5909,N_5898);
or U6157 (N_6157,N_5972,N_5971);
xnor U6158 (N_6158,N_5826,N_5839);
nand U6159 (N_6159,N_5791,N_5820);
nand U6160 (N_6160,N_5886,N_5922);
and U6161 (N_6161,N_5805,N_5751);
nand U6162 (N_6162,N_5857,N_5866);
or U6163 (N_6163,N_5815,N_5808);
or U6164 (N_6164,N_5852,N_5847);
and U6165 (N_6165,N_5949,N_5859);
nor U6166 (N_6166,N_5858,N_5977);
or U6167 (N_6167,N_5989,N_5782);
nand U6168 (N_6168,N_5753,N_5805);
nor U6169 (N_6169,N_5750,N_5975);
nor U6170 (N_6170,N_5982,N_5975);
and U6171 (N_6171,N_5777,N_5871);
nand U6172 (N_6172,N_5872,N_5996);
and U6173 (N_6173,N_5968,N_5980);
nand U6174 (N_6174,N_5991,N_5778);
xnor U6175 (N_6175,N_5979,N_5765);
nor U6176 (N_6176,N_5932,N_5918);
or U6177 (N_6177,N_5758,N_5892);
and U6178 (N_6178,N_5874,N_5968);
nor U6179 (N_6179,N_5865,N_5812);
or U6180 (N_6180,N_5936,N_5754);
or U6181 (N_6181,N_5841,N_5963);
and U6182 (N_6182,N_5809,N_5759);
nand U6183 (N_6183,N_5802,N_5872);
nor U6184 (N_6184,N_5938,N_5923);
nor U6185 (N_6185,N_5938,N_5895);
nand U6186 (N_6186,N_5843,N_5819);
nand U6187 (N_6187,N_5873,N_5939);
nand U6188 (N_6188,N_5889,N_5886);
nand U6189 (N_6189,N_5850,N_5907);
nor U6190 (N_6190,N_5808,N_5900);
nor U6191 (N_6191,N_5951,N_5810);
or U6192 (N_6192,N_5821,N_5790);
nor U6193 (N_6193,N_5916,N_5823);
or U6194 (N_6194,N_5754,N_5900);
or U6195 (N_6195,N_5979,N_5948);
and U6196 (N_6196,N_5900,N_5994);
and U6197 (N_6197,N_5871,N_5837);
and U6198 (N_6198,N_5873,N_5931);
and U6199 (N_6199,N_5898,N_5929);
or U6200 (N_6200,N_5840,N_5859);
nor U6201 (N_6201,N_5799,N_5992);
nand U6202 (N_6202,N_5873,N_5954);
nor U6203 (N_6203,N_5990,N_5859);
and U6204 (N_6204,N_5927,N_5773);
and U6205 (N_6205,N_5946,N_5985);
or U6206 (N_6206,N_5755,N_5763);
or U6207 (N_6207,N_5762,N_5946);
or U6208 (N_6208,N_5822,N_5878);
nand U6209 (N_6209,N_5753,N_5951);
nor U6210 (N_6210,N_5769,N_5800);
nand U6211 (N_6211,N_5828,N_5931);
and U6212 (N_6212,N_5942,N_5753);
and U6213 (N_6213,N_5986,N_5818);
and U6214 (N_6214,N_5856,N_5774);
nand U6215 (N_6215,N_5801,N_5982);
nand U6216 (N_6216,N_5750,N_5878);
or U6217 (N_6217,N_5965,N_5952);
xor U6218 (N_6218,N_5814,N_5863);
nand U6219 (N_6219,N_5841,N_5851);
xnor U6220 (N_6220,N_5947,N_5839);
or U6221 (N_6221,N_5991,N_5983);
nor U6222 (N_6222,N_5996,N_5805);
nand U6223 (N_6223,N_5836,N_5975);
and U6224 (N_6224,N_5937,N_5928);
nor U6225 (N_6225,N_5920,N_5833);
or U6226 (N_6226,N_5799,N_5873);
nor U6227 (N_6227,N_5761,N_5883);
nor U6228 (N_6228,N_5813,N_5960);
nand U6229 (N_6229,N_5825,N_5843);
and U6230 (N_6230,N_5815,N_5947);
or U6231 (N_6231,N_5945,N_5939);
nor U6232 (N_6232,N_5753,N_5807);
nand U6233 (N_6233,N_5911,N_5951);
and U6234 (N_6234,N_5870,N_5830);
nand U6235 (N_6235,N_5905,N_5755);
and U6236 (N_6236,N_5815,N_5764);
and U6237 (N_6237,N_5862,N_5823);
or U6238 (N_6238,N_5774,N_5954);
nand U6239 (N_6239,N_5886,N_5910);
or U6240 (N_6240,N_5948,N_5917);
and U6241 (N_6241,N_5928,N_5809);
or U6242 (N_6242,N_5982,N_5913);
nor U6243 (N_6243,N_5964,N_5810);
nor U6244 (N_6244,N_5915,N_5979);
nor U6245 (N_6245,N_5878,N_5949);
nor U6246 (N_6246,N_5833,N_5962);
or U6247 (N_6247,N_5997,N_5844);
and U6248 (N_6248,N_5751,N_5975);
and U6249 (N_6249,N_5946,N_5866);
nor U6250 (N_6250,N_6230,N_6120);
nand U6251 (N_6251,N_6071,N_6238);
and U6252 (N_6252,N_6186,N_6132);
and U6253 (N_6253,N_6170,N_6050);
nand U6254 (N_6254,N_6061,N_6097);
nand U6255 (N_6255,N_6072,N_6003);
and U6256 (N_6256,N_6048,N_6029);
or U6257 (N_6257,N_6066,N_6176);
xor U6258 (N_6258,N_6147,N_6167);
nand U6259 (N_6259,N_6156,N_6245);
xnor U6260 (N_6260,N_6084,N_6222);
nor U6261 (N_6261,N_6031,N_6127);
nand U6262 (N_6262,N_6190,N_6121);
nand U6263 (N_6263,N_6145,N_6104);
or U6264 (N_6264,N_6129,N_6049);
nand U6265 (N_6265,N_6064,N_6028);
nand U6266 (N_6266,N_6098,N_6125);
or U6267 (N_6267,N_6198,N_6158);
nand U6268 (N_6268,N_6200,N_6201);
and U6269 (N_6269,N_6134,N_6149);
nor U6270 (N_6270,N_6012,N_6192);
nor U6271 (N_6271,N_6101,N_6246);
nand U6272 (N_6272,N_6093,N_6067);
nand U6273 (N_6273,N_6089,N_6039);
and U6274 (N_6274,N_6138,N_6148);
and U6275 (N_6275,N_6209,N_6207);
or U6276 (N_6276,N_6194,N_6117);
nand U6277 (N_6277,N_6103,N_6030);
xor U6278 (N_6278,N_6151,N_6159);
nand U6279 (N_6279,N_6100,N_6063);
or U6280 (N_6280,N_6099,N_6218);
nand U6281 (N_6281,N_6140,N_6017);
xor U6282 (N_6282,N_6062,N_6105);
or U6283 (N_6283,N_6199,N_6080);
xnor U6284 (N_6284,N_6183,N_6113);
or U6285 (N_6285,N_6070,N_6131);
nor U6286 (N_6286,N_6024,N_6051);
nor U6287 (N_6287,N_6095,N_6092);
or U6288 (N_6288,N_6204,N_6075);
nor U6289 (N_6289,N_6189,N_6032);
nand U6290 (N_6290,N_6009,N_6136);
or U6291 (N_6291,N_6087,N_6079);
nor U6292 (N_6292,N_6005,N_6130);
and U6293 (N_6293,N_6135,N_6122);
or U6294 (N_6294,N_6053,N_6011);
and U6295 (N_6295,N_6019,N_6241);
nand U6296 (N_6296,N_6188,N_6180);
nand U6297 (N_6297,N_6239,N_6077);
nand U6298 (N_6298,N_6018,N_6133);
nor U6299 (N_6299,N_6119,N_6060);
and U6300 (N_6300,N_6074,N_6193);
nor U6301 (N_6301,N_6157,N_6016);
or U6302 (N_6302,N_6088,N_6248);
or U6303 (N_6303,N_6237,N_6171);
nand U6304 (N_6304,N_6034,N_6173);
or U6305 (N_6305,N_6083,N_6006);
and U6306 (N_6306,N_6056,N_6211);
or U6307 (N_6307,N_6205,N_6219);
nor U6308 (N_6308,N_6021,N_6227);
and U6309 (N_6309,N_6187,N_6141);
and U6310 (N_6310,N_6114,N_6115);
and U6311 (N_6311,N_6078,N_6178);
nand U6312 (N_6312,N_6073,N_6068);
nand U6313 (N_6313,N_6181,N_6226);
nor U6314 (N_6314,N_6144,N_6242);
or U6315 (N_6315,N_6228,N_6065);
nor U6316 (N_6316,N_6054,N_6111);
nand U6317 (N_6317,N_6164,N_6212);
or U6318 (N_6318,N_6220,N_6015);
nor U6319 (N_6319,N_6243,N_6094);
nand U6320 (N_6320,N_6000,N_6214);
or U6321 (N_6321,N_6076,N_6184);
and U6322 (N_6322,N_6169,N_6043);
nand U6323 (N_6323,N_6247,N_6107);
nand U6324 (N_6324,N_6161,N_6160);
xor U6325 (N_6325,N_6202,N_6213);
nor U6326 (N_6326,N_6059,N_6231);
or U6327 (N_6327,N_6223,N_6081);
nand U6328 (N_6328,N_6042,N_6152);
nand U6329 (N_6329,N_6150,N_6110);
nand U6330 (N_6330,N_6037,N_6045);
nor U6331 (N_6331,N_6052,N_6002);
and U6332 (N_6332,N_6069,N_6154);
or U6333 (N_6333,N_6162,N_6046);
and U6334 (N_6334,N_6109,N_6102);
nand U6335 (N_6335,N_6010,N_6038);
nor U6336 (N_6336,N_6143,N_6208);
or U6337 (N_6337,N_6118,N_6007);
nor U6338 (N_6338,N_6085,N_6196);
and U6339 (N_6339,N_6036,N_6232);
nor U6340 (N_6340,N_6179,N_6197);
and U6341 (N_6341,N_6026,N_6240);
nand U6342 (N_6342,N_6155,N_6008);
and U6343 (N_6343,N_6233,N_6004);
and U6344 (N_6344,N_6022,N_6027);
or U6345 (N_6345,N_6082,N_6203);
nand U6346 (N_6346,N_6035,N_6221);
nor U6347 (N_6347,N_6216,N_6055);
or U6348 (N_6348,N_6025,N_6236);
or U6349 (N_6349,N_6210,N_6124);
and U6350 (N_6350,N_6168,N_6139);
and U6351 (N_6351,N_6153,N_6185);
and U6352 (N_6352,N_6225,N_6195);
and U6353 (N_6353,N_6234,N_6172);
and U6354 (N_6354,N_6116,N_6041);
and U6355 (N_6355,N_6126,N_6174);
and U6356 (N_6356,N_6137,N_6108);
or U6357 (N_6357,N_6001,N_6175);
and U6358 (N_6358,N_6014,N_6229);
xor U6359 (N_6359,N_6040,N_6191);
and U6360 (N_6360,N_6106,N_6112);
nor U6361 (N_6361,N_6182,N_6146);
nor U6362 (N_6362,N_6224,N_6090);
nand U6363 (N_6363,N_6235,N_6163);
and U6364 (N_6364,N_6217,N_6086);
nand U6365 (N_6365,N_6215,N_6177);
nand U6366 (N_6366,N_6249,N_6023);
xnor U6367 (N_6367,N_6044,N_6166);
nor U6368 (N_6368,N_6165,N_6058);
nand U6369 (N_6369,N_6047,N_6142);
nand U6370 (N_6370,N_6244,N_6020);
nand U6371 (N_6371,N_6057,N_6123);
nand U6372 (N_6372,N_6096,N_6091);
and U6373 (N_6373,N_6013,N_6033);
and U6374 (N_6374,N_6128,N_6206);
and U6375 (N_6375,N_6122,N_6235);
nor U6376 (N_6376,N_6079,N_6033);
nor U6377 (N_6377,N_6147,N_6060);
or U6378 (N_6378,N_6078,N_6127);
nand U6379 (N_6379,N_6102,N_6096);
and U6380 (N_6380,N_6097,N_6090);
and U6381 (N_6381,N_6191,N_6209);
or U6382 (N_6382,N_6128,N_6058);
nand U6383 (N_6383,N_6209,N_6224);
nand U6384 (N_6384,N_6181,N_6238);
or U6385 (N_6385,N_6227,N_6096);
nor U6386 (N_6386,N_6159,N_6004);
nand U6387 (N_6387,N_6133,N_6084);
or U6388 (N_6388,N_6243,N_6005);
and U6389 (N_6389,N_6000,N_6205);
nand U6390 (N_6390,N_6159,N_6209);
and U6391 (N_6391,N_6097,N_6207);
nand U6392 (N_6392,N_6045,N_6083);
nor U6393 (N_6393,N_6068,N_6198);
nand U6394 (N_6394,N_6030,N_6167);
nor U6395 (N_6395,N_6168,N_6190);
or U6396 (N_6396,N_6103,N_6057);
or U6397 (N_6397,N_6237,N_6189);
nor U6398 (N_6398,N_6137,N_6176);
or U6399 (N_6399,N_6124,N_6185);
or U6400 (N_6400,N_6140,N_6133);
or U6401 (N_6401,N_6147,N_6009);
nand U6402 (N_6402,N_6070,N_6191);
and U6403 (N_6403,N_6035,N_6030);
nand U6404 (N_6404,N_6063,N_6218);
nand U6405 (N_6405,N_6035,N_6052);
or U6406 (N_6406,N_6159,N_6227);
nand U6407 (N_6407,N_6190,N_6098);
nor U6408 (N_6408,N_6123,N_6172);
and U6409 (N_6409,N_6155,N_6184);
and U6410 (N_6410,N_6085,N_6088);
nor U6411 (N_6411,N_6071,N_6069);
or U6412 (N_6412,N_6025,N_6168);
or U6413 (N_6413,N_6166,N_6026);
and U6414 (N_6414,N_6245,N_6018);
nand U6415 (N_6415,N_6104,N_6095);
nand U6416 (N_6416,N_6058,N_6211);
nor U6417 (N_6417,N_6126,N_6191);
nand U6418 (N_6418,N_6127,N_6147);
and U6419 (N_6419,N_6215,N_6165);
or U6420 (N_6420,N_6114,N_6069);
or U6421 (N_6421,N_6013,N_6105);
nand U6422 (N_6422,N_6144,N_6095);
and U6423 (N_6423,N_6173,N_6094);
or U6424 (N_6424,N_6025,N_6046);
nor U6425 (N_6425,N_6193,N_6220);
xnor U6426 (N_6426,N_6108,N_6070);
nand U6427 (N_6427,N_6004,N_6236);
nand U6428 (N_6428,N_6128,N_6111);
nor U6429 (N_6429,N_6000,N_6073);
nor U6430 (N_6430,N_6223,N_6050);
nor U6431 (N_6431,N_6017,N_6175);
nor U6432 (N_6432,N_6157,N_6239);
or U6433 (N_6433,N_6126,N_6185);
or U6434 (N_6434,N_6039,N_6166);
nor U6435 (N_6435,N_6133,N_6022);
or U6436 (N_6436,N_6166,N_6004);
xor U6437 (N_6437,N_6033,N_6138);
nor U6438 (N_6438,N_6024,N_6203);
nand U6439 (N_6439,N_6004,N_6229);
nand U6440 (N_6440,N_6001,N_6022);
nor U6441 (N_6441,N_6020,N_6017);
and U6442 (N_6442,N_6192,N_6116);
or U6443 (N_6443,N_6216,N_6021);
or U6444 (N_6444,N_6163,N_6013);
or U6445 (N_6445,N_6062,N_6090);
nor U6446 (N_6446,N_6191,N_6233);
or U6447 (N_6447,N_6147,N_6244);
and U6448 (N_6448,N_6068,N_6085);
or U6449 (N_6449,N_6076,N_6122);
nor U6450 (N_6450,N_6238,N_6151);
and U6451 (N_6451,N_6113,N_6050);
and U6452 (N_6452,N_6172,N_6129);
or U6453 (N_6453,N_6056,N_6054);
and U6454 (N_6454,N_6036,N_6038);
nand U6455 (N_6455,N_6016,N_6060);
and U6456 (N_6456,N_6067,N_6234);
nor U6457 (N_6457,N_6012,N_6014);
nand U6458 (N_6458,N_6152,N_6001);
nor U6459 (N_6459,N_6019,N_6209);
and U6460 (N_6460,N_6142,N_6073);
nor U6461 (N_6461,N_6099,N_6163);
nand U6462 (N_6462,N_6152,N_6157);
and U6463 (N_6463,N_6064,N_6117);
nand U6464 (N_6464,N_6131,N_6029);
nor U6465 (N_6465,N_6185,N_6201);
nand U6466 (N_6466,N_6179,N_6065);
and U6467 (N_6467,N_6096,N_6110);
nand U6468 (N_6468,N_6175,N_6224);
nor U6469 (N_6469,N_6041,N_6082);
and U6470 (N_6470,N_6187,N_6183);
or U6471 (N_6471,N_6008,N_6119);
and U6472 (N_6472,N_6196,N_6090);
nor U6473 (N_6473,N_6188,N_6101);
or U6474 (N_6474,N_6163,N_6181);
and U6475 (N_6475,N_6148,N_6185);
nand U6476 (N_6476,N_6164,N_6170);
or U6477 (N_6477,N_6143,N_6135);
nand U6478 (N_6478,N_6114,N_6202);
and U6479 (N_6479,N_6016,N_6119);
or U6480 (N_6480,N_6072,N_6191);
nor U6481 (N_6481,N_6070,N_6061);
or U6482 (N_6482,N_6175,N_6220);
and U6483 (N_6483,N_6240,N_6245);
or U6484 (N_6484,N_6204,N_6248);
nor U6485 (N_6485,N_6205,N_6119);
or U6486 (N_6486,N_6246,N_6083);
and U6487 (N_6487,N_6225,N_6047);
and U6488 (N_6488,N_6050,N_6192);
nor U6489 (N_6489,N_6010,N_6160);
nand U6490 (N_6490,N_6241,N_6080);
and U6491 (N_6491,N_6015,N_6108);
nor U6492 (N_6492,N_6218,N_6157);
nor U6493 (N_6493,N_6216,N_6205);
nor U6494 (N_6494,N_6009,N_6241);
nand U6495 (N_6495,N_6138,N_6107);
or U6496 (N_6496,N_6050,N_6013);
nand U6497 (N_6497,N_6130,N_6238);
and U6498 (N_6498,N_6140,N_6193);
nand U6499 (N_6499,N_6158,N_6102);
and U6500 (N_6500,N_6410,N_6406);
nand U6501 (N_6501,N_6377,N_6364);
nor U6502 (N_6502,N_6319,N_6432);
nor U6503 (N_6503,N_6433,N_6408);
or U6504 (N_6504,N_6384,N_6378);
nor U6505 (N_6505,N_6351,N_6389);
nor U6506 (N_6506,N_6369,N_6496);
and U6507 (N_6507,N_6425,N_6276);
and U6508 (N_6508,N_6405,N_6255);
or U6509 (N_6509,N_6388,N_6420);
or U6510 (N_6510,N_6485,N_6392);
and U6511 (N_6511,N_6262,N_6365);
or U6512 (N_6512,N_6346,N_6459);
and U6513 (N_6513,N_6350,N_6301);
nand U6514 (N_6514,N_6292,N_6320);
or U6515 (N_6515,N_6417,N_6329);
xor U6516 (N_6516,N_6285,N_6316);
nor U6517 (N_6517,N_6330,N_6488);
nor U6518 (N_6518,N_6360,N_6254);
or U6519 (N_6519,N_6470,N_6422);
nand U6520 (N_6520,N_6274,N_6297);
and U6521 (N_6521,N_6415,N_6357);
nand U6522 (N_6522,N_6339,N_6426);
nor U6523 (N_6523,N_6493,N_6436);
nand U6524 (N_6524,N_6340,N_6312);
or U6525 (N_6525,N_6321,N_6413);
and U6526 (N_6526,N_6468,N_6454);
or U6527 (N_6527,N_6476,N_6372);
nor U6528 (N_6528,N_6282,N_6299);
and U6529 (N_6529,N_6441,N_6445);
nand U6530 (N_6530,N_6483,N_6469);
nand U6531 (N_6531,N_6491,N_6331);
and U6532 (N_6532,N_6374,N_6379);
nand U6533 (N_6533,N_6337,N_6421);
nand U6534 (N_6534,N_6479,N_6314);
and U6535 (N_6535,N_6451,N_6250);
nand U6536 (N_6536,N_6309,N_6261);
nand U6537 (N_6537,N_6407,N_6411);
nand U6538 (N_6538,N_6387,N_6322);
and U6539 (N_6539,N_6290,N_6391);
and U6540 (N_6540,N_6298,N_6327);
and U6541 (N_6541,N_6423,N_6326);
and U6542 (N_6542,N_6455,N_6318);
nor U6543 (N_6543,N_6341,N_6484);
nand U6544 (N_6544,N_6295,N_6435);
nor U6545 (N_6545,N_6363,N_6283);
and U6546 (N_6546,N_6460,N_6368);
nand U6547 (N_6547,N_6253,N_6296);
nor U6548 (N_6548,N_6278,N_6434);
or U6549 (N_6549,N_6272,N_6307);
nor U6550 (N_6550,N_6464,N_6315);
and U6551 (N_6551,N_6303,N_6490);
and U6552 (N_6552,N_6323,N_6265);
nand U6553 (N_6553,N_6343,N_6430);
and U6554 (N_6554,N_6338,N_6440);
nor U6555 (N_6555,N_6284,N_6251);
or U6556 (N_6556,N_6328,N_6416);
and U6557 (N_6557,N_6317,N_6302);
nand U6558 (N_6558,N_6475,N_6336);
nand U6559 (N_6559,N_6263,N_6489);
or U6560 (N_6560,N_6306,N_6481);
nor U6561 (N_6561,N_6448,N_6449);
xor U6562 (N_6562,N_6443,N_6444);
and U6563 (N_6563,N_6492,N_6452);
or U6564 (N_6564,N_6332,N_6259);
nor U6565 (N_6565,N_6347,N_6264);
nor U6566 (N_6566,N_6359,N_6442);
and U6567 (N_6567,N_6487,N_6308);
nand U6568 (N_6568,N_6271,N_6279);
or U6569 (N_6569,N_6352,N_6333);
nor U6570 (N_6570,N_6472,N_6401);
or U6571 (N_6571,N_6461,N_6256);
nand U6572 (N_6572,N_6258,N_6463);
and U6573 (N_6573,N_6438,N_6412);
or U6574 (N_6574,N_6376,N_6371);
nor U6575 (N_6575,N_6396,N_6345);
and U6576 (N_6576,N_6370,N_6431);
or U6577 (N_6577,N_6462,N_6275);
or U6578 (N_6578,N_6375,N_6394);
nor U6579 (N_6579,N_6467,N_6355);
nand U6580 (N_6580,N_6381,N_6288);
nor U6581 (N_6581,N_6356,N_6429);
nand U6582 (N_6582,N_6287,N_6499);
nor U6583 (N_6583,N_6403,N_6427);
nand U6584 (N_6584,N_6439,N_6478);
and U6585 (N_6585,N_6428,N_6270);
nand U6586 (N_6586,N_6325,N_6313);
and U6587 (N_6587,N_6397,N_6456);
or U6588 (N_6588,N_6294,N_6437);
nand U6589 (N_6589,N_6466,N_6494);
nor U6590 (N_6590,N_6373,N_6398);
or U6591 (N_6591,N_6358,N_6260);
or U6592 (N_6592,N_6273,N_6383);
and U6593 (N_6593,N_6286,N_6471);
nand U6594 (N_6594,N_6362,N_6385);
and U6595 (N_6595,N_6414,N_6404);
nand U6596 (N_6596,N_6366,N_6393);
nand U6597 (N_6597,N_6281,N_6497);
nor U6598 (N_6598,N_6446,N_6293);
nor U6599 (N_6599,N_6486,N_6482);
and U6600 (N_6600,N_6402,N_6419);
or U6601 (N_6601,N_6390,N_6450);
nand U6602 (N_6602,N_6304,N_6342);
xnor U6603 (N_6603,N_6311,N_6458);
or U6604 (N_6604,N_6447,N_6400);
nor U6605 (N_6605,N_6480,N_6335);
or U6606 (N_6606,N_6349,N_6289);
and U6607 (N_6607,N_6495,N_6257);
or U6608 (N_6608,N_6477,N_6399);
or U6609 (N_6609,N_6268,N_6395);
nand U6610 (N_6610,N_6418,N_6291);
or U6611 (N_6611,N_6457,N_6277);
or U6612 (N_6612,N_6324,N_6252);
or U6613 (N_6613,N_6310,N_6465);
or U6614 (N_6614,N_6498,N_6280);
and U6615 (N_6615,N_6367,N_6380);
nand U6616 (N_6616,N_6348,N_6382);
or U6617 (N_6617,N_6453,N_6473);
and U6618 (N_6618,N_6305,N_6269);
nand U6619 (N_6619,N_6344,N_6424);
nor U6620 (N_6620,N_6361,N_6300);
nand U6621 (N_6621,N_6474,N_6266);
nor U6622 (N_6622,N_6409,N_6354);
nor U6623 (N_6623,N_6353,N_6386);
nor U6624 (N_6624,N_6267,N_6334);
nand U6625 (N_6625,N_6446,N_6409);
xnor U6626 (N_6626,N_6364,N_6450);
and U6627 (N_6627,N_6494,N_6469);
or U6628 (N_6628,N_6439,N_6411);
and U6629 (N_6629,N_6486,N_6383);
nand U6630 (N_6630,N_6255,N_6459);
nand U6631 (N_6631,N_6413,N_6299);
nor U6632 (N_6632,N_6287,N_6286);
or U6633 (N_6633,N_6330,N_6381);
nor U6634 (N_6634,N_6441,N_6307);
or U6635 (N_6635,N_6447,N_6441);
or U6636 (N_6636,N_6425,N_6388);
nand U6637 (N_6637,N_6327,N_6328);
and U6638 (N_6638,N_6366,N_6384);
nand U6639 (N_6639,N_6255,N_6335);
nor U6640 (N_6640,N_6383,N_6391);
and U6641 (N_6641,N_6250,N_6483);
nand U6642 (N_6642,N_6285,N_6374);
nand U6643 (N_6643,N_6428,N_6421);
or U6644 (N_6644,N_6294,N_6277);
or U6645 (N_6645,N_6458,N_6264);
and U6646 (N_6646,N_6252,N_6495);
nand U6647 (N_6647,N_6451,N_6338);
or U6648 (N_6648,N_6362,N_6381);
nor U6649 (N_6649,N_6369,N_6488);
and U6650 (N_6650,N_6308,N_6421);
and U6651 (N_6651,N_6290,N_6384);
nor U6652 (N_6652,N_6446,N_6493);
nor U6653 (N_6653,N_6302,N_6361);
nand U6654 (N_6654,N_6487,N_6299);
or U6655 (N_6655,N_6493,N_6454);
and U6656 (N_6656,N_6291,N_6285);
or U6657 (N_6657,N_6498,N_6329);
nand U6658 (N_6658,N_6467,N_6359);
xnor U6659 (N_6659,N_6423,N_6382);
or U6660 (N_6660,N_6385,N_6476);
nor U6661 (N_6661,N_6343,N_6289);
nand U6662 (N_6662,N_6406,N_6474);
nand U6663 (N_6663,N_6461,N_6455);
and U6664 (N_6664,N_6344,N_6397);
or U6665 (N_6665,N_6441,N_6278);
or U6666 (N_6666,N_6356,N_6345);
and U6667 (N_6667,N_6347,N_6383);
xor U6668 (N_6668,N_6274,N_6426);
or U6669 (N_6669,N_6476,N_6480);
nand U6670 (N_6670,N_6319,N_6398);
nand U6671 (N_6671,N_6377,N_6357);
or U6672 (N_6672,N_6485,N_6448);
nand U6673 (N_6673,N_6355,N_6496);
nand U6674 (N_6674,N_6348,N_6262);
or U6675 (N_6675,N_6324,N_6414);
and U6676 (N_6676,N_6382,N_6384);
nor U6677 (N_6677,N_6283,N_6315);
nor U6678 (N_6678,N_6307,N_6359);
and U6679 (N_6679,N_6377,N_6382);
and U6680 (N_6680,N_6447,N_6343);
or U6681 (N_6681,N_6271,N_6349);
nor U6682 (N_6682,N_6430,N_6465);
nand U6683 (N_6683,N_6269,N_6258);
nand U6684 (N_6684,N_6472,N_6431);
nor U6685 (N_6685,N_6391,N_6285);
and U6686 (N_6686,N_6362,N_6301);
and U6687 (N_6687,N_6370,N_6302);
or U6688 (N_6688,N_6320,N_6283);
or U6689 (N_6689,N_6254,N_6383);
and U6690 (N_6690,N_6399,N_6423);
and U6691 (N_6691,N_6389,N_6296);
and U6692 (N_6692,N_6443,N_6309);
or U6693 (N_6693,N_6415,N_6451);
or U6694 (N_6694,N_6256,N_6285);
nor U6695 (N_6695,N_6458,N_6472);
and U6696 (N_6696,N_6323,N_6435);
and U6697 (N_6697,N_6253,N_6298);
nand U6698 (N_6698,N_6310,N_6393);
or U6699 (N_6699,N_6498,N_6296);
and U6700 (N_6700,N_6385,N_6443);
or U6701 (N_6701,N_6447,N_6456);
and U6702 (N_6702,N_6325,N_6254);
nor U6703 (N_6703,N_6385,N_6273);
and U6704 (N_6704,N_6346,N_6362);
and U6705 (N_6705,N_6312,N_6390);
or U6706 (N_6706,N_6253,N_6499);
and U6707 (N_6707,N_6337,N_6435);
and U6708 (N_6708,N_6300,N_6492);
nor U6709 (N_6709,N_6362,N_6387);
nand U6710 (N_6710,N_6456,N_6469);
or U6711 (N_6711,N_6338,N_6320);
and U6712 (N_6712,N_6379,N_6443);
and U6713 (N_6713,N_6370,N_6374);
xor U6714 (N_6714,N_6275,N_6315);
nor U6715 (N_6715,N_6332,N_6319);
nand U6716 (N_6716,N_6411,N_6349);
nor U6717 (N_6717,N_6381,N_6305);
nand U6718 (N_6718,N_6390,N_6306);
nand U6719 (N_6719,N_6350,N_6254);
or U6720 (N_6720,N_6338,N_6483);
or U6721 (N_6721,N_6332,N_6385);
nand U6722 (N_6722,N_6339,N_6251);
nand U6723 (N_6723,N_6330,N_6428);
nand U6724 (N_6724,N_6457,N_6297);
nor U6725 (N_6725,N_6329,N_6411);
nor U6726 (N_6726,N_6367,N_6304);
or U6727 (N_6727,N_6423,N_6259);
and U6728 (N_6728,N_6490,N_6327);
nor U6729 (N_6729,N_6464,N_6401);
and U6730 (N_6730,N_6346,N_6492);
nand U6731 (N_6731,N_6356,N_6441);
xor U6732 (N_6732,N_6292,N_6427);
or U6733 (N_6733,N_6409,N_6283);
nor U6734 (N_6734,N_6380,N_6280);
or U6735 (N_6735,N_6426,N_6446);
nand U6736 (N_6736,N_6326,N_6486);
or U6737 (N_6737,N_6464,N_6285);
and U6738 (N_6738,N_6493,N_6357);
nand U6739 (N_6739,N_6440,N_6258);
or U6740 (N_6740,N_6280,N_6275);
nand U6741 (N_6741,N_6324,N_6481);
xnor U6742 (N_6742,N_6376,N_6453);
or U6743 (N_6743,N_6395,N_6458);
nand U6744 (N_6744,N_6283,N_6375);
and U6745 (N_6745,N_6378,N_6437);
or U6746 (N_6746,N_6462,N_6368);
nor U6747 (N_6747,N_6393,N_6262);
nor U6748 (N_6748,N_6292,N_6356);
xor U6749 (N_6749,N_6374,N_6289);
and U6750 (N_6750,N_6589,N_6718);
nor U6751 (N_6751,N_6743,N_6620);
nor U6752 (N_6752,N_6606,N_6553);
xor U6753 (N_6753,N_6622,N_6657);
nor U6754 (N_6754,N_6633,N_6719);
nand U6755 (N_6755,N_6660,N_6698);
nand U6756 (N_6756,N_6680,N_6616);
nor U6757 (N_6757,N_6598,N_6571);
or U6758 (N_6758,N_6639,N_6576);
and U6759 (N_6759,N_6610,N_6720);
xnor U6760 (N_6760,N_6645,N_6686);
or U6761 (N_6761,N_6659,N_6525);
and U6762 (N_6762,N_6600,N_6629);
or U6763 (N_6763,N_6684,N_6510);
or U6764 (N_6764,N_6537,N_6575);
nor U6765 (N_6765,N_6584,N_6527);
nor U6766 (N_6766,N_6617,N_6564);
nor U6767 (N_6767,N_6634,N_6685);
or U6768 (N_6768,N_6710,N_6565);
nand U6769 (N_6769,N_6627,N_6592);
and U6770 (N_6770,N_6672,N_6649);
or U6771 (N_6771,N_6585,N_6513);
nor U6772 (N_6772,N_6574,N_6563);
nand U6773 (N_6773,N_6745,N_6579);
and U6774 (N_6774,N_6604,N_6688);
nor U6775 (N_6775,N_6643,N_6562);
nand U6776 (N_6776,N_6665,N_6702);
or U6777 (N_6777,N_6524,N_6742);
nor U6778 (N_6778,N_6637,N_6542);
and U6779 (N_6779,N_6550,N_6729);
or U6780 (N_6780,N_6614,N_6601);
or U6781 (N_6781,N_6667,N_6648);
or U6782 (N_6782,N_6568,N_6518);
xor U6783 (N_6783,N_6597,N_6652);
nor U6784 (N_6784,N_6683,N_6746);
or U6785 (N_6785,N_6551,N_6586);
nor U6786 (N_6786,N_6572,N_6739);
and U6787 (N_6787,N_6544,N_6695);
or U6788 (N_6788,N_6632,N_6594);
nand U6789 (N_6789,N_6694,N_6658);
nand U6790 (N_6790,N_6602,N_6500);
nor U6791 (N_6791,N_6512,N_6609);
or U6792 (N_6792,N_6715,N_6504);
nor U6793 (N_6793,N_6635,N_6619);
or U6794 (N_6794,N_6740,N_6555);
nor U6795 (N_6795,N_6613,N_6734);
nor U6796 (N_6796,N_6728,N_6726);
nor U6797 (N_6797,N_6663,N_6717);
nor U6798 (N_6798,N_6681,N_6590);
or U6799 (N_6799,N_6674,N_6661);
nor U6800 (N_6800,N_6559,N_6650);
and U6801 (N_6801,N_6538,N_6607);
or U6802 (N_6802,N_6647,N_6541);
or U6803 (N_6803,N_6546,N_6682);
xor U6804 (N_6804,N_6503,N_6515);
nor U6805 (N_6805,N_6519,N_6588);
nor U6806 (N_6806,N_6548,N_6630);
or U6807 (N_6807,N_6547,N_6511);
nor U6808 (N_6808,N_6703,N_6711);
and U6809 (N_6809,N_6516,N_6611);
nor U6810 (N_6810,N_6706,N_6696);
nor U6811 (N_6811,N_6505,N_6520);
and U6812 (N_6812,N_6501,N_6733);
nand U6813 (N_6813,N_6699,N_6693);
nand U6814 (N_6814,N_6705,N_6725);
and U6815 (N_6815,N_6689,N_6608);
or U6816 (N_6816,N_6673,N_6552);
and U6817 (N_6817,N_6536,N_6612);
nand U6818 (N_6818,N_6531,N_6721);
or U6819 (N_6819,N_6664,N_6567);
and U6820 (N_6820,N_6596,N_6549);
nand U6821 (N_6821,N_6566,N_6646);
and U6822 (N_6822,N_6662,N_6626);
nor U6823 (N_6823,N_6535,N_6605);
nor U6824 (N_6824,N_6692,N_6624);
and U6825 (N_6825,N_6533,N_6603);
or U6826 (N_6826,N_6507,N_6561);
and U6827 (N_6827,N_6671,N_6628);
and U6828 (N_6828,N_6625,N_6655);
or U6829 (N_6829,N_6560,N_6528);
nand U6830 (N_6830,N_6723,N_6523);
and U6831 (N_6831,N_6631,N_6716);
or U6832 (N_6832,N_6508,N_6690);
nor U6833 (N_6833,N_6534,N_6582);
and U6834 (N_6834,N_6540,N_6581);
nand U6835 (N_6835,N_6687,N_6545);
nand U6836 (N_6836,N_6678,N_6744);
or U6837 (N_6837,N_6618,N_6591);
xnor U6838 (N_6838,N_6653,N_6595);
and U6839 (N_6839,N_6509,N_6735);
and U6840 (N_6840,N_6641,N_6707);
nor U6841 (N_6841,N_6676,N_6670);
nor U6842 (N_6842,N_6656,N_6517);
or U6843 (N_6843,N_6691,N_6677);
or U6844 (N_6844,N_6701,N_6526);
nor U6845 (N_6845,N_6741,N_6668);
nand U6846 (N_6846,N_6714,N_6640);
or U6847 (N_6847,N_6724,N_6654);
nor U6848 (N_6848,N_6569,N_6578);
nor U6849 (N_6849,N_6679,N_6736);
and U6850 (N_6850,N_6530,N_6539);
nor U6851 (N_6851,N_6713,N_6712);
and U6852 (N_6852,N_6583,N_6573);
or U6853 (N_6853,N_6666,N_6732);
and U6854 (N_6854,N_6543,N_6556);
nor U6855 (N_6855,N_6737,N_6554);
and U6856 (N_6856,N_6532,N_6558);
or U6857 (N_6857,N_6502,N_6506);
nand U6858 (N_6858,N_6521,N_6621);
nand U6859 (N_6859,N_6577,N_6731);
or U6860 (N_6860,N_6738,N_6636);
nor U6861 (N_6861,N_6638,N_6747);
nand U6862 (N_6862,N_6749,N_6587);
and U6863 (N_6863,N_6709,N_6748);
nor U6864 (N_6864,N_6580,N_6599);
or U6865 (N_6865,N_6651,N_6522);
nand U6866 (N_6866,N_6730,N_6570);
and U6867 (N_6867,N_6697,N_6615);
and U6868 (N_6868,N_6529,N_6708);
or U6869 (N_6869,N_6557,N_6593);
nand U6870 (N_6870,N_6722,N_6675);
nor U6871 (N_6871,N_6644,N_6623);
nand U6872 (N_6872,N_6704,N_6727);
or U6873 (N_6873,N_6669,N_6514);
or U6874 (N_6874,N_6642,N_6700);
nand U6875 (N_6875,N_6739,N_6710);
and U6876 (N_6876,N_6662,N_6695);
nand U6877 (N_6877,N_6643,N_6535);
nor U6878 (N_6878,N_6520,N_6608);
nand U6879 (N_6879,N_6696,N_6560);
nor U6880 (N_6880,N_6563,N_6508);
nand U6881 (N_6881,N_6613,N_6709);
and U6882 (N_6882,N_6636,N_6727);
nor U6883 (N_6883,N_6607,N_6726);
nor U6884 (N_6884,N_6639,N_6556);
nor U6885 (N_6885,N_6578,N_6550);
and U6886 (N_6886,N_6676,N_6698);
nand U6887 (N_6887,N_6643,N_6675);
nor U6888 (N_6888,N_6722,N_6546);
nand U6889 (N_6889,N_6551,N_6573);
nand U6890 (N_6890,N_6543,N_6659);
or U6891 (N_6891,N_6590,N_6677);
or U6892 (N_6892,N_6636,N_6730);
and U6893 (N_6893,N_6558,N_6662);
and U6894 (N_6894,N_6603,N_6613);
or U6895 (N_6895,N_6570,N_6501);
nand U6896 (N_6896,N_6678,N_6710);
nand U6897 (N_6897,N_6729,N_6674);
or U6898 (N_6898,N_6732,N_6690);
and U6899 (N_6899,N_6700,N_6567);
and U6900 (N_6900,N_6510,N_6656);
nand U6901 (N_6901,N_6543,N_6612);
nand U6902 (N_6902,N_6526,N_6582);
nor U6903 (N_6903,N_6540,N_6548);
or U6904 (N_6904,N_6581,N_6544);
nor U6905 (N_6905,N_6518,N_6722);
and U6906 (N_6906,N_6598,N_6674);
or U6907 (N_6907,N_6627,N_6640);
nor U6908 (N_6908,N_6633,N_6592);
nand U6909 (N_6909,N_6508,N_6687);
or U6910 (N_6910,N_6665,N_6566);
and U6911 (N_6911,N_6522,N_6598);
nor U6912 (N_6912,N_6739,N_6707);
nor U6913 (N_6913,N_6630,N_6636);
or U6914 (N_6914,N_6739,N_6708);
nand U6915 (N_6915,N_6591,N_6542);
xnor U6916 (N_6916,N_6626,N_6701);
nor U6917 (N_6917,N_6597,N_6683);
or U6918 (N_6918,N_6649,N_6602);
nor U6919 (N_6919,N_6690,N_6615);
or U6920 (N_6920,N_6702,N_6729);
and U6921 (N_6921,N_6671,N_6682);
nor U6922 (N_6922,N_6714,N_6614);
or U6923 (N_6923,N_6644,N_6741);
nand U6924 (N_6924,N_6594,N_6536);
nand U6925 (N_6925,N_6658,N_6620);
or U6926 (N_6926,N_6634,N_6674);
nor U6927 (N_6927,N_6628,N_6537);
nor U6928 (N_6928,N_6595,N_6542);
and U6929 (N_6929,N_6669,N_6529);
nand U6930 (N_6930,N_6701,N_6659);
and U6931 (N_6931,N_6743,N_6740);
nand U6932 (N_6932,N_6506,N_6584);
or U6933 (N_6933,N_6606,N_6576);
nand U6934 (N_6934,N_6532,N_6676);
xor U6935 (N_6935,N_6538,N_6537);
and U6936 (N_6936,N_6570,N_6557);
nor U6937 (N_6937,N_6515,N_6645);
nor U6938 (N_6938,N_6503,N_6513);
or U6939 (N_6939,N_6547,N_6586);
nand U6940 (N_6940,N_6627,N_6572);
and U6941 (N_6941,N_6534,N_6539);
nand U6942 (N_6942,N_6719,N_6652);
nand U6943 (N_6943,N_6649,N_6659);
nand U6944 (N_6944,N_6544,N_6749);
or U6945 (N_6945,N_6644,N_6607);
nand U6946 (N_6946,N_6611,N_6638);
nor U6947 (N_6947,N_6701,N_6538);
nor U6948 (N_6948,N_6577,N_6560);
or U6949 (N_6949,N_6661,N_6514);
nor U6950 (N_6950,N_6624,N_6665);
nand U6951 (N_6951,N_6696,N_6702);
nand U6952 (N_6952,N_6623,N_6548);
nor U6953 (N_6953,N_6608,N_6571);
and U6954 (N_6954,N_6660,N_6686);
and U6955 (N_6955,N_6692,N_6672);
xnor U6956 (N_6956,N_6668,N_6574);
xor U6957 (N_6957,N_6595,N_6643);
nand U6958 (N_6958,N_6713,N_6515);
nor U6959 (N_6959,N_6685,N_6638);
nand U6960 (N_6960,N_6547,N_6724);
nor U6961 (N_6961,N_6556,N_6643);
nor U6962 (N_6962,N_6729,N_6570);
nand U6963 (N_6963,N_6681,N_6624);
and U6964 (N_6964,N_6546,N_6550);
nand U6965 (N_6965,N_6729,N_6633);
nor U6966 (N_6966,N_6637,N_6521);
or U6967 (N_6967,N_6626,N_6549);
and U6968 (N_6968,N_6537,N_6541);
nand U6969 (N_6969,N_6517,N_6687);
or U6970 (N_6970,N_6519,N_6746);
and U6971 (N_6971,N_6655,N_6567);
or U6972 (N_6972,N_6513,N_6630);
or U6973 (N_6973,N_6697,N_6636);
and U6974 (N_6974,N_6636,N_6510);
nor U6975 (N_6975,N_6650,N_6628);
or U6976 (N_6976,N_6525,N_6506);
nor U6977 (N_6977,N_6746,N_6626);
nor U6978 (N_6978,N_6613,N_6521);
nand U6979 (N_6979,N_6528,N_6706);
xor U6980 (N_6980,N_6574,N_6731);
or U6981 (N_6981,N_6536,N_6554);
nor U6982 (N_6982,N_6548,N_6743);
xor U6983 (N_6983,N_6708,N_6530);
nand U6984 (N_6984,N_6686,N_6571);
and U6985 (N_6985,N_6731,N_6533);
nor U6986 (N_6986,N_6637,N_6689);
or U6987 (N_6987,N_6557,N_6715);
nor U6988 (N_6988,N_6518,N_6684);
or U6989 (N_6989,N_6665,N_6727);
nand U6990 (N_6990,N_6526,N_6702);
nor U6991 (N_6991,N_6646,N_6657);
nor U6992 (N_6992,N_6620,N_6714);
or U6993 (N_6993,N_6740,N_6698);
nor U6994 (N_6994,N_6599,N_6586);
nor U6995 (N_6995,N_6600,N_6689);
nor U6996 (N_6996,N_6589,N_6623);
or U6997 (N_6997,N_6713,N_6695);
or U6998 (N_6998,N_6542,N_6648);
nand U6999 (N_6999,N_6546,N_6718);
or U7000 (N_7000,N_6870,N_6940);
nor U7001 (N_7001,N_6766,N_6802);
and U7002 (N_7002,N_6964,N_6996);
nand U7003 (N_7003,N_6763,N_6975);
and U7004 (N_7004,N_6862,N_6791);
nand U7005 (N_7005,N_6769,N_6851);
nand U7006 (N_7006,N_6965,N_6859);
and U7007 (N_7007,N_6815,N_6987);
nor U7008 (N_7008,N_6918,N_6788);
or U7009 (N_7009,N_6784,N_6972);
and U7010 (N_7010,N_6892,N_6895);
nand U7011 (N_7011,N_6782,N_6982);
nand U7012 (N_7012,N_6807,N_6830);
and U7013 (N_7013,N_6871,N_6900);
nand U7014 (N_7014,N_6818,N_6772);
nand U7015 (N_7015,N_6989,N_6935);
nand U7016 (N_7016,N_6875,N_6909);
nor U7017 (N_7017,N_6865,N_6777);
or U7018 (N_7018,N_6798,N_6752);
nand U7019 (N_7019,N_6923,N_6957);
xor U7020 (N_7020,N_6755,N_6829);
nand U7021 (N_7021,N_6959,N_6955);
nand U7022 (N_7022,N_6898,N_6878);
and U7023 (N_7023,N_6894,N_6917);
or U7024 (N_7024,N_6781,N_6757);
and U7025 (N_7025,N_6933,N_6966);
nor U7026 (N_7026,N_6961,N_6984);
or U7027 (N_7027,N_6879,N_6799);
nand U7028 (N_7028,N_6953,N_6845);
nor U7029 (N_7029,N_6942,N_6974);
and U7030 (N_7030,N_6805,N_6794);
nand U7031 (N_7031,N_6843,N_6817);
or U7032 (N_7032,N_6868,N_6911);
nand U7033 (N_7033,N_6978,N_6992);
nand U7034 (N_7034,N_6759,N_6967);
nand U7035 (N_7035,N_6867,N_6880);
nor U7036 (N_7036,N_6834,N_6920);
nand U7037 (N_7037,N_6869,N_6764);
or U7038 (N_7038,N_6842,N_6884);
nand U7039 (N_7039,N_6927,N_6952);
or U7040 (N_7040,N_6886,N_6991);
nand U7041 (N_7041,N_6821,N_6872);
and U7042 (N_7042,N_6806,N_6928);
or U7043 (N_7043,N_6994,N_6810);
nor U7044 (N_7044,N_6753,N_6812);
or U7045 (N_7045,N_6931,N_6841);
nor U7046 (N_7046,N_6941,N_6877);
or U7047 (N_7047,N_6932,N_6874);
nand U7048 (N_7048,N_6924,N_6919);
nor U7049 (N_7049,N_6760,N_6770);
and U7050 (N_7050,N_6863,N_6793);
or U7051 (N_7051,N_6993,N_6887);
nand U7052 (N_7052,N_6826,N_6925);
and U7053 (N_7053,N_6885,N_6979);
nand U7054 (N_7054,N_6990,N_6896);
and U7055 (N_7055,N_6881,N_6997);
and U7056 (N_7056,N_6891,N_6903);
nor U7057 (N_7057,N_6803,N_6801);
nand U7058 (N_7058,N_6944,N_6751);
or U7059 (N_7059,N_6850,N_6762);
nor U7060 (N_7060,N_6939,N_6837);
nor U7061 (N_7061,N_6767,N_6902);
nor U7062 (N_7062,N_6789,N_6840);
or U7063 (N_7063,N_6914,N_6866);
nor U7064 (N_7064,N_6983,N_6838);
and U7065 (N_7065,N_6824,N_6936);
nor U7066 (N_7066,N_6882,N_6930);
nor U7067 (N_7067,N_6937,N_6949);
and U7068 (N_7068,N_6980,N_6943);
and U7069 (N_7069,N_6778,N_6853);
nand U7070 (N_7070,N_6827,N_6904);
and U7071 (N_7071,N_6861,N_6999);
nor U7072 (N_7072,N_6883,N_6795);
and U7073 (N_7073,N_6948,N_6796);
or U7074 (N_7074,N_6906,N_6846);
or U7075 (N_7075,N_6934,N_6968);
nand U7076 (N_7076,N_6986,N_6776);
and U7077 (N_7077,N_6787,N_6773);
nor U7078 (N_7078,N_6962,N_6988);
or U7079 (N_7079,N_6831,N_6901);
or U7080 (N_7080,N_6908,N_6783);
or U7081 (N_7081,N_6971,N_6907);
or U7082 (N_7082,N_6864,N_6780);
and U7083 (N_7083,N_6956,N_6844);
or U7084 (N_7084,N_6893,N_6808);
nor U7085 (N_7085,N_6820,N_6899);
nor U7086 (N_7086,N_6958,N_6779);
nand U7087 (N_7087,N_6897,N_6819);
and U7088 (N_7088,N_6774,N_6910);
nor U7089 (N_7089,N_6889,N_6848);
nand U7090 (N_7090,N_6938,N_6954);
and U7091 (N_7091,N_6945,N_6970);
nor U7092 (N_7092,N_6790,N_6761);
and U7093 (N_7093,N_6951,N_6922);
nor U7094 (N_7094,N_6832,N_6855);
and U7095 (N_7095,N_6768,N_6756);
nand U7096 (N_7096,N_6976,N_6985);
or U7097 (N_7097,N_6828,N_6792);
or U7098 (N_7098,N_6811,N_6809);
or U7099 (N_7099,N_6804,N_6981);
nor U7100 (N_7100,N_6916,N_6977);
and U7101 (N_7101,N_6950,N_6814);
nand U7102 (N_7102,N_6960,N_6946);
or U7103 (N_7103,N_6926,N_6888);
nor U7104 (N_7104,N_6849,N_6890);
nand U7105 (N_7105,N_6785,N_6856);
nand U7106 (N_7106,N_6825,N_6775);
and U7107 (N_7107,N_6912,N_6847);
nor U7108 (N_7108,N_6873,N_6823);
or U7109 (N_7109,N_6813,N_6822);
nand U7110 (N_7110,N_6771,N_6913);
nor U7111 (N_7111,N_6929,N_6876);
nor U7112 (N_7112,N_6852,N_6750);
nand U7113 (N_7113,N_6835,N_6998);
and U7114 (N_7114,N_6854,N_6969);
nor U7115 (N_7115,N_6963,N_6947);
and U7116 (N_7116,N_6839,N_6860);
or U7117 (N_7117,N_6921,N_6857);
or U7118 (N_7118,N_6858,N_6915);
nand U7119 (N_7119,N_6833,N_6797);
and U7120 (N_7120,N_6758,N_6995);
and U7121 (N_7121,N_6765,N_6816);
xnor U7122 (N_7122,N_6905,N_6754);
nand U7123 (N_7123,N_6836,N_6800);
or U7124 (N_7124,N_6973,N_6786);
nor U7125 (N_7125,N_6914,N_6860);
nand U7126 (N_7126,N_6972,N_6910);
nand U7127 (N_7127,N_6753,N_6798);
and U7128 (N_7128,N_6914,N_6840);
nand U7129 (N_7129,N_6922,N_6783);
or U7130 (N_7130,N_6977,N_6837);
and U7131 (N_7131,N_6807,N_6841);
nand U7132 (N_7132,N_6809,N_6871);
nor U7133 (N_7133,N_6942,N_6987);
nand U7134 (N_7134,N_6956,N_6778);
or U7135 (N_7135,N_6924,N_6827);
and U7136 (N_7136,N_6977,N_6955);
or U7137 (N_7137,N_6884,N_6776);
or U7138 (N_7138,N_6770,N_6836);
and U7139 (N_7139,N_6777,N_6981);
nor U7140 (N_7140,N_6801,N_6841);
or U7141 (N_7141,N_6986,N_6859);
nor U7142 (N_7142,N_6804,N_6953);
and U7143 (N_7143,N_6976,N_6885);
or U7144 (N_7144,N_6906,N_6945);
or U7145 (N_7145,N_6802,N_6976);
nor U7146 (N_7146,N_6875,N_6801);
or U7147 (N_7147,N_6883,N_6881);
and U7148 (N_7148,N_6848,N_6894);
and U7149 (N_7149,N_6761,N_6924);
and U7150 (N_7150,N_6992,N_6844);
and U7151 (N_7151,N_6972,N_6926);
nor U7152 (N_7152,N_6947,N_6768);
nor U7153 (N_7153,N_6790,N_6897);
and U7154 (N_7154,N_6951,N_6994);
and U7155 (N_7155,N_6979,N_6884);
and U7156 (N_7156,N_6760,N_6992);
nor U7157 (N_7157,N_6882,N_6941);
or U7158 (N_7158,N_6900,N_6920);
xnor U7159 (N_7159,N_6890,N_6764);
nor U7160 (N_7160,N_6829,N_6831);
or U7161 (N_7161,N_6993,N_6862);
and U7162 (N_7162,N_6753,N_6790);
nor U7163 (N_7163,N_6912,N_6999);
or U7164 (N_7164,N_6989,N_6820);
nor U7165 (N_7165,N_6822,N_6828);
xor U7166 (N_7166,N_6895,N_6920);
or U7167 (N_7167,N_6903,N_6897);
nand U7168 (N_7168,N_6903,N_6851);
nand U7169 (N_7169,N_6785,N_6916);
or U7170 (N_7170,N_6845,N_6929);
or U7171 (N_7171,N_6766,N_6818);
and U7172 (N_7172,N_6816,N_6961);
and U7173 (N_7173,N_6849,N_6974);
nor U7174 (N_7174,N_6801,N_6775);
and U7175 (N_7175,N_6758,N_6767);
or U7176 (N_7176,N_6999,N_6771);
nand U7177 (N_7177,N_6795,N_6859);
or U7178 (N_7178,N_6914,N_6867);
nand U7179 (N_7179,N_6814,N_6797);
and U7180 (N_7180,N_6913,N_6842);
or U7181 (N_7181,N_6997,N_6849);
and U7182 (N_7182,N_6871,N_6778);
and U7183 (N_7183,N_6798,N_6986);
xnor U7184 (N_7184,N_6857,N_6757);
nor U7185 (N_7185,N_6837,N_6875);
nand U7186 (N_7186,N_6977,N_6779);
and U7187 (N_7187,N_6813,N_6982);
nor U7188 (N_7188,N_6986,N_6909);
nor U7189 (N_7189,N_6835,N_6973);
nor U7190 (N_7190,N_6909,N_6806);
or U7191 (N_7191,N_6842,N_6885);
nor U7192 (N_7192,N_6897,N_6937);
xnor U7193 (N_7193,N_6972,N_6799);
and U7194 (N_7194,N_6832,N_6764);
or U7195 (N_7195,N_6806,N_6950);
xnor U7196 (N_7196,N_6876,N_6852);
or U7197 (N_7197,N_6995,N_6877);
and U7198 (N_7198,N_6963,N_6986);
and U7199 (N_7199,N_6902,N_6935);
and U7200 (N_7200,N_6839,N_6974);
or U7201 (N_7201,N_6954,N_6905);
nand U7202 (N_7202,N_6902,N_6776);
or U7203 (N_7203,N_6879,N_6792);
or U7204 (N_7204,N_6960,N_6883);
or U7205 (N_7205,N_6962,N_6858);
and U7206 (N_7206,N_6954,N_6922);
nand U7207 (N_7207,N_6813,N_6884);
xnor U7208 (N_7208,N_6918,N_6962);
nor U7209 (N_7209,N_6931,N_6925);
nand U7210 (N_7210,N_6898,N_6927);
nor U7211 (N_7211,N_6950,N_6927);
or U7212 (N_7212,N_6916,N_6959);
nand U7213 (N_7213,N_6915,N_6889);
and U7214 (N_7214,N_6961,N_6848);
or U7215 (N_7215,N_6854,N_6857);
and U7216 (N_7216,N_6797,N_6869);
nor U7217 (N_7217,N_6917,N_6866);
nor U7218 (N_7218,N_6936,N_6922);
or U7219 (N_7219,N_6932,N_6768);
and U7220 (N_7220,N_6840,N_6750);
or U7221 (N_7221,N_6983,N_6866);
nor U7222 (N_7222,N_6756,N_6909);
nor U7223 (N_7223,N_6893,N_6928);
nor U7224 (N_7224,N_6891,N_6934);
or U7225 (N_7225,N_6888,N_6850);
nand U7226 (N_7226,N_6842,N_6875);
or U7227 (N_7227,N_6995,N_6950);
nand U7228 (N_7228,N_6756,N_6806);
nand U7229 (N_7229,N_6787,N_6842);
or U7230 (N_7230,N_6950,N_6812);
and U7231 (N_7231,N_6762,N_6869);
xnor U7232 (N_7232,N_6785,N_6931);
and U7233 (N_7233,N_6953,N_6806);
and U7234 (N_7234,N_6939,N_6904);
and U7235 (N_7235,N_6951,N_6875);
nor U7236 (N_7236,N_6759,N_6939);
nand U7237 (N_7237,N_6955,N_6796);
nor U7238 (N_7238,N_6879,N_6813);
nand U7239 (N_7239,N_6855,N_6856);
nand U7240 (N_7240,N_6967,N_6762);
or U7241 (N_7241,N_6852,N_6895);
or U7242 (N_7242,N_6936,N_6875);
nand U7243 (N_7243,N_6883,N_6963);
or U7244 (N_7244,N_6997,N_6978);
or U7245 (N_7245,N_6855,N_6996);
or U7246 (N_7246,N_6992,N_6817);
nand U7247 (N_7247,N_6844,N_6919);
nor U7248 (N_7248,N_6887,N_6966);
or U7249 (N_7249,N_6887,N_6900);
or U7250 (N_7250,N_7180,N_7198);
and U7251 (N_7251,N_7227,N_7195);
or U7252 (N_7252,N_7147,N_7154);
or U7253 (N_7253,N_7030,N_7202);
nand U7254 (N_7254,N_7112,N_7185);
nand U7255 (N_7255,N_7183,N_7146);
nor U7256 (N_7256,N_7001,N_7222);
nand U7257 (N_7257,N_7208,N_7033);
and U7258 (N_7258,N_7246,N_7170);
nor U7259 (N_7259,N_7068,N_7017);
nor U7260 (N_7260,N_7213,N_7187);
or U7261 (N_7261,N_7144,N_7150);
and U7262 (N_7262,N_7124,N_7020);
nor U7263 (N_7263,N_7091,N_7133);
nand U7264 (N_7264,N_7045,N_7101);
nand U7265 (N_7265,N_7070,N_7142);
or U7266 (N_7266,N_7216,N_7244);
nor U7267 (N_7267,N_7240,N_7184);
and U7268 (N_7268,N_7005,N_7140);
nand U7269 (N_7269,N_7156,N_7158);
nor U7270 (N_7270,N_7046,N_7115);
or U7271 (N_7271,N_7127,N_7120);
nand U7272 (N_7272,N_7074,N_7160);
nor U7273 (N_7273,N_7152,N_7040);
or U7274 (N_7274,N_7036,N_7097);
and U7275 (N_7275,N_7118,N_7065);
nand U7276 (N_7276,N_7137,N_7110);
nand U7277 (N_7277,N_7194,N_7229);
or U7278 (N_7278,N_7052,N_7159);
and U7279 (N_7279,N_7196,N_7089);
nand U7280 (N_7280,N_7051,N_7149);
xor U7281 (N_7281,N_7123,N_7131);
nor U7282 (N_7282,N_7027,N_7225);
nor U7283 (N_7283,N_7230,N_7226);
nor U7284 (N_7284,N_7143,N_7069);
and U7285 (N_7285,N_7199,N_7206);
nor U7286 (N_7286,N_7163,N_7009);
and U7287 (N_7287,N_7145,N_7129);
or U7288 (N_7288,N_7031,N_7054);
or U7289 (N_7289,N_7197,N_7073);
nor U7290 (N_7290,N_7011,N_7077);
or U7291 (N_7291,N_7221,N_7168);
nand U7292 (N_7292,N_7016,N_7004);
nor U7293 (N_7293,N_7214,N_7105);
or U7294 (N_7294,N_7039,N_7037);
or U7295 (N_7295,N_7201,N_7026);
and U7296 (N_7296,N_7042,N_7003);
nor U7297 (N_7297,N_7023,N_7243);
nor U7298 (N_7298,N_7058,N_7122);
nor U7299 (N_7299,N_7109,N_7116);
or U7300 (N_7300,N_7192,N_7095);
nand U7301 (N_7301,N_7041,N_7162);
nor U7302 (N_7302,N_7151,N_7044);
and U7303 (N_7303,N_7075,N_7107);
nand U7304 (N_7304,N_7203,N_7241);
and U7305 (N_7305,N_7157,N_7093);
nand U7306 (N_7306,N_7130,N_7234);
nand U7307 (N_7307,N_7181,N_7148);
and U7308 (N_7308,N_7237,N_7153);
and U7309 (N_7309,N_7238,N_7248);
nand U7310 (N_7310,N_7071,N_7247);
nand U7311 (N_7311,N_7078,N_7114);
nor U7312 (N_7312,N_7135,N_7191);
nand U7313 (N_7313,N_7066,N_7060);
or U7314 (N_7314,N_7007,N_7028);
and U7315 (N_7315,N_7220,N_7128);
nand U7316 (N_7316,N_7174,N_7102);
or U7317 (N_7317,N_7175,N_7249);
or U7318 (N_7318,N_7098,N_7165);
nor U7319 (N_7319,N_7164,N_7090);
nor U7320 (N_7320,N_7121,N_7218);
or U7321 (N_7321,N_7108,N_7186);
nand U7322 (N_7322,N_7032,N_7106);
nor U7323 (N_7323,N_7207,N_7067);
nor U7324 (N_7324,N_7022,N_7053);
nand U7325 (N_7325,N_7057,N_7119);
nand U7326 (N_7326,N_7200,N_7092);
nand U7327 (N_7327,N_7002,N_7166);
nand U7328 (N_7328,N_7013,N_7193);
nand U7329 (N_7329,N_7204,N_7233);
and U7330 (N_7330,N_7217,N_7178);
nor U7331 (N_7331,N_7048,N_7035);
or U7332 (N_7332,N_7094,N_7043);
nor U7333 (N_7333,N_7117,N_7008);
or U7334 (N_7334,N_7096,N_7161);
nor U7335 (N_7335,N_7072,N_7099);
or U7336 (N_7336,N_7000,N_7083);
and U7337 (N_7337,N_7215,N_7239);
nand U7338 (N_7338,N_7080,N_7061);
or U7339 (N_7339,N_7006,N_7113);
or U7340 (N_7340,N_7103,N_7029);
nand U7341 (N_7341,N_7019,N_7138);
nor U7342 (N_7342,N_7111,N_7212);
and U7343 (N_7343,N_7219,N_7169);
and U7344 (N_7344,N_7167,N_7055);
nor U7345 (N_7345,N_7173,N_7176);
nor U7346 (N_7346,N_7232,N_7228);
nand U7347 (N_7347,N_7014,N_7236);
nor U7348 (N_7348,N_7079,N_7125);
and U7349 (N_7349,N_7209,N_7085);
nand U7350 (N_7350,N_7171,N_7038);
nor U7351 (N_7351,N_7021,N_7104);
or U7352 (N_7352,N_7081,N_7224);
and U7353 (N_7353,N_7063,N_7132);
nor U7354 (N_7354,N_7179,N_7015);
xnor U7355 (N_7355,N_7231,N_7205);
and U7356 (N_7356,N_7088,N_7018);
nor U7357 (N_7357,N_7050,N_7012);
or U7358 (N_7358,N_7062,N_7155);
or U7359 (N_7359,N_7126,N_7024);
nor U7360 (N_7360,N_7136,N_7082);
nor U7361 (N_7361,N_7100,N_7134);
nor U7362 (N_7362,N_7010,N_7242);
or U7363 (N_7363,N_7182,N_7025);
or U7364 (N_7364,N_7086,N_7034);
nor U7365 (N_7365,N_7049,N_7087);
nand U7366 (N_7366,N_7235,N_7211);
nor U7367 (N_7367,N_7190,N_7223);
xnor U7368 (N_7368,N_7189,N_7084);
nand U7369 (N_7369,N_7177,N_7059);
nor U7370 (N_7370,N_7245,N_7076);
or U7371 (N_7371,N_7056,N_7172);
and U7372 (N_7372,N_7210,N_7139);
or U7373 (N_7373,N_7188,N_7064);
or U7374 (N_7374,N_7047,N_7141);
nand U7375 (N_7375,N_7059,N_7078);
nand U7376 (N_7376,N_7056,N_7217);
nor U7377 (N_7377,N_7027,N_7223);
or U7378 (N_7378,N_7002,N_7027);
nand U7379 (N_7379,N_7199,N_7085);
and U7380 (N_7380,N_7099,N_7240);
or U7381 (N_7381,N_7127,N_7248);
nor U7382 (N_7382,N_7022,N_7088);
and U7383 (N_7383,N_7190,N_7074);
nand U7384 (N_7384,N_7241,N_7176);
and U7385 (N_7385,N_7218,N_7216);
and U7386 (N_7386,N_7097,N_7083);
or U7387 (N_7387,N_7152,N_7191);
nor U7388 (N_7388,N_7226,N_7212);
and U7389 (N_7389,N_7101,N_7047);
nor U7390 (N_7390,N_7106,N_7153);
or U7391 (N_7391,N_7063,N_7045);
nor U7392 (N_7392,N_7156,N_7040);
nor U7393 (N_7393,N_7141,N_7224);
and U7394 (N_7394,N_7062,N_7134);
or U7395 (N_7395,N_7073,N_7170);
or U7396 (N_7396,N_7053,N_7238);
or U7397 (N_7397,N_7141,N_7199);
nor U7398 (N_7398,N_7248,N_7165);
nor U7399 (N_7399,N_7011,N_7214);
nor U7400 (N_7400,N_7083,N_7129);
nor U7401 (N_7401,N_7018,N_7050);
nor U7402 (N_7402,N_7229,N_7000);
and U7403 (N_7403,N_7214,N_7025);
and U7404 (N_7404,N_7071,N_7001);
or U7405 (N_7405,N_7107,N_7138);
or U7406 (N_7406,N_7220,N_7092);
xor U7407 (N_7407,N_7068,N_7069);
xnor U7408 (N_7408,N_7024,N_7087);
nor U7409 (N_7409,N_7234,N_7056);
and U7410 (N_7410,N_7008,N_7054);
nand U7411 (N_7411,N_7073,N_7221);
or U7412 (N_7412,N_7190,N_7101);
or U7413 (N_7413,N_7153,N_7193);
nor U7414 (N_7414,N_7180,N_7188);
or U7415 (N_7415,N_7079,N_7049);
nand U7416 (N_7416,N_7197,N_7101);
xnor U7417 (N_7417,N_7238,N_7201);
and U7418 (N_7418,N_7109,N_7183);
or U7419 (N_7419,N_7228,N_7021);
or U7420 (N_7420,N_7102,N_7181);
nor U7421 (N_7421,N_7096,N_7014);
nand U7422 (N_7422,N_7074,N_7183);
nand U7423 (N_7423,N_7105,N_7207);
nand U7424 (N_7424,N_7238,N_7152);
nand U7425 (N_7425,N_7005,N_7135);
nand U7426 (N_7426,N_7081,N_7039);
nor U7427 (N_7427,N_7177,N_7051);
xor U7428 (N_7428,N_7110,N_7002);
and U7429 (N_7429,N_7142,N_7003);
or U7430 (N_7430,N_7115,N_7203);
nand U7431 (N_7431,N_7052,N_7055);
nand U7432 (N_7432,N_7038,N_7060);
nand U7433 (N_7433,N_7113,N_7070);
and U7434 (N_7434,N_7233,N_7141);
nand U7435 (N_7435,N_7156,N_7201);
and U7436 (N_7436,N_7219,N_7007);
and U7437 (N_7437,N_7065,N_7246);
or U7438 (N_7438,N_7189,N_7067);
nor U7439 (N_7439,N_7142,N_7085);
nor U7440 (N_7440,N_7205,N_7122);
or U7441 (N_7441,N_7213,N_7117);
and U7442 (N_7442,N_7201,N_7155);
or U7443 (N_7443,N_7079,N_7038);
and U7444 (N_7444,N_7123,N_7115);
and U7445 (N_7445,N_7136,N_7033);
and U7446 (N_7446,N_7063,N_7231);
or U7447 (N_7447,N_7190,N_7181);
and U7448 (N_7448,N_7068,N_7168);
or U7449 (N_7449,N_7238,N_7039);
or U7450 (N_7450,N_7049,N_7233);
and U7451 (N_7451,N_7029,N_7121);
nand U7452 (N_7452,N_7151,N_7169);
or U7453 (N_7453,N_7181,N_7242);
nor U7454 (N_7454,N_7081,N_7203);
nand U7455 (N_7455,N_7220,N_7043);
or U7456 (N_7456,N_7047,N_7005);
nor U7457 (N_7457,N_7110,N_7172);
or U7458 (N_7458,N_7193,N_7057);
or U7459 (N_7459,N_7210,N_7177);
nor U7460 (N_7460,N_7138,N_7002);
and U7461 (N_7461,N_7017,N_7103);
or U7462 (N_7462,N_7219,N_7239);
and U7463 (N_7463,N_7106,N_7200);
and U7464 (N_7464,N_7189,N_7223);
or U7465 (N_7465,N_7110,N_7234);
or U7466 (N_7466,N_7071,N_7002);
or U7467 (N_7467,N_7245,N_7180);
or U7468 (N_7468,N_7217,N_7171);
xnor U7469 (N_7469,N_7075,N_7181);
and U7470 (N_7470,N_7081,N_7208);
and U7471 (N_7471,N_7190,N_7025);
nand U7472 (N_7472,N_7176,N_7065);
nor U7473 (N_7473,N_7140,N_7216);
and U7474 (N_7474,N_7220,N_7167);
nand U7475 (N_7475,N_7086,N_7209);
and U7476 (N_7476,N_7187,N_7037);
nor U7477 (N_7477,N_7013,N_7080);
nand U7478 (N_7478,N_7120,N_7208);
or U7479 (N_7479,N_7007,N_7082);
nand U7480 (N_7480,N_7191,N_7142);
nand U7481 (N_7481,N_7167,N_7076);
nor U7482 (N_7482,N_7017,N_7211);
and U7483 (N_7483,N_7125,N_7072);
and U7484 (N_7484,N_7214,N_7171);
and U7485 (N_7485,N_7065,N_7170);
or U7486 (N_7486,N_7114,N_7167);
and U7487 (N_7487,N_7212,N_7129);
nor U7488 (N_7488,N_7215,N_7199);
nand U7489 (N_7489,N_7156,N_7079);
or U7490 (N_7490,N_7101,N_7064);
and U7491 (N_7491,N_7244,N_7192);
xor U7492 (N_7492,N_7189,N_7005);
or U7493 (N_7493,N_7060,N_7113);
or U7494 (N_7494,N_7184,N_7160);
nor U7495 (N_7495,N_7127,N_7173);
or U7496 (N_7496,N_7207,N_7059);
or U7497 (N_7497,N_7241,N_7128);
nor U7498 (N_7498,N_7148,N_7104);
nor U7499 (N_7499,N_7213,N_7054);
and U7500 (N_7500,N_7272,N_7403);
and U7501 (N_7501,N_7326,N_7370);
or U7502 (N_7502,N_7349,N_7319);
nand U7503 (N_7503,N_7427,N_7499);
or U7504 (N_7504,N_7463,N_7454);
xnor U7505 (N_7505,N_7285,N_7381);
nand U7506 (N_7506,N_7417,N_7460);
or U7507 (N_7507,N_7447,N_7317);
nor U7508 (N_7508,N_7462,N_7306);
and U7509 (N_7509,N_7377,N_7327);
or U7510 (N_7510,N_7257,N_7281);
nor U7511 (N_7511,N_7411,N_7428);
nor U7512 (N_7512,N_7311,N_7414);
and U7513 (N_7513,N_7290,N_7404);
nor U7514 (N_7514,N_7343,N_7416);
nand U7515 (N_7515,N_7400,N_7340);
nand U7516 (N_7516,N_7379,N_7264);
and U7517 (N_7517,N_7421,N_7487);
xor U7518 (N_7518,N_7456,N_7358);
nand U7519 (N_7519,N_7347,N_7333);
nor U7520 (N_7520,N_7442,N_7321);
nor U7521 (N_7521,N_7424,N_7284);
and U7522 (N_7522,N_7304,N_7483);
and U7523 (N_7523,N_7301,N_7478);
nor U7524 (N_7524,N_7318,N_7369);
nand U7525 (N_7525,N_7313,N_7291);
nand U7526 (N_7526,N_7316,N_7477);
and U7527 (N_7527,N_7361,N_7455);
or U7528 (N_7528,N_7328,N_7268);
nand U7529 (N_7529,N_7394,N_7299);
or U7530 (N_7530,N_7367,N_7375);
nand U7531 (N_7531,N_7498,N_7443);
nand U7532 (N_7532,N_7439,N_7265);
and U7533 (N_7533,N_7386,N_7325);
and U7534 (N_7534,N_7354,N_7279);
and U7535 (N_7535,N_7280,N_7338);
nand U7536 (N_7536,N_7276,N_7310);
nand U7537 (N_7537,N_7429,N_7438);
nor U7538 (N_7538,N_7362,N_7385);
nand U7539 (N_7539,N_7436,N_7382);
or U7540 (N_7540,N_7351,N_7300);
or U7541 (N_7541,N_7465,N_7292);
nand U7542 (N_7542,N_7485,N_7355);
nand U7543 (N_7543,N_7479,N_7302);
nand U7544 (N_7544,N_7263,N_7359);
nor U7545 (N_7545,N_7278,N_7261);
nand U7546 (N_7546,N_7378,N_7345);
nor U7547 (N_7547,N_7446,N_7476);
and U7548 (N_7548,N_7346,N_7286);
and U7549 (N_7549,N_7356,N_7474);
nand U7550 (N_7550,N_7252,N_7352);
and U7551 (N_7551,N_7402,N_7374);
nor U7552 (N_7552,N_7398,N_7387);
xor U7553 (N_7553,N_7357,N_7255);
or U7554 (N_7554,N_7256,N_7266);
nor U7555 (N_7555,N_7419,N_7467);
nor U7556 (N_7556,N_7253,N_7481);
and U7557 (N_7557,N_7434,N_7344);
and U7558 (N_7558,N_7287,N_7295);
and U7559 (N_7559,N_7409,N_7408);
and U7560 (N_7560,N_7492,N_7453);
nand U7561 (N_7561,N_7469,N_7405);
and U7562 (N_7562,N_7293,N_7431);
and U7563 (N_7563,N_7353,N_7360);
and U7564 (N_7564,N_7273,N_7277);
or U7565 (N_7565,N_7488,N_7372);
nand U7566 (N_7566,N_7399,N_7380);
nand U7567 (N_7567,N_7373,N_7461);
or U7568 (N_7568,N_7486,N_7441);
and U7569 (N_7569,N_7475,N_7466);
xor U7570 (N_7570,N_7395,N_7258);
nand U7571 (N_7571,N_7368,N_7297);
or U7572 (N_7572,N_7450,N_7412);
nor U7573 (N_7573,N_7298,N_7271);
and U7574 (N_7574,N_7432,N_7480);
and U7575 (N_7575,N_7496,N_7471);
nor U7576 (N_7576,N_7384,N_7322);
nor U7577 (N_7577,N_7420,N_7444);
and U7578 (N_7578,N_7388,N_7350);
or U7579 (N_7579,N_7335,N_7376);
nand U7580 (N_7580,N_7459,N_7296);
or U7581 (N_7581,N_7342,N_7445);
nand U7582 (N_7582,N_7371,N_7490);
or U7583 (N_7583,N_7440,N_7294);
and U7584 (N_7584,N_7425,N_7423);
and U7585 (N_7585,N_7307,N_7314);
xor U7586 (N_7586,N_7418,N_7449);
nor U7587 (N_7587,N_7391,N_7435);
nand U7588 (N_7588,N_7267,N_7426);
and U7589 (N_7589,N_7348,N_7288);
and U7590 (N_7590,N_7329,N_7303);
nand U7591 (N_7591,N_7495,N_7482);
nor U7592 (N_7592,N_7366,N_7308);
nand U7593 (N_7593,N_7275,N_7392);
nor U7594 (N_7594,N_7383,N_7312);
nand U7595 (N_7595,N_7254,N_7330);
and U7596 (N_7596,N_7259,N_7282);
nand U7597 (N_7597,N_7397,N_7415);
nand U7598 (N_7598,N_7472,N_7413);
nor U7599 (N_7599,N_7334,N_7464);
xor U7600 (N_7600,N_7457,N_7484);
or U7601 (N_7601,N_7491,N_7451);
and U7602 (N_7602,N_7393,N_7389);
or U7603 (N_7603,N_7262,N_7315);
or U7604 (N_7604,N_7433,N_7401);
and U7605 (N_7605,N_7363,N_7407);
or U7606 (N_7606,N_7260,N_7324);
or U7607 (N_7607,N_7406,N_7283);
and U7608 (N_7608,N_7390,N_7493);
and U7609 (N_7609,N_7250,N_7448);
and U7610 (N_7610,N_7331,N_7270);
and U7611 (N_7611,N_7274,N_7473);
and U7612 (N_7612,N_7305,N_7489);
or U7613 (N_7613,N_7396,N_7337);
or U7614 (N_7614,N_7468,N_7309);
or U7615 (N_7615,N_7365,N_7494);
and U7616 (N_7616,N_7364,N_7320);
nor U7617 (N_7617,N_7323,N_7341);
nor U7618 (N_7618,N_7470,N_7497);
or U7619 (N_7619,N_7452,N_7289);
or U7620 (N_7620,N_7422,N_7269);
and U7621 (N_7621,N_7339,N_7430);
nand U7622 (N_7622,N_7251,N_7410);
and U7623 (N_7623,N_7336,N_7458);
or U7624 (N_7624,N_7437,N_7332);
or U7625 (N_7625,N_7385,N_7265);
or U7626 (N_7626,N_7387,N_7492);
nor U7627 (N_7627,N_7392,N_7385);
nor U7628 (N_7628,N_7373,N_7410);
nand U7629 (N_7629,N_7265,N_7325);
and U7630 (N_7630,N_7362,N_7464);
or U7631 (N_7631,N_7458,N_7404);
and U7632 (N_7632,N_7419,N_7295);
and U7633 (N_7633,N_7455,N_7276);
or U7634 (N_7634,N_7300,N_7361);
or U7635 (N_7635,N_7280,N_7302);
nand U7636 (N_7636,N_7330,N_7292);
or U7637 (N_7637,N_7406,N_7301);
nor U7638 (N_7638,N_7422,N_7287);
nor U7639 (N_7639,N_7287,N_7257);
or U7640 (N_7640,N_7313,N_7495);
nor U7641 (N_7641,N_7313,N_7455);
or U7642 (N_7642,N_7274,N_7328);
nor U7643 (N_7643,N_7475,N_7293);
nor U7644 (N_7644,N_7270,N_7278);
nand U7645 (N_7645,N_7460,N_7397);
xor U7646 (N_7646,N_7486,N_7306);
nor U7647 (N_7647,N_7309,N_7413);
or U7648 (N_7648,N_7280,N_7403);
nand U7649 (N_7649,N_7256,N_7451);
nand U7650 (N_7650,N_7368,N_7257);
and U7651 (N_7651,N_7266,N_7448);
nor U7652 (N_7652,N_7480,N_7279);
nor U7653 (N_7653,N_7253,N_7494);
nand U7654 (N_7654,N_7264,N_7411);
or U7655 (N_7655,N_7432,N_7426);
or U7656 (N_7656,N_7489,N_7288);
nand U7657 (N_7657,N_7463,N_7411);
nor U7658 (N_7658,N_7325,N_7499);
nand U7659 (N_7659,N_7301,N_7293);
and U7660 (N_7660,N_7366,N_7293);
nand U7661 (N_7661,N_7319,N_7394);
or U7662 (N_7662,N_7336,N_7331);
or U7663 (N_7663,N_7363,N_7311);
or U7664 (N_7664,N_7279,N_7416);
and U7665 (N_7665,N_7342,N_7317);
or U7666 (N_7666,N_7256,N_7302);
or U7667 (N_7667,N_7381,N_7373);
nand U7668 (N_7668,N_7280,N_7394);
nand U7669 (N_7669,N_7431,N_7446);
or U7670 (N_7670,N_7471,N_7458);
nand U7671 (N_7671,N_7422,N_7480);
nor U7672 (N_7672,N_7377,N_7250);
nand U7673 (N_7673,N_7364,N_7367);
nand U7674 (N_7674,N_7478,N_7442);
or U7675 (N_7675,N_7295,N_7308);
nor U7676 (N_7676,N_7387,N_7346);
nor U7677 (N_7677,N_7399,N_7300);
nand U7678 (N_7678,N_7492,N_7375);
nand U7679 (N_7679,N_7449,N_7363);
nor U7680 (N_7680,N_7395,N_7253);
nand U7681 (N_7681,N_7304,N_7442);
or U7682 (N_7682,N_7300,N_7273);
nand U7683 (N_7683,N_7430,N_7288);
nor U7684 (N_7684,N_7300,N_7366);
nand U7685 (N_7685,N_7271,N_7420);
and U7686 (N_7686,N_7410,N_7384);
nand U7687 (N_7687,N_7483,N_7477);
nand U7688 (N_7688,N_7446,N_7433);
and U7689 (N_7689,N_7345,N_7322);
nand U7690 (N_7690,N_7352,N_7393);
nand U7691 (N_7691,N_7275,N_7489);
or U7692 (N_7692,N_7408,N_7350);
or U7693 (N_7693,N_7430,N_7469);
nor U7694 (N_7694,N_7311,N_7339);
nand U7695 (N_7695,N_7426,N_7473);
nor U7696 (N_7696,N_7284,N_7269);
or U7697 (N_7697,N_7251,N_7380);
nand U7698 (N_7698,N_7480,N_7387);
or U7699 (N_7699,N_7286,N_7281);
and U7700 (N_7700,N_7428,N_7371);
or U7701 (N_7701,N_7280,N_7423);
or U7702 (N_7702,N_7493,N_7355);
nor U7703 (N_7703,N_7262,N_7379);
xor U7704 (N_7704,N_7420,N_7414);
and U7705 (N_7705,N_7394,N_7457);
or U7706 (N_7706,N_7264,N_7461);
nor U7707 (N_7707,N_7398,N_7352);
nand U7708 (N_7708,N_7280,N_7323);
nand U7709 (N_7709,N_7335,N_7427);
or U7710 (N_7710,N_7256,N_7329);
or U7711 (N_7711,N_7273,N_7342);
or U7712 (N_7712,N_7405,N_7457);
or U7713 (N_7713,N_7321,N_7334);
and U7714 (N_7714,N_7357,N_7481);
and U7715 (N_7715,N_7277,N_7260);
nand U7716 (N_7716,N_7310,N_7457);
or U7717 (N_7717,N_7304,N_7347);
nor U7718 (N_7718,N_7415,N_7488);
nor U7719 (N_7719,N_7263,N_7262);
nand U7720 (N_7720,N_7268,N_7387);
nand U7721 (N_7721,N_7465,N_7383);
nor U7722 (N_7722,N_7494,N_7327);
and U7723 (N_7723,N_7482,N_7387);
nand U7724 (N_7724,N_7280,N_7416);
or U7725 (N_7725,N_7328,N_7495);
and U7726 (N_7726,N_7459,N_7466);
or U7727 (N_7727,N_7373,N_7379);
and U7728 (N_7728,N_7309,N_7499);
and U7729 (N_7729,N_7454,N_7374);
and U7730 (N_7730,N_7380,N_7369);
and U7731 (N_7731,N_7379,N_7439);
and U7732 (N_7732,N_7340,N_7280);
nor U7733 (N_7733,N_7454,N_7330);
and U7734 (N_7734,N_7295,N_7331);
nor U7735 (N_7735,N_7475,N_7348);
and U7736 (N_7736,N_7441,N_7304);
nor U7737 (N_7737,N_7423,N_7476);
nand U7738 (N_7738,N_7340,N_7342);
and U7739 (N_7739,N_7441,N_7335);
or U7740 (N_7740,N_7302,N_7293);
and U7741 (N_7741,N_7338,N_7296);
nor U7742 (N_7742,N_7324,N_7375);
nor U7743 (N_7743,N_7472,N_7485);
nand U7744 (N_7744,N_7303,N_7328);
nand U7745 (N_7745,N_7481,N_7497);
or U7746 (N_7746,N_7423,N_7327);
or U7747 (N_7747,N_7364,N_7343);
nor U7748 (N_7748,N_7406,N_7306);
nand U7749 (N_7749,N_7407,N_7449);
or U7750 (N_7750,N_7565,N_7500);
nor U7751 (N_7751,N_7630,N_7635);
or U7752 (N_7752,N_7584,N_7554);
nand U7753 (N_7753,N_7684,N_7700);
nor U7754 (N_7754,N_7509,N_7605);
nor U7755 (N_7755,N_7691,N_7716);
or U7756 (N_7756,N_7532,N_7632);
nor U7757 (N_7757,N_7693,N_7662);
nand U7758 (N_7758,N_7588,N_7510);
xor U7759 (N_7759,N_7613,N_7521);
and U7760 (N_7760,N_7661,N_7671);
or U7761 (N_7761,N_7650,N_7653);
nor U7762 (N_7762,N_7525,N_7651);
and U7763 (N_7763,N_7726,N_7604);
nor U7764 (N_7764,N_7522,N_7536);
nand U7765 (N_7765,N_7520,N_7595);
or U7766 (N_7766,N_7713,N_7699);
or U7767 (N_7767,N_7586,N_7637);
nand U7768 (N_7768,N_7591,N_7593);
nand U7769 (N_7769,N_7569,N_7687);
and U7770 (N_7770,N_7608,N_7672);
nor U7771 (N_7771,N_7545,N_7623);
nor U7772 (N_7772,N_7643,N_7704);
nand U7773 (N_7773,N_7535,N_7534);
and U7774 (N_7774,N_7703,N_7668);
and U7775 (N_7775,N_7677,N_7607);
nand U7776 (N_7776,N_7701,N_7705);
nand U7777 (N_7777,N_7616,N_7567);
or U7778 (N_7778,N_7743,N_7720);
and U7779 (N_7779,N_7559,N_7737);
and U7780 (N_7780,N_7746,N_7528);
or U7781 (N_7781,N_7731,N_7621);
nor U7782 (N_7782,N_7537,N_7736);
and U7783 (N_7783,N_7708,N_7640);
nand U7784 (N_7784,N_7560,N_7549);
nor U7785 (N_7785,N_7652,N_7572);
nand U7786 (N_7786,N_7527,N_7624);
or U7787 (N_7787,N_7678,N_7542);
nand U7788 (N_7788,N_7690,N_7502);
nor U7789 (N_7789,N_7666,N_7694);
nor U7790 (N_7790,N_7501,N_7550);
and U7791 (N_7791,N_7524,N_7642);
or U7792 (N_7792,N_7599,N_7709);
nand U7793 (N_7793,N_7507,N_7674);
nand U7794 (N_7794,N_7739,N_7626);
nor U7795 (N_7795,N_7552,N_7629);
or U7796 (N_7796,N_7675,N_7742);
or U7797 (N_7797,N_7654,N_7740);
nand U7798 (N_7798,N_7513,N_7646);
and U7799 (N_7799,N_7574,N_7617);
nor U7800 (N_7800,N_7628,N_7614);
and U7801 (N_7801,N_7619,N_7538);
nand U7802 (N_7802,N_7667,N_7540);
and U7803 (N_7803,N_7663,N_7648);
nor U7804 (N_7804,N_7680,N_7719);
nor U7805 (N_7805,N_7573,N_7717);
nor U7806 (N_7806,N_7634,N_7715);
or U7807 (N_7807,N_7610,N_7718);
and U7808 (N_7808,N_7683,N_7681);
nand U7809 (N_7809,N_7689,N_7585);
and U7810 (N_7810,N_7644,N_7732);
and U7811 (N_7811,N_7695,N_7733);
xor U7812 (N_7812,N_7696,N_7548);
and U7813 (N_7813,N_7529,N_7566);
and U7814 (N_7814,N_7673,N_7580);
nor U7815 (N_7815,N_7505,N_7639);
nand U7816 (N_7816,N_7658,N_7575);
nor U7817 (N_7817,N_7656,N_7725);
and U7818 (N_7818,N_7557,N_7508);
and U7819 (N_7819,N_7601,N_7546);
or U7820 (N_7820,N_7747,N_7721);
nand U7821 (N_7821,N_7512,N_7581);
nand U7822 (N_7822,N_7697,N_7612);
and U7823 (N_7823,N_7749,N_7597);
and U7824 (N_7824,N_7519,N_7636);
or U7825 (N_7825,N_7564,N_7609);
xnor U7826 (N_7826,N_7523,N_7543);
xnor U7827 (N_7827,N_7741,N_7723);
and U7828 (N_7828,N_7657,N_7511);
nor U7829 (N_7829,N_7638,N_7526);
and U7830 (N_7830,N_7665,N_7647);
and U7831 (N_7831,N_7531,N_7506);
nor U7832 (N_7832,N_7539,N_7551);
nand U7833 (N_7833,N_7603,N_7576);
and U7834 (N_7834,N_7633,N_7562);
and U7835 (N_7835,N_7714,N_7724);
nand U7836 (N_7836,N_7606,N_7711);
nand U7837 (N_7837,N_7504,N_7579);
nand U7838 (N_7838,N_7515,N_7730);
nand U7839 (N_7839,N_7533,N_7707);
nand U7840 (N_7840,N_7571,N_7517);
and U7841 (N_7841,N_7649,N_7602);
nand U7842 (N_7842,N_7611,N_7706);
or U7843 (N_7843,N_7556,N_7702);
or U7844 (N_7844,N_7570,N_7547);
or U7845 (N_7845,N_7745,N_7600);
or U7846 (N_7846,N_7738,N_7660);
or U7847 (N_7847,N_7592,N_7686);
and U7848 (N_7848,N_7748,N_7555);
nand U7849 (N_7849,N_7553,N_7530);
and U7850 (N_7850,N_7582,N_7561);
nand U7851 (N_7851,N_7729,N_7728);
or U7852 (N_7852,N_7655,N_7578);
nor U7853 (N_7853,N_7710,N_7735);
and U7854 (N_7854,N_7676,N_7627);
or U7855 (N_7855,N_7688,N_7563);
nor U7856 (N_7856,N_7558,N_7670);
and U7857 (N_7857,N_7590,N_7615);
or U7858 (N_7858,N_7568,N_7685);
or U7859 (N_7859,N_7503,N_7682);
and U7860 (N_7860,N_7577,N_7625);
and U7861 (N_7861,N_7712,N_7544);
nor U7862 (N_7862,N_7598,N_7692);
nor U7863 (N_7863,N_7618,N_7744);
and U7864 (N_7864,N_7587,N_7727);
and U7865 (N_7865,N_7641,N_7664);
nand U7866 (N_7866,N_7516,N_7645);
or U7867 (N_7867,N_7669,N_7698);
nor U7868 (N_7868,N_7631,N_7659);
and U7869 (N_7869,N_7620,N_7589);
nand U7870 (N_7870,N_7734,N_7679);
or U7871 (N_7871,N_7622,N_7594);
nand U7872 (N_7872,N_7518,N_7514);
and U7873 (N_7873,N_7541,N_7583);
nand U7874 (N_7874,N_7596,N_7722);
nor U7875 (N_7875,N_7648,N_7733);
nand U7876 (N_7876,N_7721,N_7577);
and U7877 (N_7877,N_7626,N_7517);
nand U7878 (N_7878,N_7525,N_7578);
nand U7879 (N_7879,N_7689,N_7512);
nor U7880 (N_7880,N_7600,N_7626);
nand U7881 (N_7881,N_7525,N_7699);
nor U7882 (N_7882,N_7542,N_7588);
xnor U7883 (N_7883,N_7515,N_7560);
nor U7884 (N_7884,N_7576,N_7632);
nor U7885 (N_7885,N_7533,N_7532);
or U7886 (N_7886,N_7600,N_7696);
nor U7887 (N_7887,N_7727,N_7621);
and U7888 (N_7888,N_7677,N_7575);
and U7889 (N_7889,N_7644,N_7609);
or U7890 (N_7890,N_7676,N_7547);
nor U7891 (N_7891,N_7590,N_7653);
and U7892 (N_7892,N_7673,N_7717);
nand U7893 (N_7893,N_7516,N_7515);
or U7894 (N_7894,N_7627,N_7733);
nor U7895 (N_7895,N_7546,N_7747);
xor U7896 (N_7896,N_7676,N_7536);
nand U7897 (N_7897,N_7512,N_7505);
nor U7898 (N_7898,N_7734,N_7622);
nand U7899 (N_7899,N_7600,N_7622);
nand U7900 (N_7900,N_7727,N_7533);
and U7901 (N_7901,N_7738,N_7714);
nand U7902 (N_7902,N_7725,N_7677);
and U7903 (N_7903,N_7626,N_7502);
nor U7904 (N_7904,N_7581,N_7648);
or U7905 (N_7905,N_7524,N_7670);
and U7906 (N_7906,N_7555,N_7655);
nor U7907 (N_7907,N_7571,N_7508);
nor U7908 (N_7908,N_7531,N_7697);
nor U7909 (N_7909,N_7664,N_7556);
or U7910 (N_7910,N_7649,N_7542);
and U7911 (N_7911,N_7618,N_7712);
and U7912 (N_7912,N_7663,N_7698);
and U7913 (N_7913,N_7633,N_7610);
and U7914 (N_7914,N_7691,N_7596);
nor U7915 (N_7915,N_7566,N_7540);
xor U7916 (N_7916,N_7591,N_7560);
or U7917 (N_7917,N_7705,N_7714);
nand U7918 (N_7918,N_7594,N_7674);
and U7919 (N_7919,N_7509,N_7622);
or U7920 (N_7920,N_7715,N_7670);
nand U7921 (N_7921,N_7551,N_7584);
nor U7922 (N_7922,N_7635,N_7673);
nor U7923 (N_7923,N_7705,N_7676);
and U7924 (N_7924,N_7669,N_7645);
nand U7925 (N_7925,N_7633,N_7501);
and U7926 (N_7926,N_7742,N_7560);
and U7927 (N_7927,N_7559,N_7631);
and U7928 (N_7928,N_7644,N_7561);
nor U7929 (N_7929,N_7729,N_7578);
and U7930 (N_7930,N_7608,N_7601);
nor U7931 (N_7931,N_7707,N_7715);
or U7932 (N_7932,N_7653,N_7724);
nand U7933 (N_7933,N_7689,N_7618);
nand U7934 (N_7934,N_7704,N_7705);
and U7935 (N_7935,N_7603,N_7708);
and U7936 (N_7936,N_7508,N_7728);
and U7937 (N_7937,N_7512,N_7621);
nor U7938 (N_7938,N_7745,N_7659);
nand U7939 (N_7939,N_7531,N_7594);
xnor U7940 (N_7940,N_7629,N_7720);
and U7941 (N_7941,N_7618,N_7720);
nand U7942 (N_7942,N_7707,N_7716);
and U7943 (N_7943,N_7627,N_7560);
and U7944 (N_7944,N_7604,N_7632);
and U7945 (N_7945,N_7684,N_7511);
nand U7946 (N_7946,N_7740,N_7562);
nor U7947 (N_7947,N_7629,N_7595);
and U7948 (N_7948,N_7513,N_7502);
or U7949 (N_7949,N_7545,N_7526);
nand U7950 (N_7950,N_7727,N_7502);
nor U7951 (N_7951,N_7562,N_7667);
nand U7952 (N_7952,N_7658,N_7685);
and U7953 (N_7953,N_7634,N_7737);
nand U7954 (N_7954,N_7505,N_7632);
or U7955 (N_7955,N_7681,N_7538);
and U7956 (N_7956,N_7653,N_7647);
nor U7957 (N_7957,N_7641,N_7691);
or U7958 (N_7958,N_7512,N_7554);
or U7959 (N_7959,N_7535,N_7690);
or U7960 (N_7960,N_7693,N_7694);
or U7961 (N_7961,N_7703,N_7528);
nand U7962 (N_7962,N_7720,N_7563);
and U7963 (N_7963,N_7549,N_7641);
or U7964 (N_7964,N_7654,N_7563);
or U7965 (N_7965,N_7569,N_7742);
nand U7966 (N_7966,N_7728,N_7541);
nor U7967 (N_7967,N_7691,N_7608);
and U7968 (N_7968,N_7575,N_7602);
or U7969 (N_7969,N_7729,N_7576);
or U7970 (N_7970,N_7628,N_7692);
nand U7971 (N_7971,N_7548,N_7590);
nand U7972 (N_7972,N_7533,N_7548);
or U7973 (N_7973,N_7514,N_7505);
or U7974 (N_7974,N_7671,N_7637);
nor U7975 (N_7975,N_7659,N_7648);
or U7976 (N_7976,N_7715,N_7722);
and U7977 (N_7977,N_7516,N_7711);
nand U7978 (N_7978,N_7584,N_7700);
nor U7979 (N_7979,N_7552,N_7641);
or U7980 (N_7980,N_7638,N_7737);
and U7981 (N_7981,N_7620,N_7717);
nand U7982 (N_7982,N_7531,N_7629);
and U7983 (N_7983,N_7652,N_7547);
nand U7984 (N_7984,N_7710,N_7679);
nand U7985 (N_7985,N_7624,N_7606);
and U7986 (N_7986,N_7660,N_7580);
nand U7987 (N_7987,N_7557,N_7558);
nand U7988 (N_7988,N_7721,N_7643);
or U7989 (N_7989,N_7549,N_7707);
and U7990 (N_7990,N_7592,N_7683);
and U7991 (N_7991,N_7677,N_7628);
or U7992 (N_7992,N_7559,N_7602);
nor U7993 (N_7993,N_7576,N_7641);
nor U7994 (N_7994,N_7506,N_7703);
nor U7995 (N_7995,N_7704,N_7579);
and U7996 (N_7996,N_7582,N_7612);
nor U7997 (N_7997,N_7644,N_7511);
and U7998 (N_7998,N_7698,N_7735);
and U7999 (N_7999,N_7529,N_7637);
or U8000 (N_8000,N_7854,N_7895);
nand U8001 (N_8001,N_7842,N_7860);
or U8002 (N_8002,N_7777,N_7846);
nand U8003 (N_8003,N_7814,N_7967);
or U8004 (N_8004,N_7843,N_7824);
and U8005 (N_8005,N_7801,N_7912);
or U8006 (N_8006,N_7856,N_7831);
nand U8007 (N_8007,N_7828,N_7980);
nand U8008 (N_8008,N_7813,N_7809);
nand U8009 (N_8009,N_7753,N_7780);
nand U8010 (N_8010,N_7888,N_7838);
nand U8011 (N_8011,N_7858,N_7887);
and U8012 (N_8012,N_7876,N_7865);
or U8013 (N_8013,N_7982,N_7821);
nand U8014 (N_8014,N_7944,N_7919);
nand U8015 (N_8015,N_7981,N_7805);
nand U8016 (N_8016,N_7991,N_7788);
and U8017 (N_8017,N_7841,N_7771);
nand U8018 (N_8018,N_7953,N_7752);
and U8019 (N_8019,N_7815,N_7884);
nand U8020 (N_8020,N_7959,N_7983);
and U8021 (N_8021,N_7794,N_7978);
and U8022 (N_8022,N_7871,N_7907);
nor U8023 (N_8023,N_7826,N_7800);
nand U8024 (N_8024,N_7762,N_7774);
or U8025 (N_8025,N_7807,N_7974);
nand U8026 (N_8026,N_7881,N_7941);
nand U8027 (N_8027,N_7761,N_7916);
and U8028 (N_8028,N_7885,N_7882);
or U8029 (N_8029,N_7797,N_7954);
nor U8030 (N_8030,N_7866,N_7886);
or U8031 (N_8031,N_7950,N_7853);
nand U8032 (N_8032,N_7823,N_7946);
or U8033 (N_8033,N_7973,N_7966);
nor U8034 (N_8034,N_7785,N_7986);
nor U8035 (N_8035,N_7851,N_7963);
and U8036 (N_8036,N_7929,N_7874);
nand U8037 (N_8037,N_7905,N_7808);
nand U8038 (N_8038,N_7879,N_7911);
nand U8039 (N_8039,N_7918,N_7931);
or U8040 (N_8040,N_7934,N_7909);
or U8041 (N_8041,N_7758,N_7868);
nand U8042 (N_8042,N_7971,N_7837);
nor U8043 (N_8043,N_7773,N_7812);
nor U8044 (N_8044,N_7993,N_7751);
nand U8045 (N_8045,N_7827,N_7822);
nor U8046 (N_8046,N_7811,N_7772);
xnor U8047 (N_8047,N_7962,N_7817);
nand U8048 (N_8048,N_7952,N_7880);
and U8049 (N_8049,N_7775,N_7975);
nand U8050 (N_8050,N_7913,N_7917);
nor U8051 (N_8051,N_7786,N_7940);
nor U8052 (N_8052,N_7850,N_7898);
nor U8053 (N_8053,N_7901,N_7765);
nor U8054 (N_8054,N_7987,N_7942);
nand U8055 (N_8055,N_7960,N_7989);
nor U8056 (N_8056,N_7789,N_7939);
or U8057 (N_8057,N_7859,N_7755);
or U8058 (N_8058,N_7922,N_7764);
nand U8059 (N_8059,N_7829,N_7903);
or U8060 (N_8060,N_7985,N_7867);
nand U8061 (N_8061,N_7900,N_7820);
nand U8062 (N_8062,N_7864,N_7924);
nand U8063 (N_8063,N_7995,N_7957);
nand U8064 (N_8064,N_7976,N_7969);
or U8065 (N_8065,N_7839,N_7862);
nand U8066 (N_8066,N_7872,N_7869);
nand U8067 (N_8067,N_7833,N_7943);
nand U8068 (N_8068,N_7908,N_7899);
or U8069 (N_8069,N_7926,N_7945);
nor U8070 (N_8070,N_7834,N_7877);
and U8071 (N_8071,N_7970,N_7766);
nor U8072 (N_8072,N_7921,N_7767);
nor U8073 (N_8073,N_7923,N_7855);
or U8074 (N_8074,N_7852,N_7795);
nor U8075 (N_8075,N_7818,N_7902);
nand U8076 (N_8076,N_7782,N_7798);
nand U8077 (N_8077,N_7878,N_7873);
nand U8078 (N_8078,N_7990,N_7896);
or U8079 (N_8079,N_7832,N_7897);
nor U8080 (N_8080,N_7769,N_7955);
or U8081 (N_8081,N_7784,N_7998);
nor U8082 (N_8082,N_7870,N_7948);
nand U8083 (N_8083,N_7875,N_7927);
nor U8084 (N_8084,N_7810,N_7793);
nor U8085 (N_8085,N_7906,N_7933);
nor U8086 (N_8086,N_7894,N_7979);
and U8087 (N_8087,N_7750,N_7996);
or U8088 (N_8088,N_7935,N_7863);
nor U8089 (N_8089,N_7891,N_7792);
or U8090 (N_8090,N_7763,N_7988);
nand U8091 (N_8091,N_7779,N_7968);
nand U8092 (N_8092,N_7791,N_7778);
and U8093 (N_8093,N_7892,N_7890);
and U8094 (N_8094,N_7893,N_7925);
nor U8095 (N_8095,N_7760,N_7849);
nor U8096 (N_8096,N_7883,N_7857);
or U8097 (N_8097,N_7759,N_7787);
nor U8098 (N_8098,N_7836,N_7757);
nor U8099 (N_8099,N_7848,N_7756);
or U8100 (N_8100,N_7847,N_7958);
nor U8101 (N_8101,N_7781,N_7951);
or U8102 (N_8102,N_7889,N_7936);
nor U8103 (N_8103,N_7910,N_7915);
and U8104 (N_8104,N_7796,N_7776);
and U8105 (N_8105,N_7816,N_7972);
or U8106 (N_8106,N_7799,N_7845);
or U8107 (N_8107,N_7844,N_7992);
and U8108 (N_8108,N_7754,N_7790);
nor U8109 (N_8109,N_7930,N_7840);
nand U8110 (N_8110,N_7932,N_7928);
and U8111 (N_8111,N_7861,N_7904);
nand U8112 (N_8112,N_7825,N_7804);
nand U8113 (N_8113,N_7937,N_7997);
or U8114 (N_8114,N_7977,N_7768);
or U8115 (N_8115,N_7802,N_7961);
xor U8116 (N_8116,N_7938,N_7819);
nor U8117 (N_8117,N_7964,N_7999);
and U8118 (N_8118,N_7783,N_7947);
or U8119 (N_8119,N_7965,N_7956);
and U8120 (N_8120,N_7835,N_7949);
nand U8121 (N_8121,N_7920,N_7806);
nor U8122 (N_8122,N_7984,N_7994);
or U8123 (N_8123,N_7770,N_7914);
and U8124 (N_8124,N_7803,N_7830);
nor U8125 (N_8125,N_7911,N_7789);
xor U8126 (N_8126,N_7771,N_7945);
nor U8127 (N_8127,N_7752,N_7885);
and U8128 (N_8128,N_7829,N_7955);
or U8129 (N_8129,N_7905,N_7953);
and U8130 (N_8130,N_7986,N_7765);
nand U8131 (N_8131,N_7954,N_7802);
and U8132 (N_8132,N_7890,N_7846);
nor U8133 (N_8133,N_7949,N_7992);
or U8134 (N_8134,N_7988,N_7876);
nor U8135 (N_8135,N_7826,N_7842);
and U8136 (N_8136,N_7804,N_7924);
or U8137 (N_8137,N_7808,N_7897);
nor U8138 (N_8138,N_7788,N_7763);
and U8139 (N_8139,N_7990,N_7857);
and U8140 (N_8140,N_7990,N_7989);
nor U8141 (N_8141,N_7756,N_7819);
nor U8142 (N_8142,N_7797,N_7757);
or U8143 (N_8143,N_7973,N_7833);
and U8144 (N_8144,N_7850,N_7931);
or U8145 (N_8145,N_7762,N_7896);
nor U8146 (N_8146,N_7987,N_7902);
or U8147 (N_8147,N_7863,N_7772);
and U8148 (N_8148,N_7943,N_7988);
or U8149 (N_8149,N_7944,N_7836);
nand U8150 (N_8150,N_7976,N_7884);
nor U8151 (N_8151,N_7992,N_7899);
and U8152 (N_8152,N_7852,N_7925);
or U8153 (N_8153,N_7891,N_7858);
nor U8154 (N_8154,N_7758,N_7804);
nor U8155 (N_8155,N_7976,N_7834);
or U8156 (N_8156,N_7805,N_7876);
xnor U8157 (N_8157,N_7788,N_7894);
and U8158 (N_8158,N_7988,N_7946);
and U8159 (N_8159,N_7879,N_7902);
and U8160 (N_8160,N_7926,N_7947);
and U8161 (N_8161,N_7840,N_7781);
nand U8162 (N_8162,N_7939,N_7773);
and U8163 (N_8163,N_7863,N_7876);
nand U8164 (N_8164,N_7777,N_7882);
nand U8165 (N_8165,N_7982,N_7990);
or U8166 (N_8166,N_7982,N_7795);
nor U8167 (N_8167,N_7809,N_7773);
nor U8168 (N_8168,N_7846,N_7857);
nor U8169 (N_8169,N_7826,N_7888);
and U8170 (N_8170,N_7986,N_7775);
and U8171 (N_8171,N_7825,N_7802);
and U8172 (N_8172,N_7919,N_7939);
nor U8173 (N_8173,N_7836,N_7964);
nor U8174 (N_8174,N_7843,N_7905);
xor U8175 (N_8175,N_7896,N_7874);
nand U8176 (N_8176,N_7808,N_7807);
nand U8177 (N_8177,N_7840,N_7867);
or U8178 (N_8178,N_7970,N_7759);
nor U8179 (N_8179,N_7906,N_7908);
nor U8180 (N_8180,N_7770,N_7793);
and U8181 (N_8181,N_7999,N_7985);
nor U8182 (N_8182,N_7949,N_7891);
nor U8183 (N_8183,N_7953,N_7961);
nor U8184 (N_8184,N_7966,N_7879);
and U8185 (N_8185,N_7792,N_7782);
nand U8186 (N_8186,N_7862,N_7879);
nor U8187 (N_8187,N_7975,N_7929);
nor U8188 (N_8188,N_7753,N_7904);
nor U8189 (N_8189,N_7823,N_7870);
nand U8190 (N_8190,N_7957,N_7978);
or U8191 (N_8191,N_7807,N_7861);
nand U8192 (N_8192,N_7861,N_7827);
nor U8193 (N_8193,N_7854,N_7754);
or U8194 (N_8194,N_7969,N_7951);
nor U8195 (N_8195,N_7782,N_7882);
and U8196 (N_8196,N_7838,N_7952);
and U8197 (N_8197,N_7783,N_7895);
or U8198 (N_8198,N_7949,N_7932);
nand U8199 (N_8199,N_7952,N_7755);
nand U8200 (N_8200,N_7768,N_7928);
nand U8201 (N_8201,N_7876,N_7943);
nor U8202 (N_8202,N_7856,N_7766);
nor U8203 (N_8203,N_7940,N_7938);
or U8204 (N_8204,N_7824,N_7996);
xnor U8205 (N_8205,N_7796,N_7827);
and U8206 (N_8206,N_7858,N_7965);
nor U8207 (N_8207,N_7872,N_7907);
and U8208 (N_8208,N_7996,N_7994);
and U8209 (N_8209,N_7929,N_7757);
and U8210 (N_8210,N_7894,N_7965);
nand U8211 (N_8211,N_7839,N_7932);
and U8212 (N_8212,N_7919,N_7823);
xor U8213 (N_8213,N_7907,N_7834);
nor U8214 (N_8214,N_7771,N_7847);
and U8215 (N_8215,N_7920,N_7788);
nand U8216 (N_8216,N_7836,N_7906);
or U8217 (N_8217,N_7758,N_7974);
nand U8218 (N_8218,N_7866,N_7994);
or U8219 (N_8219,N_7999,N_7812);
nand U8220 (N_8220,N_7752,N_7950);
or U8221 (N_8221,N_7755,N_7759);
nand U8222 (N_8222,N_7946,N_7843);
or U8223 (N_8223,N_7990,N_7870);
nor U8224 (N_8224,N_7812,N_7921);
and U8225 (N_8225,N_7852,N_7849);
nor U8226 (N_8226,N_7918,N_7976);
nand U8227 (N_8227,N_7754,N_7827);
or U8228 (N_8228,N_7994,N_7770);
nand U8229 (N_8229,N_7867,N_7818);
xor U8230 (N_8230,N_7834,N_7987);
or U8231 (N_8231,N_7977,N_7787);
and U8232 (N_8232,N_7768,N_7869);
nor U8233 (N_8233,N_7893,N_7944);
nand U8234 (N_8234,N_7770,N_7999);
or U8235 (N_8235,N_7846,N_7773);
nand U8236 (N_8236,N_7830,N_7974);
and U8237 (N_8237,N_7879,N_7920);
and U8238 (N_8238,N_7844,N_7896);
nor U8239 (N_8239,N_7853,N_7960);
nor U8240 (N_8240,N_7845,N_7917);
or U8241 (N_8241,N_7968,N_7925);
or U8242 (N_8242,N_7854,N_7884);
and U8243 (N_8243,N_7835,N_7828);
nor U8244 (N_8244,N_7891,N_7991);
or U8245 (N_8245,N_7750,N_7784);
and U8246 (N_8246,N_7771,N_7792);
and U8247 (N_8247,N_7914,N_7898);
nand U8248 (N_8248,N_7882,N_7964);
nor U8249 (N_8249,N_7859,N_7987);
and U8250 (N_8250,N_8247,N_8043);
nor U8251 (N_8251,N_8130,N_8208);
nand U8252 (N_8252,N_8095,N_8053);
and U8253 (N_8253,N_8142,N_8180);
nand U8254 (N_8254,N_8110,N_8038);
nor U8255 (N_8255,N_8115,N_8241);
nor U8256 (N_8256,N_8137,N_8139);
xor U8257 (N_8257,N_8222,N_8062);
nor U8258 (N_8258,N_8085,N_8188);
and U8259 (N_8259,N_8163,N_8172);
and U8260 (N_8260,N_8230,N_8225);
nand U8261 (N_8261,N_8133,N_8019);
nor U8262 (N_8262,N_8091,N_8217);
nand U8263 (N_8263,N_8081,N_8194);
and U8264 (N_8264,N_8226,N_8151);
or U8265 (N_8265,N_8202,N_8159);
nor U8266 (N_8266,N_8134,N_8145);
nand U8267 (N_8267,N_8213,N_8071);
nor U8268 (N_8268,N_8079,N_8068);
nand U8269 (N_8269,N_8032,N_8051);
or U8270 (N_8270,N_8209,N_8138);
nor U8271 (N_8271,N_8034,N_8146);
nor U8272 (N_8272,N_8047,N_8057);
or U8273 (N_8273,N_8177,N_8107);
and U8274 (N_8274,N_8195,N_8153);
or U8275 (N_8275,N_8129,N_8097);
and U8276 (N_8276,N_8244,N_8124);
xnor U8277 (N_8277,N_8132,N_8179);
nor U8278 (N_8278,N_8105,N_8144);
nor U8279 (N_8279,N_8212,N_8009);
and U8280 (N_8280,N_8196,N_8109);
nor U8281 (N_8281,N_8036,N_8100);
nand U8282 (N_8282,N_8223,N_8184);
or U8283 (N_8283,N_8096,N_8245);
nand U8284 (N_8284,N_8012,N_8084);
or U8285 (N_8285,N_8065,N_8067);
nand U8286 (N_8286,N_8122,N_8136);
or U8287 (N_8287,N_8198,N_8015);
nand U8288 (N_8288,N_8077,N_8089);
nor U8289 (N_8289,N_8014,N_8033);
nor U8290 (N_8290,N_8236,N_8157);
or U8291 (N_8291,N_8006,N_8117);
and U8292 (N_8292,N_8165,N_8182);
or U8293 (N_8293,N_8018,N_8114);
nor U8294 (N_8294,N_8126,N_8017);
and U8295 (N_8295,N_8169,N_8123);
xnor U8296 (N_8296,N_8027,N_8049);
or U8297 (N_8297,N_8207,N_8078);
or U8298 (N_8298,N_8166,N_8238);
or U8299 (N_8299,N_8059,N_8023);
nand U8300 (N_8300,N_8200,N_8242);
and U8301 (N_8301,N_8003,N_8221);
nand U8302 (N_8302,N_8187,N_8025);
nor U8303 (N_8303,N_8204,N_8218);
or U8304 (N_8304,N_8060,N_8052);
nand U8305 (N_8305,N_8099,N_8041);
or U8306 (N_8306,N_8094,N_8080);
or U8307 (N_8307,N_8205,N_8227);
nor U8308 (N_8308,N_8073,N_8185);
and U8309 (N_8309,N_8090,N_8083);
or U8310 (N_8310,N_8149,N_8106);
xor U8311 (N_8311,N_8229,N_8183);
nand U8312 (N_8312,N_8008,N_8224);
or U8313 (N_8313,N_8013,N_8118);
and U8314 (N_8314,N_8040,N_8020);
nand U8315 (N_8315,N_8127,N_8055);
nor U8316 (N_8316,N_8181,N_8239);
xor U8317 (N_8317,N_8066,N_8178);
nor U8318 (N_8318,N_8190,N_8088);
nand U8319 (N_8319,N_8233,N_8193);
and U8320 (N_8320,N_8167,N_8037);
and U8321 (N_8321,N_8092,N_8050);
nor U8322 (N_8322,N_8243,N_8016);
and U8323 (N_8323,N_8143,N_8192);
and U8324 (N_8324,N_8064,N_8237);
and U8325 (N_8325,N_8155,N_8141);
or U8326 (N_8326,N_8168,N_8001);
nor U8327 (N_8327,N_8005,N_8199);
nand U8328 (N_8328,N_8219,N_8161);
and U8329 (N_8329,N_8069,N_8175);
nor U8330 (N_8330,N_8074,N_8216);
and U8331 (N_8331,N_8191,N_8021);
and U8332 (N_8332,N_8173,N_8240);
and U8333 (N_8333,N_8148,N_8054);
and U8334 (N_8334,N_8072,N_8087);
and U8335 (N_8335,N_8048,N_8170);
nand U8336 (N_8336,N_8022,N_8220);
and U8337 (N_8337,N_8004,N_8045);
or U8338 (N_8338,N_8000,N_8135);
or U8339 (N_8339,N_8171,N_8002);
xor U8340 (N_8340,N_8101,N_8160);
nand U8341 (N_8341,N_8056,N_8010);
or U8342 (N_8342,N_8112,N_8211);
xor U8343 (N_8343,N_8031,N_8058);
and U8344 (N_8344,N_8156,N_8120);
and U8345 (N_8345,N_8044,N_8150);
or U8346 (N_8346,N_8162,N_8075);
and U8347 (N_8347,N_8104,N_8024);
nor U8348 (N_8348,N_8206,N_8186);
nand U8349 (N_8349,N_8214,N_8039);
or U8350 (N_8350,N_8232,N_8108);
nor U8351 (N_8351,N_8076,N_8007);
or U8352 (N_8352,N_8234,N_8128);
or U8353 (N_8353,N_8035,N_8125);
nand U8354 (N_8354,N_8093,N_8116);
and U8355 (N_8355,N_8176,N_8046);
nor U8356 (N_8356,N_8197,N_8086);
nor U8357 (N_8357,N_8098,N_8131);
and U8358 (N_8358,N_8026,N_8140);
nand U8359 (N_8359,N_8174,N_8103);
and U8360 (N_8360,N_8121,N_8228);
and U8361 (N_8361,N_8029,N_8189);
nand U8362 (N_8362,N_8042,N_8063);
and U8363 (N_8363,N_8147,N_8201);
nor U8364 (N_8364,N_8011,N_8164);
and U8365 (N_8365,N_8154,N_8152);
nand U8366 (N_8366,N_8210,N_8215);
nor U8367 (N_8367,N_8235,N_8203);
or U8368 (N_8368,N_8102,N_8248);
or U8369 (N_8369,N_8246,N_8158);
or U8370 (N_8370,N_8119,N_8030);
or U8371 (N_8371,N_8061,N_8231);
xnor U8372 (N_8372,N_8082,N_8070);
nor U8373 (N_8373,N_8028,N_8249);
or U8374 (N_8374,N_8111,N_8113);
and U8375 (N_8375,N_8104,N_8041);
nor U8376 (N_8376,N_8061,N_8056);
and U8377 (N_8377,N_8138,N_8104);
and U8378 (N_8378,N_8199,N_8152);
or U8379 (N_8379,N_8093,N_8173);
or U8380 (N_8380,N_8123,N_8212);
or U8381 (N_8381,N_8047,N_8149);
or U8382 (N_8382,N_8169,N_8181);
and U8383 (N_8383,N_8238,N_8033);
or U8384 (N_8384,N_8191,N_8113);
or U8385 (N_8385,N_8083,N_8102);
nand U8386 (N_8386,N_8182,N_8214);
nor U8387 (N_8387,N_8091,N_8011);
and U8388 (N_8388,N_8191,N_8168);
nand U8389 (N_8389,N_8184,N_8203);
nand U8390 (N_8390,N_8051,N_8048);
nand U8391 (N_8391,N_8196,N_8242);
nor U8392 (N_8392,N_8218,N_8009);
nand U8393 (N_8393,N_8077,N_8058);
or U8394 (N_8394,N_8107,N_8085);
and U8395 (N_8395,N_8056,N_8193);
nand U8396 (N_8396,N_8115,N_8173);
or U8397 (N_8397,N_8077,N_8199);
or U8398 (N_8398,N_8066,N_8195);
or U8399 (N_8399,N_8014,N_8125);
or U8400 (N_8400,N_8157,N_8196);
nand U8401 (N_8401,N_8126,N_8013);
and U8402 (N_8402,N_8050,N_8128);
nand U8403 (N_8403,N_8121,N_8171);
nand U8404 (N_8404,N_8193,N_8170);
or U8405 (N_8405,N_8093,N_8209);
and U8406 (N_8406,N_8220,N_8014);
nand U8407 (N_8407,N_8146,N_8049);
nor U8408 (N_8408,N_8155,N_8028);
nand U8409 (N_8409,N_8099,N_8149);
nor U8410 (N_8410,N_8188,N_8100);
nand U8411 (N_8411,N_8137,N_8015);
and U8412 (N_8412,N_8155,N_8006);
nor U8413 (N_8413,N_8050,N_8192);
or U8414 (N_8414,N_8066,N_8054);
and U8415 (N_8415,N_8029,N_8091);
nor U8416 (N_8416,N_8165,N_8249);
nor U8417 (N_8417,N_8029,N_8225);
or U8418 (N_8418,N_8000,N_8193);
or U8419 (N_8419,N_8073,N_8088);
nand U8420 (N_8420,N_8086,N_8129);
and U8421 (N_8421,N_8013,N_8192);
or U8422 (N_8422,N_8101,N_8249);
nand U8423 (N_8423,N_8242,N_8152);
nor U8424 (N_8424,N_8191,N_8162);
nand U8425 (N_8425,N_8177,N_8055);
and U8426 (N_8426,N_8191,N_8142);
or U8427 (N_8427,N_8201,N_8149);
or U8428 (N_8428,N_8077,N_8134);
or U8429 (N_8429,N_8036,N_8216);
or U8430 (N_8430,N_8124,N_8135);
nand U8431 (N_8431,N_8191,N_8213);
or U8432 (N_8432,N_8121,N_8077);
nor U8433 (N_8433,N_8111,N_8122);
and U8434 (N_8434,N_8212,N_8238);
nand U8435 (N_8435,N_8212,N_8125);
and U8436 (N_8436,N_8146,N_8219);
nand U8437 (N_8437,N_8209,N_8122);
or U8438 (N_8438,N_8055,N_8079);
or U8439 (N_8439,N_8236,N_8127);
or U8440 (N_8440,N_8197,N_8241);
nand U8441 (N_8441,N_8115,N_8114);
nor U8442 (N_8442,N_8064,N_8232);
and U8443 (N_8443,N_8025,N_8235);
nand U8444 (N_8444,N_8074,N_8080);
nand U8445 (N_8445,N_8074,N_8244);
or U8446 (N_8446,N_8212,N_8037);
nor U8447 (N_8447,N_8176,N_8207);
and U8448 (N_8448,N_8184,N_8122);
or U8449 (N_8449,N_8043,N_8011);
nand U8450 (N_8450,N_8162,N_8114);
nor U8451 (N_8451,N_8187,N_8118);
or U8452 (N_8452,N_8211,N_8048);
nand U8453 (N_8453,N_8096,N_8242);
and U8454 (N_8454,N_8029,N_8049);
nor U8455 (N_8455,N_8072,N_8066);
nand U8456 (N_8456,N_8215,N_8080);
and U8457 (N_8457,N_8111,N_8046);
and U8458 (N_8458,N_8100,N_8193);
or U8459 (N_8459,N_8187,N_8240);
nand U8460 (N_8460,N_8169,N_8141);
or U8461 (N_8461,N_8236,N_8193);
and U8462 (N_8462,N_8179,N_8112);
and U8463 (N_8463,N_8162,N_8037);
and U8464 (N_8464,N_8029,N_8147);
and U8465 (N_8465,N_8150,N_8214);
and U8466 (N_8466,N_8232,N_8063);
nor U8467 (N_8467,N_8240,N_8079);
and U8468 (N_8468,N_8093,N_8062);
nand U8469 (N_8469,N_8154,N_8131);
xnor U8470 (N_8470,N_8238,N_8214);
and U8471 (N_8471,N_8008,N_8156);
or U8472 (N_8472,N_8057,N_8248);
nand U8473 (N_8473,N_8212,N_8081);
nor U8474 (N_8474,N_8208,N_8191);
nand U8475 (N_8475,N_8180,N_8171);
or U8476 (N_8476,N_8116,N_8232);
or U8477 (N_8477,N_8227,N_8156);
and U8478 (N_8478,N_8241,N_8173);
nand U8479 (N_8479,N_8164,N_8096);
nor U8480 (N_8480,N_8056,N_8007);
nand U8481 (N_8481,N_8246,N_8191);
or U8482 (N_8482,N_8218,N_8158);
nand U8483 (N_8483,N_8191,N_8017);
nor U8484 (N_8484,N_8052,N_8007);
and U8485 (N_8485,N_8032,N_8106);
nand U8486 (N_8486,N_8008,N_8163);
and U8487 (N_8487,N_8071,N_8086);
nor U8488 (N_8488,N_8015,N_8203);
nand U8489 (N_8489,N_8177,N_8101);
or U8490 (N_8490,N_8130,N_8025);
or U8491 (N_8491,N_8094,N_8177);
or U8492 (N_8492,N_8232,N_8103);
and U8493 (N_8493,N_8155,N_8072);
or U8494 (N_8494,N_8241,N_8165);
or U8495 (N_8495,N_8025,N_8023);
nand U8496 (N_8496,N_8098,N_8154);
or U8497 (N_8497,N_8074,N_8157);
nand U8498 (N_8498,N_8194,N_8159);
nand U8499 (N_8499,N_8213,N_8207);
or U8500 (N_8500,N_8445,N_8443);
nor U8501 (N_8501,N_8263,N_8359);
or U8502 (N_8502,N_8490,N_8414);
nor U8503 (N_8503,N_8396,N_8293);
xnor U8504 (N_8504,N_8413,N_8322);
nor U8505 (N_8505,N_8465,N_8300);
or U8506 (N_8506,N_8261,N_8323);
nor U8507 (N_8507,N_8495,N_8301);
nand U8508 (N_8508,N_8266,N_8402);
and U8509 (N_8509,N_8478,N_8365);
nor U8510 (N_8510,N_8388,N_8356);
nand U8511 (N_8511,N_8255,N_8376);
nor U8512 (N_8512,N_8307,N_8260);
nor U8513 (N_8513,N_8433,N_8363);
or U8514 (N_8514,N_8448,N_8308);
and U8515 (N_8515,N_8417,N_8406);
nor U8516 (N_8516,N_8277,N_8418);
and U8517 (N_8517,N_8434,N_8497);
nor U8518 (N_8518,N_8428,N_8367);
and U8519 (N_8519,N_8267,N_8390);
nand U8520 (N_8520,N_8327,N_8355);
or U8521 (N_8521,N_8253,N_8400);
nand U8522 (N_8522,N_8421,N_8286);
and U8523 (N_8523,N_8274,N_8262);
and U8524 (N_8524,N_8310,N_8462);
nor U8525 (N_8525,N_8362,N_8250);
and U8526 (N_8526,N_8299,N_8449);
nand U8527 (N_8527,N_8284,N_8389);
nand U8528 (N_8528,N_8252,N_8279);
xnor U8529 (N_8529,N_8473,N_8344);
nor U8530 (N_8530,N_8429,N_8387);
nor U8531 (N_8531,N_8306,N_8437);
nor U8532 (N_8532,N_8385,N_8334);
nor U8533 (N_8533,N_8394,N_8482);
nand U8534 (N_8534,N_8439,N_8460);
and U8535 (N_8535,N_8276,N_8316);
nor U8536 (N_8536,N_8283,N_8313);
or U8537 (N_8537,N_8487,N_8422);
and U8538 (N_8538,N_8412,N_8265);
nand U8539 (N_8539,N_8295,N_8351);
nor U8540 (N_8540,N_8494,N_8458);
nor U8541 (N_8541,N_8309,N_8288);
nor U8542 (N_8542,N_8304,N_8420);
nand U8543 (N_8543,N_8268,N_8453);
or U8544 (N_8544,N_8492,N_8264);
and U8545 (N_8545,N_8432,N_8319);
and U8546 (N_8546,N_8461,N_8446);
nand U8547 (N_8547,N_8383,N_8269);
or U8548 (N_8548,N_8399,N_8315);
or U8549 (N_8549,N_8426,N_8486);
and U8550 (N_8550,N_8484,N_8342);
nor U8551 (N_8551,N_8324,N_8350);
xnor U8552 (N_8552,N_8303,N_8290);
nor U8553 (N_8553,N_8404,N_8393);
and U8554 (N_8554,N_8476,N_8364);
or U8555 (N_8555,N_8401,N_8328);
nand U8556 (N_8556,N_8441,N_8357);
or U8557 (N_8557,N_8358,N_8361);
or U8558 (N_8558,N_8493,N_8371);
or U8559 (N_8559,N_8373,N_8257);
nand U8560 (N_8560,N_8331,N_8392);
or U8561 (N_8561,N_8477,N_8489);
or U8562 (N_8562,N_8294,N_8287);
nor U8563 (N_8563,N_8470,N_8272);
nand U8564 (N_8564,N_8353,N_8275);
nand U8565 (N_8565,N_8397,N_8410);
nor U8566 (N_8566,N_8280,N_8370);
or U8567 (N_8567,N_8326,N_8491);
nor U8568 (N_8568,N_8352,N_8498);
nand U8569 (N_8569,N_8488,N_8481);
nand U8570 (N_8570,N_8297,N_8440);
nor U8571 (N_8571,N_8474,N_8475);
nand U8572 (N_8572,N_8339,N_8338);
and U8573 (N_8573,N_8336,N_8403);
nand U8574 (N_8574,N_8292,N_8354);
nor U8575 (N_8575,N_8472,N_8348);
or U8576 (N_8576,N_8411,N_8471);
or U8577 (N_8577,N_8450,N_8291);
nor U8578 (N_8578,N_8374,N_8258);
nor U8579 (N_8579,N_8408,N_8395);
nand U8580 (N_8580,N_8464,N_8347);
nor U8581 (N_8581,N_8329,N_8271);
and U8582 (N_8582,N_8379,N_8337);
or U8583 (N_8583,N_8372,N_8270);
nor U8584 (N_8584,N_8431,N_8330);
or U8585 (N_8585,N_8427,N_8483);
nor U8586 (N_8586,N_8442,N_8479);
and U8587 (N_8587,N_8375,N_8377);
nand U8588 (N_8588,N_8282,N_8407);
and U8589 (N_8589,N_8451,N_8296);
or U8590 (N_8590,N_8466,N_8391);
nand U8591 (N_8591,N_8314,N_8368);
or U8592 (N_8592,N_8312,N_8318);
and U8593 (N_8593,N_8380,N_8321);
or U8594 (N_8594,N_8317,N_8278);
nor U8595 (N_8595,N_8468,N_8469);
and U8596 (N_8596,N_8333,N_8305);
nand U8597 (N_8597,N_8340,N_8384);
and U8598 (N_8598,N_8254,N_8405);
nand U8599 (N_8599,N_8447,N_8459);
and U8600 (N_8600,N_8463,N_8386);
nor U8601 (N_8601,N_8320,N_8341);
and U8602 (N_8602,N_8424,N_8281);
and U8603 (N_8603,N_8457,N_8298);
or U8604 (N_8604,N_8378,N_8423);
nor U8605 (N_8605,N_8369,N_8345);
or U8606 (N_8606,N_8302,N_8467);
nand U8607 (N_8607,N_8499,N_8381);
nor U8608 (N_8608,N_8256,N_8485);
nor U8609 (N_8609,N_8496,N_8456);
or U8610 (N_8610,N_8382,N_8360);
or U8611 (N_8611,N_8335,N_8454);
or U8612 (N_8612,N_8251,N_8325);
nor U8613 (N_8613,N_8425,N_8452);
and U8614 (N_8614,N_8415,N_8436);
nand U8615 (N_8615,N_8398,N_8435);
and U8616 (N_8616,N_8444,N_8273);
nand U8617 (N_8617,N_8409,N_8311);
nor U8618 (N_8618,N_8416,N_8346);
or U8619 (N_8619,N_8259,N_8349);
nor U8620 (N_8620,N_8419,N_8289);
nor U8621 (N_8621,N_8480,N_8438);
nor U8622 (N_8622,N_8455,N_8343);
and U8623 (N_8623,N_8430,N_8366);
and U8624 (N_8624,N_8285,N_8332);
and U8625 (N_8625,N_8376,N_8276);
or U8626 (N_8626,N_8419,N_8451);
or U8627 (N_8627,N_8309,N_8273);
or U8628 (N_8628,N_8337,N_8482);
or U8629 (N_8629,N_8377,N_8459);
nor U8630 (N_8630,N_8395,N_8391);
nor U8631 (N_8631,N_8373,N_8263);
nand U8632 (N_8632,N_8352,N_8404);
or U8633 (N_8633,N_8440,N_8390);
nand U8634 (N_8634,N_8362,N_8439);
nand U8635 (N_8635,N_8497,N_8324);
nor U8636 (N_8636,N_8253,N_8495);
or U8637 (N_8637,N_8366,N_8408);
and U8638 (N_8638,N_8405,N_8330);
or U8639 (N_8639,N_8276,N_8390);
or U8640 (N_8640,N_8274,N_8393);
and U8641 (N_8641,N_8405,N_8373);
and U8642 (N_8642,N_8313,N_8337);
and U8643 (N_8643,N_8360,N_8482);
or U8644 (N_8644,N_8305,N_8475);
nand U8645 (N_8645,N_8359,N_8418);
nand U8646 (N_8646,N_8400,N_8461);
and U8647 (N_8647,N_8396,N_8304);
nand U8648 (N_8648,N_8465,N_8261);
and U8649 (N_8649,N_8448,N_8322);
or U8650 (N_8650,N_8405,N_8412);
and U8651 (N_8651,N_8487,N_8489);
or U8652 (N_8652,N_8340,N_8468);
nand U8653 (N_8653,N_8279,N_8347);
nand U8654 (N_8654,N_8408,N_8471);
or U8655 (N_8655,N_8442,N_8293);
and U8656 (N_8656,N_8426,N_8256);
nand U8657 (N_8657,N_8471,N_8332);
and U8658 (N_8658,N_8330,N_8285);
and U8659 (N_8659,N_8467,N_8319);
or U8660 (N_8660,N_8408,N_8376);
and U8661 (N_8661,N_8335,N_8281);
nand U8662 (N_8662,N_8331,N_8311);
or U8663 (N_8663,N_8358,N_8312);
or U8664 (N_8664,N_8372,N_8492);
and U8665 (N_8665,N_8368,N_8269);
nor U8666 (N_8666,N_8376,N_8320);
or U8667 (N_8667,N_8462,N_8399);
nand U8668 (N_8668,N_8404,N_8256);
nand U8669 (N_8669,N_8292,N_8486);
nor U8670 (N_8670,N_8357,N_8462);
and U8671 (N_8671,N_8407,N_8279);
nand U8672 (N_8672,N_8361,N_8251);
or U8673 (N_8673,N_8309,N_8438);
or U8674 (N_8674,N_8406,N_8432);
and U8675 (N_8675,N_8288,N_8293);
or U8676 (N_8676,N_8375,N_8267);
nor U8677 (N_8677,N_8326,N_8315);
and U8678 (N_8678,N_8292,N_8375);
and U8679 (N_8679,N_8449,N_8269);
nor U8680 (N_8680,N_8334,N_8353);
and U8681 (N_8681,N_8479,N_8430);
nor U8682 (N_8682,N_8280,N_8314);
nand U8683 (N_8683,N_8419,N_8250);
or U8684 (N_8684,N_8328,N_8297);
nand U8685 (N_8685,N_8319,N_8476);
nor U8686 (N_8686,N_8370,N_8436);
or U8687 (N_8687,N_8440,N_8259);
nor U8688 (N_8688,N_8329,N_8327);
xnor U8689 (N_8689,N_8306,N_8377);
and U8690 (N_8690,N_8277,N_8262);
and U8691 (N_8691,N_8458,N_8417);
nand U8692 (N_8692,N_8408,N_8436);
and U8693 (N_8693,N_8433,N_8259);
and U8694 (N_8694,N_8487,N_8342);
xor U8695 (N_8695,N_8393,N_8315);
nand U8696 (N_8696,N_8359,N_8408);
or U8697 (N_8697,N_8348,N_8428);
and U8698 (N_8698,N_8485,N_8458);
or U8699 (N_8699,N_8258,N_8499);
nor U8700 (N_8700,N_8393,N_8330);
nor U8701 (N_8701,N_8362,N_8263);
nand U8702 (N_8702,N_8421,N_8345);
and U8703 (N_8703,N_8453,N_8456);
nand U8704 (N_8704,N_8278,N_8335);
and U8705 (N_8705,N_8493,N_8312);
nor U8706 (N_8706,N_8279,N_8312);
or U8707 (N_8707,N_8318,N_8362);
or U8708 (N_8708,N_8496,N_8484);
and U8709 (N_8709,N_8347,N_8498);
or U8710 (N_8710,N_8460,N_8355);
nand U8711 (N_8711,N_8316,N_8312);
xor U8712 (N_8712,N_8476,N_8467);
or U8713 (N_8713,N_8486,N_8269);
or U8714 (N_8714,N_8345,N_8488);
and U8715 (N_8715,N_8298,N_8396);
nor U8716 (N_8716,N_8478,N_8465);
or U8717 (N_8717,N_8434,N_8366);
or U8718 (N_8718,N_8342,N_8414);
or U8719 (N_8719,N_8450,N_8255);
and U8720 (N_8720,N_8491,N_8323);
or U8721 (N_8721,N_8280,N_8448);
nand U8722 (N_8722,N_8272,N_8488);
or U8723 (N_8723,N_8485,N_8491);
nor U8724 (N_8724,N_8465,N_8484);
or U8725 (N_8725,N_8313,N_8413);
and U8726 (N_8726,N_8423,N_8422);
and U8727 (N_8727,N_8428,N_8495);
nand U8728 (N_8728,N_8457,N_8417);
and U8729 (N_8729,N_8471,N_8328);
and U8730 (N_8730,N_8390,N_8476);
nand U8731 (N_8731,N_8370,N_8488);
nand U8732 (N_8732,N_8462,N_8385);
nand U8733 (N_8733,N_8288,N_8482);
or U8734 (N_8734,N_8378,N_8449);
and U8735 (N_8735,N_8420,N_8433);
and U8736 (N_8736,N_8271,N_8424);
nand U8737 (N_8737,N_8458,N_8462);
and U8738 (N_8738,N_8472,N_8487);
nor U8739 (N_8739,N_8423,N_8282);
and U8740 (N_8740,N_8458,N_8366);
nor U8741 (N_8741,N_8429,N_8317);
nor U8742 (N_8742,N_8256,N_8265);
nand U8743 (N_8743,N_8420,N_8297);
and U8744 (N_8744,N_8345,N_8440);
or U8745 (N_8745,N_8394,N_8356);
xor U8746 (N_8746,N_8465,N_8352);
nand U8747 (N_8747,N_8441,N_8338);
nor U8748 (N_8748,N_8457,N_8482);
nor U8749 (N_8749,N_8403,N_8416);
nand U8750 (N_8750,N_8688,N_8529);
nor U8751 (N_8751,N_8721,N_8503);
or U8752 (N_8752,N_8510,N_8728);
and U8753 (N_8753,N_8559,N_8674);
nor U8754 (N_8754,N_8689,N_8504);
nand U8755 (N_8755,N_8604,N_8725);
nor U8756 (N_8756,N_8702,N_8592);
nand U8757 (N_8757,N_8653,N_8623);
or U8758 (N_8758,N_8744,N_8556);
nor U8759 (N_8759,N_8703,N_8534);
nor U8760 (N_8760,N_8584,N_8745);
nor U8761 (N_8761,N_8566,N_8543);
nand U8762 (N_8762,N_8719,N_8730);
or U8763 (N_8763,N_8644,N_8746);
nand U8764 (N_8764,N_8572,N_8546);
or U8765 (N_8765,N_8642,N_8723);
and U8766 (N_8766,N_8588,N_8673);
nand U8767 (N_8767,N_8564,N_8562);
or U8768 (N_8768,N_8524,N_8538);
and U8769 (N_8769,N_8545,N_8657);
nand U8770 (N_8770,N_8722,N_8521);
and U8771 (N_8771,N_8511,N_8651);
and U8772 (N_8772,N_8732,N_8636);
nand U8773 (N_8773,N_8647,N_8551);
nor U8774 (N_8774,N_8549,N_8539);
xnor U8775 (N_8775,N_8649,N_8639);
nor U8776 (N_8776,N_8656,N_8720);
nor U8777 (N_8777,N_8669,N_8740);
and U8778 (N_8778,N_8571,N_8742);
and U8779 (N_8779,N_8668,N_8659);
xnor U8780 (N_8780,N_8518,N_8523);
or U8781 (N_8781,N_8747,N_8590);
nand U8782 (N_8782,N_8614,N_8563);
nand U8783 (N_8783,N_8617,N_8627);
nand U8784 (N_8784,N_8734,N_8696);
nand U8785 (N_8785,N_8569,N_8579);
and U8786 (N_8786,N_8519,N_8603);
or U8787 (N_8787,N_8692,N_8567);
or U8788 (N_8788,N_8568,N_8690);
nand U8789 (N_8789,N_8654,N_8535);
nor U8790 (N_8790,N_8516,N_8686);
and U8791 (N_8791,N_8502,N_8508);
nor U8792 (N_8792,N_8713,N_8514);
and U8793 (N_8793,N_8718,N_8607);
and U8794 (N_8794,N_8715,N_8735);
and U8795 (N_8795,N_8638,N_8698);
and U8796 (N_8796,N_8682,N_8678);
and U8797 (N_8797,N_8599,N_8550);
or U8798 (N_8798,N_8605,N_8600);
nor U8799 (N_8799,N_8573,N_8506);
or U8800 (N_8800,N_8611,N_8581);
or U8801 (N_8801,N_8711,N_8509);
nand U8802 (N_8802,N_8501,N_8741);
nand U8803 (N_8803,N_8641,N_8574);
nand U8804 (N_8804,N_8716,N_8706);
or U8805 (N_8805,N_8602,N_8632);
nor U8806 (N_8806,N_8743,N_8515);
nor U8807 (N_8807,N_8680,N_8666);
nor U8808 (N_8808,N_8652,N_8726);
or U8809 (N_8809,N_8687,N_8695);
or U8810 (N_8810,N_8575,N_8526);
nor U8811 (N_8811,N_8561,N_8548);
nand U8812 (N_8812,N_8655,N_8700);
nand U8813 (N_8813,N_8595,N_8681);
nor U8814 (N_8814,N_8712,N_8645);
nor U8815 (N_8815,N_8547,N_8525);
and U8816 (N_8816,N_8512,N_8739);
or U8817 (N_8817,N_8646,N_8662);
nand U8818 (N_8818,N_8593,N_8621);
or U8819 (N_8819,N_8554,N_8637);
nand U8820 (N_8820,N_8522,N_8594);
nor U8821 (N_8821,N_8717,N_8701);
nor U8822 (N_8822,N_8634,N_8625);
nor U8823 (N_8823,N_8542,N_8731);
nor U8824 (N_8824,N_8667,N_8694);
and U8825 (N_8825,N_8505,N_8576);
or U8826 (N_8826,N_8693,N_8714);
or U8827 (N_8827,N_8587,N_8620);
nor U8828 (N_8828,N_8676,N_8643);
and U8829 (N_8829,N_8533,N_8660);
nor U8830 (N_8830,N_8537,N_8624);
nand U8831 (N_8831,N_8619,N_8565);
nor U8832 (N_8832,N_8513,N_8749);
and U8833 (N_8833,N_8532,N_8531);
nor U8834 (N_8834,N_8635,N_8648);
or U8835 (N_8835,N_8670,N_8628);
and U8836 (N_8836,N_8558,N_8528);
and U8837 (N_8837,N_8626,N_8658);
nand U8838 (N_8838,N_8540,N_8672);
or U8839 (N_8839,N_8597,N_8578);
or U8840 (N_8840,N_8609,N_8629);
and U8841 (N_8841,N_8738,N_8517);
nor U8842 (N_8842,N_8633,N_8613);
nor U8843 (N_8843,N_8598,N_8596);
nor U8844 (N_8844,N_8709,N_8560);
or U8845 (N_8845,N_8733,N_8729);
nor U8846 (N_8846,N_8679,N_8557);
or U8847 (N_8847,N_8631,N_8684);
nand U8848 (N_8848,N_8555,N_8727);
or U8849 (N_8849,N_8683,N_8591);
or U8850 (N_8850,N_8553,N_8650);
or U8851 (N_8851,N_8586,N_8601);
and U8852 (N_8852,N_8616,N_8507);
and U8853 (N_8853,N_8608,N_8748);
nand U8854 (N_8854,N_8699,N_8736);
nand U8855 (N_8855,N_8582,N_8685);
or U8856 (N_8856,N_8724,N_8541);
or U8857 (N_8857,N_8630,N_8737);
nor U8858 (N_8858,N_8708,N_8610);
nor U8859 (N_8859,N_8585,N_8530);
or U8860 (N_8860,N_8661,N_8697);
or U8861 (N_8861,N_8612,N_8536);
nor U8862 (N_8862,N_8664,N_8663);
nand U8863 (N_8863,N_8707,N_8677);
nand U8864 (N_8864,N_8665,N_8640);
or U8865 (N_8865,N_8671,N_8705);
and U8866 (N_8866,N_8606,N_8552);
and U8867 (N_8867,N_8704,N_8675);
xnor U8868 (N_8868,N_8527,N_8580);
nor U8869 (N_8869,N_8544,N_8500);
nor U8870 (N_8870,N_8691,N_8577);
nor U8871 (N_8871,N_8589,N_8622);
and U8872 (N_8872,N_8710,N_8583);
nand U8873 (N_8873,N_8618,N_8615);
nand U8874 (N_8874,N_8520,N_8570);
or U8875 (N_8875,N_8507,N_8630);
nand U8876 (N_8876,N_8531,N_8668);
and U8877 (N_8877,N_8702,N_8647);
or U8878 (N_8878,N_8566,N_8698);
nand U8879 (N_8879,N_8627,N_8553);
or U8880 (N_8880,N_8747,N_8595);
and U8881 (N_8881,N_8521,N_8620);
or U8882 (N_8882,N_8689,N_8517);
nand U8883 (N_8883,N_8542,N_8588);
and U8884 (N_8884,N_8593,N_8571);
or U8885 (N_8885,N_8509,N_8603);
or U8886 (N_8886,N_8642,N_8685);
xor U8887 (N_8887,N_8727,N_8559);
nor U8888 (N_8888,N_8646,N_8700);
nor U8889 (N_8889,N_8524,N_8742);
nor U8890 (N_8890,N_8651,N_8697);
or U8891 (N_8891,N_8605,N_8515);
or U8892 (N_8892,N_8508,N_8524);
and U8893 (N_8893,N_8616,N_8606);
and U8894 (N_8894,N_8678,N_8716);
and U8895 (N_8895,N_8636,N_8743);
nor U8896 (N_8896,N_8553,N_8718);
nand U8897 (N_8897,N_8646,N_8554);
and U8898 (N_8898,N_8630,N_8616);
nor U8899 (N_8899,N_8535,N_8747);
xor U8900 (N_8900,N_8717,N_8676);
xnor U8901 (N_8901,N_8541,N_8651);
nand U8902 (N_8902,N_8617,N_8681);
nand U8903 (N_8903,N_8610,N_8613);
and U8904 (N_8904,N_8596,N_8581);
nor U8905 (N_8905,N_8567,N_8582);
and U8906 (N_8906,N_8587,N_8692);
or U8907 (N_8907,N_8668,N_8501);
xor U8908 (N_8908,N_8728,N_8515);
or U8909 (N_8909,N_8709,N_8671);
nand U8910 (N_8910,N_8665,N_8683);
nor U8911 (N_8911,N_8545,N_8660);
or U8912 (N_8912,N_8719,N_8710);
and U8913 (N_8913,N_8567,N_8602);
nand U8914 (N_8914,N_8604,N_8505);
nand U8915 (N_8915,N_8652,N_8629);
or U8916 (N_8916,N_8641,N_8556);
nand U8917 (N_8917,N_8679,N_8688);
xnor U8918 (N_8918,N_8701,N_8628);
and U8919 (N_8919,N_8507,N_8573);
nand U8920 (N_8920,N_8528,N_8579);
nor U8921 (N_8921,N_8568,N_8593);
nand U8922 (N_8922,N_8511,N_8695);
nand U8923 (N_8923,N_8744,N_8679);
nor U8924 (N_8924,N_8689,N_8608);
nand U8925 (N_8925,N_8706,N_8711);
or U8926 (N_8926,N_8567,N_8534);
nand U8927 (N_8927,N_8526,N_8572);
nor U8928 (N_8928,N_8514,N_8712);
nand U8929 (N_8929,N_8673,N_8602);
nor U8930 (N_8930,N_8523,N_8658);
xnor U8931 (N_8931,N_8681,N_8584);
nor U8932 (N_8932,N_8709,N_8602);
nand U8933 (N_8933,N_8529,N_8720);
nand U8934 (N_8934,N_8700,N_8639);
xnor U8935 (N_8935,N_8713,N_8685);
nor U8936 (N_8936,N_8557,N_8655);
nand U8937 (N_8937,N_8609,N_8627);
nand U8938 (N_8938,N_8565,N_8735);
or U8939 (N_8939,N_8679,N_8732);
or U8940 (N_8940,N_8740,N_8662);
and U8941 (N_8941,N_8615,N_8644);
nor U8942 (N_8942,N_8720,N_8528);
and U8943 (N_8943,N_8612,N_8511);
nand U8944 (N_8944,N_8702,N_8502);
or U8945 (N_8945,N_8563,N_8726);
nor U8946 (N_8946,N_8733,N_8687);
and U8947 (N_8947,N_8709,N_8611);
and U8948 (N_8948,N_8679,N_8657);
and U8949 (N_8949,N_8576,N_8639);
nor U8950 (N_8950,N_8509,N_8561);
nor U8951 (N_8951,N_8528,N_8545);
nor U8952 (N_8952,N_8698,N_8650);
or U8953 (N_8953,N_8595,N_8525);
and U8954 (N_8954,N_8641,N_8508);
nand U8955 (N_8955,N_8581,N_8561);
nand U8956 (N_8956,N_8589,N_8724);
or U8957 (N_8957,N_8559,N_8691);
and U8958 (N_8958,N_8632,N_8598);
and U8959 (N_8959,N_8522,N_8727);
nand U8960 (N_8960,N_8590,N_8706);
and U8961 (N_8961,N_8710,N_8506);
and U8962 (N_8962,N_8516,N_8693);
nor U8963 (N_8963,N_8678,N_8500);
or U8964 (N_8964,N_8582,N_8544);
xor U8965 (N_8965,N_8503,N_8646);
or U8966 (N_8966,N_8730,N_8690);
or U8967 (N_8967,N_8636,N_8689);
nor U8968 (N_8968,N_8716,N_8531);
or U8969 (N_8969,N_8504,N_8603);
nand U8970 (N_8970,N_8654,N_8710);
and U8971 (N_8971,N_8519,N_8707);
nand U8972 (N_8972,N_8525,N_8710);
or U8973 (N_8973,N_8561,N_8532);
and U8974 (N_8974,N_8558,N_8524);
and U8975 (N_8975,N_8603,N_8569);
and U8976 (N_8976,N_8579,N_8526);
and U8977 (N_8977,N_8737,N_8665);
and U8978 (N_8978,N_8661,N_8720);
nor U8979 (N_8979,N_8620,N_8596);
nor U8980 (N_8980,N_8632,N_8742);
nand U8981 (N_8981,N_8609,N_8733);
nor U8982 (N_8982,N_8518,N_8700);
and U8983 (N_8983,N_8697,N_8581);
and U8984 (N_8984,N_8508,N_8673);
nor U8985 (N_8985,N_8528,N_8511);
nand U8986 (N_8986,N_8696,N_8660);
and U8987 (N_8987,N_8747,N_8527);
and U8988 (N_8988,N_8509,N_8503);
nor U8989 (N_8989,N_8719,N_8706);
and U8990 (N_8990,N_8603,N_8697);
and U8991 (N_8991,N_8668,N_8584);
and U8992 (N_8992,N_8636,N_8596);
nand U8993 (N_8993,N_8701,N_8668);
nand U8994 (N_8994,N_8677,N_8674);
nor U8995 (N_8995,N_8604,N_8671);
nor U8996 (N_8996,N_8739,N_8656);
nand U8997 (N_8997,N_8708,N_8649);
nor U8998 (N_8998,N_8633,N_8511);
or U8999 (N_8999,N_8566,N_8680);
and U9000 (N_9000,N_8910,N_8760);
or U9001 (N_9001,N_8896,N_8868);
or U9002 (N_9002,N_8862,N_8898);
or U9003 (N_9003,N_8773,N_8883);
and U9004 (N_9004,N_8823,N_8916);
and U9005 (N_9005,N_8765,N_8884);
or U9006 (N_9006,N_8946,N_8864);
and U9007 (N_9007,N_8956,N_8912);
nand U9008 (N_9008,N_8997,N_8928);
or U9009 (N_9009,N_8787,N_8942);
nor U9010 (N_9010,N_8887,N_8797);
and U9011 (N_9011,N_8816,N_8799);
xor U9012 (N_9012,N_8899,N_8962);
nand U9013 (N_9013,N_8891,N_8959);
and U9014 (N_9014,N_8929,N_8813);
or U9015 (N_9015,N_8978,N_8781);
nand U9016 (N_9016,N_8763,N_8996);
nand U9017 (N_9017,N_8839,N_8963);
and U9018 (N_9018,N_8919,N_8828);
or U9019 (N_9019,N_8972,N_8885);
nor U9020 (N_9020,N_8917,N_8844);
nor U9021 (N_9021,N_8991,N_8779);
nor U9022 (N_9022,N_8834,N_8918);
and U9023 (N_9023,N_8922,N_8937);
nand U9024 (N_9024,N_8842,N_8855);
and U9025 (N_9025,N_8758,N_8971);
nand U9026 (N_9026,N_8854,N_8968);
nor U9027 (N_9027,N_8945,N_8788);
and U9028 (N_9028,N_8914,N_8821);
or U9029 (N_9029,N_8960,N_8908);
nor U9030 (N_9030,N_8833,N_8761);
or U9031 (N_9031,N_8984,N_8987);
nor U9032 (N_9032,N_8951,N_8785);
nor U9033 (N_9033,N_8811,N_8802);
nor U9034 (N_9034,N_8764,N_8766);
and U9035 (N_9035,N_8871,N_8931);
nand U9036 (N_9036,N_8870,N_8830);
nor U9037 (N_9037,N_8801,N_8909);
and U9038 (N_9038,N_8974,N_8815);
or U9039 (N_9039,N_8966,N_8882);
or U9040 (N_9040,N_8762,N_8933);
or U9041 (N_9041,N_8965,N_8940);
nand U9042 (N_9042,N_8867,N_8953);
nor U9043 (N_9043,N_8961,N_8893);
or U9044 (N_9044,N_8944,N_8925);
nand U9045 (N_9045,N_8999,N_8983);
nand U9046 (N_9046,N_8806,N_8750);
and U9047 (N_9047,N_8789,N_8778);
xnor U9048 (N_9048,N_8767,N_8905);
nand U9049 (N_9049,N_8881,N_8992);
nand U9050 (N_9050,N_8783,N_8792);
nand U9051 (N_9051,N_8793,N_8849);
and U9052 (N_9052,N_8993,N_8814);
or U9053 (N_9053,N_8865,N_8994);
nor U9054 (N_9054,N_8784,N_8822);
or U9055 (N_9055,N_8847,N_8936);
or U9056 (N_9056,N_8782,N_8795);
and U9057 (N_9057,N_8930,N_8901);
nand U9058 (N_9058,N_8810,N_8895);
or U9059 (N_9059,N_8866,N_8955);
or U9060 (N_9060,N_8958,N_8818);
and U9061 (N_9061,N_8973,N_8804);
or U9062 (N_9062,N_8894,N_8857);
nand U9063 (N_9063,N_8923,N_8976);
or U9064 (N_9064,N_8776,N_8886);
and U9065 (N_9065,N_8935,N_8875);
nor U9066 (N_9066,N_8863,N_8879);
or U9067 (N_9067,N_8751,N_8780);
or U9068 (N_9068,N_8981,N_8954);
and U9069 (N_9069,N_8990,N_8812);
or U9070 (N_9070,N_8790,N_8995);
nand U9071 (N_9071,N_8920,N_8775);
nand U9072 (N_9072,N_8820,N_8851);
or U9073 (N_9073,N_8756,N_8924);
nand U9074 (N_9074,N_8943,N_8846);
and U9075 (N_9075,N_8998,N_8808);
nand U9076 (N_9076,N_8800,N_8938);
and U9077 (N_9077,N_8948,N_8827);
nor U9078 (N_9078,N_8835,N_8859);
nand U9079 (N_9079,N_8969,N_8807);
or U9080 (N_9080,N_8869,N_8975);
nand U9081 (N_9081,N_8902,N_8932);
nor U9082 (N_9082,N_8843,N_8982);
and U9083 (N_9083,N_8786,N_8888);
nor U9084 (N_9084,N_8877,N_8826);
nor U9085 (N_9085,N_8825,N_8829);
and U9086 (N_9086,N_8915,N_8988);
and U9087 (N_9087,N_8805,N_8853);
and U9088 (N_9088,N_8831,N_8913);
xor U9089 (N_9089,N_8757,N_8770);
nor U9090 (N_9090,N_8980,N_8900);
or U9091 (N_9091,N_8819,N_8809);
or U9092 (N_9092,N_8777,N_8840);
nand U9093 (N_9093,N_8874,N_8967);
nor U9094 (N_9094,N_8759,N_8771);
nor U9095 (N_9095,N_8986,N_8768);
nor U9096 (N_9096,N_8832,N_8845);
nand U9097 (N_9097,N_8752,N_8911);
nor U9098 (N_9098,N_8860,N_8824);
nand U9099 (N_9099,N_8796,N_8964);
or U9100 (N_9100,N_8878,N_8861);
or U9101 (N_9101,N_8939,N_8949);
nor U9102 (N_9102,N_8841,N_8798);
xor U9103 (N_9103,N_8957,N_8794);
nand U9104 (N_9104,N_8837,N_8889);
nor U9105 (N_9105,N_8872,N_8904);
and U9106 (N_9106,N_8817,N_8906);
nand U9107 (N_9107,N_8897,N_8979);
or U9108 (N_9108,N_8836,N_8970);
nand U9109 (N_9109,N_8873,N_8890);
nor U9110 (N_9110,N_8907,N_8952);
nor U9111 (N_9111,N_8754,N_8941);
and U9112 (N_9112,N_8927,N_8838);
nand U9113 (N_9113,N_8892,N_8753);
nor U9114 (N_9114,N_8880,N_8858);
or U9115 (N_9115,N_8755,N_8989);
or U9116 (N_9116,N_8926,N_8791);
nor U9117 (N_9117,N_8769,N_8856);
nor U9118 (N_9118,N_8848,N_8774);
or U9119 (N_9119,N_8903,N_8772);
nand U9120 (N_9120,N_8985,N_8977);
nand U9121 (N_9121,N_8852,N_8947);
nor U9122 (N_9122,N_8850,N_8921);
or U9123 (N_9123,N_8950,N_8934);
nand U9124 (N_9124,N_8876,N_8803);
and U9125 (N_9125,N_8846,N_8897);
nor U9126 (N_9126,N_8942,N_8932);
nand U9127 (N_9127,N_8781,N_8835);
or U9128 (N_9128,N_8995,N_8826);
nor U9129 (N_9129,N_8983,N_8769);
nor U9130 (N_9130,N_8880,N_8781);
xnor U9131 (N_9131,N_8860,N_8779);
xnor U9132 (N_9132,N_8854,N_8888);
nand U9133 (N_9133,N_8826,N_8803);
and U9134 (N_9134,N_8756,N_8951);
nand U9135 (N_9135,N_8863,N_8775);
xor U9136 (N_9136,N_8798,N_8924);
nand U9137 (N_9137,N_8841,N_8994);
and U9138 (N_9138,N_8803,N_8874);
nand U9139 (N_9139,N_8973,N_8801);
and U9140 (N_9140,N_8876,N_8895);
nand U9141 (N_9141,N_8967,N_8770);
nand U9142 (N_9142,N_8950,N_8872);
nor U9143 (N_9143,N_8820,N_8985);
nor U9144 (N_9144,N_8837,N_8828);
nor U9145 (N_9145,N_8945,N_8896);
nand U9146 (N_9146,N_8814,N_8824);
nor U9147 (N_9147,N_8825,N_8754);
and U9148 (N_9148,N_8929,N_8752);
and U9149 (N_9149,N_8755,N_8954);
and U9150 (N_9150,N_8993,N_8899);
nor U9151 (N_9151,N_8751,N_8774);
or U9152 (N_9152,N_8825,N_8962);
and U9153 (N_9153,N_8946,N_8768);
xnor U9154 (N_9154,N_8961,N_8794);
nand U9155 (N_9155,N_8928,N_8937);
nand U9156 (N_9156,N_8971,N_8970);
nor U9157 (N_9157,N_8818,N_8997);
and U9158 (N_9158,N_8922,N_8790);
or U9159 (N_9159,N_8761,N_8802);
nor U9160 (N_9160,N_8908,N_8936);
or U9161 (N_9161,N_8956,N_8754);
nor U9162 (N_9162,N_8772,N_8796);
xnor U9163 (N_9163,N_8853,N_8894);
nor U9164 (N_9164,N_8775,N_8939);
or U9165 (N_9165,N_8938,N_8849);
and U9166 (N_9166,N_8794,N_8778);
or U9167 (N_9167,N_8818,N_8946);
nand U9168 (N_9168,N_8874,N_8852);
nand U9169 (N_9169,N_8955,N_8995);
and U9170 (N_9170,N_8849,N_8988);
xor U9171 (N_9171,N_8816,N_8853);
xnor U9172 (N_9172,N_8813,N_8817);
or U9173 (N_9173,N_8975,N_8991);
nand U9174 (N_9174,N_8766,N_8867);
and U9175 (N_9175,N_8921,N_8959);
and U9176 (N_9176,N_8816,N_8761);
nor U9177 (N_9177,N_8781,N_8810);
xnor U9178 (N_9178,N_8974,N_8820);
nor U9179 (N_9179,N_8985,N_8840);
nor U9180 (N_9180,N_8750,N_8903);
or U9181 (N_9181,N_8817,N_8945);
or U9182 (N_9182,N_8954,N_8994);
and U9183 (N_9183,N_8758,N_8839);
nor U9184 (N_9184,N_8900,N_8899);
nand U9185 (N_9185,N_8774,N_8801);
nor U9186 (N_9186,N_8869,N_8874);
and U9187 (N_9187,N_8986,N_8895);
nand U9188 (N_9188,N_8877,N_8869);
or U9189 (N_9189,N_8960,N_8807);
nand U9190 (N_9190,N_8852,N_8924);
nor U9191 (N_9191,N_8944,N_8803);
nor U9192 (N_9192,N_8940,N_8902);
nand U9193 (N_9193,N_8785,N_8868);
and U9194 (N_9194,N_8817,N_8867);
or U9195 (N_9195,N_8842,N_8776);
or U9196 (N_9196,N_8939,N_8936);
and U9197 (N_9197,N_8819,N_8875);
nor U9198 (N_9198,N_8829,N_8951);
or U9199 (N_9199,N_8971,N_8868);
or U9200 (N_9200,N_8924,N_8755);
or U9201 (N_9201,N_8799,N_8878);
nand U9202 (N_9202,N_8937,N_8867);
and U9203 (N_9203,N_8825,N_8968);
or U9204 (N_9204,N_8969,N_8895);
and U9205 (N_9205,N_8988,N_8775);
nand U9206 (N_9206,N_8803,N_8930);
nor U9207 (N_9207,N_8890,N_8971);
nand U9208 (N_9208,N_8787,N_8957);
and U9209 (N_9209,N_8759,N_8765);
nor U9210 (N_9210,N_8954,N_8851);
nand U9211 (N_9211,N_8964,N_8852);
nand U9212 (N_9212,N_8788,N_8770);
or U9213 (N_9213,N_8768,N_8795);
nor U9214 (N_9214,N_8856,N_8827);
nand U9215 (N_9215,N_8916,N_8953);
nor U9216 (N_9216,N_8815,N_8753);
nand U9217 (N_9217,N_8848,N_8987);
or U9218 (N_9218,N_8951,N_8753);
nor U9219 (N_9219,N_8965,N_8962);
nand U9220 (N_9220,N_8832,N_8755);
nand U9221 (N_9221,N_8759,N_8919);
and U9222 (N_9222,N_8938,N_8992);
nor U9223 (N_9223,N_8977,N_8842);
nand U9224 (N_9224,N_8850,N_8933);
or U9225 (N_9225,N_8909,N_8857);
and U9226 (N_9226,N_8991,N_8828);
nand U9227 (N_9227,N_8789,N_8802);
or U9228 (N_9228,N_8835,N_8776);
nand U9229 (N_9229,N_8996,N_8812);
or U9230 (N_9230,N_8986,N_8796);
nand U9231 (N_9231,N_8897,N_8935);
nor U9232 (N_9232,N_8913,N_8918);
nand U9233 (N_9233,N_8777,N_8941);
or U9234 (N_9234,N_8883,N_8795);
or U9235 (N_9235,N_8988,N_8772);
or U9236 (N_9236,N_8929,N_8920);
or U9237 (N_9237,N_8800,N_8989);
nand U9238 (N_9238,N_8968,N_8945);
and U9239 (N_9239,N_8776,N_8874);
and U9240 (N_9240,N_8840,N_8889);
and U9241 (N_9241,N_8989,N_8917);
nor U9242 (N_9242,N_8996,N_8785);
or U9243 (N_9243,N_8900,N_8926);
or U9244 (N_9244,N_8774,N_8830);
nand U9245 (N_9245,N_8880,N_8925);
and U9246 (N_9246,N_8757,N_8917);
or U9247 (N_9247,N_8850,N_8826);
nor U9248 (N_9248,N_8916,N_8899);
or U9249 (N_9249,N_8961,N_8999);
nand U9250 (N_9250,N_9101,N_9010);
nand U9251 (N_9251,N_9168,N_9206);
or U9252 (N_9252,N_9005,N_9194);
and U9253 (N_9253,N_9034,N_9241);
nor U9254 (N_9254,N_9240,N_9120);
or U9255 (N_9255,N_9067,N_9243);
nor U9256 (N_9256,N_9116,N_9160);
and U9257 (N_9257,N_9114,N_9149);
nor U9258 (N_9258,N_9176,N_9202);
and U9259 (N_9259,N_9150,N_9073);
nor U9260 (N_9260,N_9175,N_9169);
nand U9261 (N_9261,N_9204,N_9135);
nand U9262 (N_9262,N_9105,N_9213);
and U9263 (N_9263,N_9155,N_9110);
nor U9264 (N_9264,N_9062,N_9173);
and U9265 (N_9265,N_9195,N_9170);
xnor U9266 (N_9266,N_9183,N_9045);
nor U9267 (N_9267,N_9222,N_9069);
nand U9268 (N_9268,N_9108,N_9248);
nor U9269 (N_9269,N_9234,N_9154);
nand U9270 (N_9270,N_9184,N_9066);
nand U9271 (N_9271,N_9079,N_9163);
and U9272 (N_9272,N_9187,N_9230);
and U9273 (N_9273,N_9221,N_9166);
nor U9274 (N_9274,N_9082,N_9092);
nand U9275 (N_9275,N_9012,N_9139);
nand U9276 (N_9276,N_9188,N_9218);
and U9277 (N_9277,N_9239,N_9203);
or U9278 (N_9278,N_9174,N_9233);
nand U9279 (N_9279,N_9137,N_9227);
nor U9280 (N_9280,N_9245,N_9162);
or U9281 (N_9281,N_9159,N_9231);
nor U9282 (N_9282,N_9236,N_9180);
or U9283 (N_9283,N_9044,N_9128);
nor U9284 (N_9284,N_9216,N_9070);
nand U9285 (N_9285,N_9145,N_9060);
and U9286 (N_9286,N_9164,N_9232);
nand U9287 (N_9287,N_9247,N_9104);
nand U9288 (N_9288,N_9096,N_9225);
and U9289 (N_9289,N_9043,N_9026);
or U9290 (N_9290,N_9085,N_9119);
or U9291 (N_9291,N_9052,N_9091);
nor U9292 (N_9292,N_9007,N_9153);
nand U9293 (N_9293,N_9013,N_9205);
nor U9294 (N_9294,N_9083,N_9215);
xor U9295 (N_9295,N_9140,N_9030);
nand U9296 (N_9296,N_9078,N_9144);
nand U9297 (N_9297,N_9212,N_9017);
nor U9298 (N_9298,N_9132,N_9041);
or U9299 (N_9299,N_9022,N_9001);
and U9300 (N_9300,N_9152,N_9037);
nor U9301 (N_9301,N_9249,N_9165);
nor U9302 (N_9302,N_9217,N_9197);
or U9303 (N_9303,N_9011,N_9042);
or U9304 (N_9304,N_9098,N_9029);
or U9305 (N_9305,N_9242,N_9109);
nand U9306 (N_9306,N_9229,N_9058);
xnor U9307 (N_9307,N_9046,N_9051);
and U9308 (N_9308,N_9002,N_9000);
nand U9309 (N_9309,N_9077,N_9090);
nand U9310 (N_9310,N_9141,N_9064);
and U9311 (N_9311,N_9056,N_9006);
nor U9312 (N_9312,N_9027,N_9228);
or U9313 (N_9313,N_9093,N_9148);
xnor U9314 (N_9314,N_9238,N_9196);
nand U9315 (N_9315,N_9038,N_9146);
nor U9316 (N_9316,N_9123,N_9057);
nand U9317 (N_9317,N_9033,N_9072);
nand U9318 (N_9318,N_9099,N_9192);
and U9319 (N_9319,N_9050,N_9179);
nor U9320 (N_9320,N_9126,N_9118);
and U9321 (N_9321,N_9015,N_9156);
nand U9322 (N_9322,N_9124,N_9003);
nor U9323 (N_9323,N_9074,N_9127);
or U9324 (N_9324,N_9063,N_9084);
or U9325 (N_9325,N_9136,N_9246);
nand U9326 (N_9326,N_9220,N_9113);
or U9327 (N_9327,N_9054,N_9181);
nor U9328 (N_9328,N_9095,N_9039);
or U9329 (N_9329,N_9122,N_9237);
nor U9330 (N_9330,N_9081,N_9224);
and U9331 (N_9331,N_9147,N_9178);
nor U9332 (N_9332,N_9076,N_9055);
and U9333 (N_9333,N_9199,N_9040);
and U9334 (N_9334,N_9191,N_9068);
and U9335 (N_9335,N_9177,N_9244);
or U9336 (N_9336,N_9129,N_9036);
or U9337 (N_9337,N_9172,N_9219);
and U9338 (N_9338,N_9214,N_9061);
and U9339 (N_9339,N_9087,N_9089);
nor U9340 (N_9340,N_9185,N_9049);
nand U9341 (N_9341,N_9024,N_9209);
and U9342 (N_9342,N_9161,N_9125);
nand U9343 (N_9343,N_9200,N_9071);
nand U9344 (N_9344,N_9053,N_9065);
and U9345 (N_9345,N_9107,N_9182);
nand U9346 (N_9346,N_9142,N_9020);
nor U9347 (N_9347,N_9115,N_9138);
and U9348 (N_9348,N_9131,N_9097);
xor U9349 (N_9349,N_9094,N_9028);
or U9350 (N_9350,N_9023,N_9117);
or U9351 (N_9351,N_9198,N_9167);
or U9352 (N_9352,N_9130,N_9151);
and U9353 (N_9353,N_9193,N_9019);
xor U9354 (N_9354,N_9025,N_9088);
and U9355 (N_9355,N_9208,N_9059);
nand U9356 (N_9356,N_9133,N_9106);
nor U9357 (N_9357,N_9080,N_9235);
or U9358 (N_9358,N_9004,N_9035);
and U9359 (N_9359,N_9016,N_9211);
or U9360 (N_9360,N_9103,N_9223);
nand U9361 (N_9361,N_9226,N_9201);
or U9362 (N_9362,N_9100,N_9134);
nand U9363 (N_9363,N_9009,N_9111);
and U9364 (N_9364,N_9190,N_9048);
nand U9365 (N_9365,N_9157,N_9210);
nand U9366 (N_9366,N_9086,N_9102);
nor U9367 (N_9367,N_9121,N_9032);
xor U9368 (N_9368,N_9018,N_9014);
or U9369 (N_9369,N_9031,N_9158);
nor U9370 (N_9370,N_9207,N_9075);
and U9371 (N_9371,N_9047,N_9143);
nor U9372 (N_9372,N_9171,N_9189);
nor U9373 (N_9373,N_9186,N_9021);
nor U9374 (N_9374,N_9008,N_9112);
and U9375 (N_9375,N_9158,N_9054);
nand U9376 (N_9376,N_9119,N_9139);
nand U9377 (N_9377,N_9126,N_9124);
nor U9378 (N_9378,N_9047,N_9029);
or U9379 (N_9379,N_9215,N_9230);
nor U9380 (N_9380,N_9079,N_9157);
or U9381 (N_9381,N_9204,N_9065);
and U9382 (N_9382,N_9153,N_9230);
or U9383 (N_9383,N_9119,N_9244);
and U9384 (N_9384,N_9206,N_9014);
nor U9385 (N_9385,N_9154,N_9102);
or U9386 (N_9386,N_9126,N_9216);
or U9387 (N_9387,N_9150,N_9197);
or U9388 (N_9388,N_9079,N_9020);
and U9389 (N_9389,N_9164,N_9073);
and U9390 (N_9390,N_9070,N_9045);
or U9391 (N_9391,N_9044,N_9145);
nand U9392 (N_9392,N_9159,N_9021);
nor U9393 (N_9393,N_9061,N_9100);
nor U9394 (N_9394,N_9082,N_9036);
nor U9395 (N_9395,N_9095,N_9160);
and U9396 (N_9396,N_9077,N_9017);
and U9397 (N_9397,N_9175,N_9071);
and U9398 (N_9398,N_9213,N_9079);
nor U9399 (N_9399,N_9015,N_9204);
and U9400 (N_9400,N_9071,N_9172);
or U9401 (N_9401,N_9209,N_9039);
nand U9402 (N_9402,N_9051,N_9207);
nor U9403 (N_9403,N_9076,N_9231);
and U9404 (N_9404,N_9217,N_9060);
nand U9405 (N_9405,N_9031,N_9057);
and U9406 (N_9406,N_9187,N_9155);
and U9407 (N_9407,N_9192,N_9011);
nor U9408 (N_9408,N_9061,N_9086);
and U9409 (N_9409,N_9061,N_9231);
nor U9410 (N_9410,N_9218,N_9140);
xnor U9411 (N_9411,N_9085,N_9054);
or U9412 (N_9412,N_9017,N_9011);
nand U9413 (N_9413,N_9063,N_9152);
and U9414 (N_9414,N_9201,N_9063);
or U9415 (N_9415,N_9087,N_9102);
or U9416 (N_9416,N_9069,N_9231);
xor U9417 (N_9417,N_9182,N_9216);
and U9418 (N_9418,N_9146,N_9149);
nand U9419 (N_9419,N_9162,N_9148);
and U9420 (N_9420,N_9003,N_9248);
nand U9421 (N_9421,N_9033,N_9016);
or U9422 (N_9422,N_9192,N_9002);
nand U9423 (N_9423,N_9227,N_9239);
nand U9424 (N_9424,N_9162,N_9128);
and U9425 (N_9425,N_9152,N_9161);
nor U9426 (N_9426,N_9062,N_9004);
or U9427 (N_9427,N_9119,N_9015);
nand U9428 (N_9428,N_9022,N_9063);
nor U9429 (N_9429,N_9248,N_9062);
nand U9430 (N_9430,N_9094,N_9106);
and U9431 (N_9431,N_9181,N_9018);
and U9432 (N_9432,N_9161,N_9084);
nand U9433 (N_9433,N_9100,N_9034);
nor U9434 (N_9434,N_9181,N_9028);
nand U9435 (N_9435,N_9018,N_9110);
or U9436 (N_9436,N_9113,N_9163);
or U9437 (N_9437,N_9051,N_9087);
or U9438 (N_9438,N_9059,N_9152);
nand U9439 (N_9439,N_9187,N_9072);
nand U9440 (N_9440,N_9019,N_9239);
and U9441 (N_9441,N_9204,N_9187);
or U9442 (N_9442,N_9022,N_9240);
nor U9443 (N_9443,N_9211,N_9062);
or U9444 (N_9444,N_9067,N_9173);
or U9445 (N_9445,N_9121,N_9219);
and U9446 (N_9446,N_9171,N_9077);
or U9447 (N_9447,N_9142,N_9201);
and U9448 (N_9448,N_9249,N_9163);
nand U9449 (N_9449,N_9080,N_9096);
and U9450 (N_9450,N_9057,N_9003);
nand U9451 (N_9451,N_9063,N_9216);
nand U9452 (N_9452,N_9095,N_9056);
or U9453 (N_9453,N_9030,N_9010);
nand U9454 (N_9454,N_9009,N_9013);
nor U9455 (N_9455,N_9225,N_9114);
and U9456 (N_9456,N_9238,N_9113);
nand U9457 (N_9457,N_9020,N_9037);
and U9458 (N_9458,N_9019,N_9203);
nand U9459 (N_9459,N_9227,N_9218);
nor U9460 (N_9460,N_9019,N_9176);
nor U9461 (N_9461,N_9148,N_9183);
nor U9462 (N_9462,N_9182,N_9170);
nand U9463 (N_9463,N_9190,N_9176);
nand U9464 (N_9464,N_9097,N_9185);
nand U9465 (N_9465,N_9216,N_9139);
and U9466 (N_9466,N_9219,N_9139);
and U9467 (N_9467,N_9067,N_9155);
nor U9468 (N_9468,N_9135,N_9227);
or U9469 (N_9469,N_9201,N_9153);
nand U9470 (N_9470,N_9123,N_9073);
and U9471 (N_9471,N_9211,N_9146);
xor U9472 (N_9472,N_9216,N_9101);
nor U9473 (N_9473,N_9153,N_9078);
or U9474 (N_9474,N_9026,N_9094);
nand U9475 (N_9475,N_9056,N_9154);
and U9476 (N_9476,N_9113,N_9013);
nor U9477 (N_9477,N_9050,N_9002);
or U9478 (N_9478,N_9188,N_9061);
nor U9479 (N_9479,N_9108,N_9006);
or U9480 (N_9480,N_9196,N_9173);
nor U9481 (N_9481,N_9118,N_9208);
or U9482 (N_9482,N_9217,N_9184);
and U9483 (N_9483,N_9149,N_9110);
nor U9484 (N_9484,N_9243,N_9047);
nor U9485 (N_9485,N_9063,N_9093);
nor U9486 (N_9486,N_9170,N_9053);
and U9487 (N_9487,N_9111,N_9161);
nor U9488 (N_9488,N_9107,N_9110);
nor U9489 (N_9489,N_9201,N_9044);
or U9490 (N_9490,N_9178,N_9143);
nand U9491 (N_9491,N_9245,N_9057);
and U9492 (N_9492,N_9141,N_9162);
nor U9493 (N_9493,N_9105,N_9203);
nor U9494 (N_9494,N_9125,N_9074);
nor U9495 (N_9495,N_9089,N_9085);
and U9496 (N_9496,N_9050,N_9109);
or U9497 (N_9497,N_9099,N_9069);
nor U9498 (N_9498,N_9073,N_9196);
and U9499 (N_9499,N_9102,N_9221);
or U9500 (N_9500,N_9407,N_9327);
nand U9501 (N_9501,N_9374,N_9284);
and U9502 (N_9502,N_9443,N_9316);
nor U9503 (N_9503,N_9317,N_9393);
or U9504 (N_9504,N_9437,N_9252);
nor U9505 (N_9505,N_9481,N_9396);
and U9506 (N_9506,N_9345,N_9277);
nor U9507 (N_9507,N_9323,N_9294);
nand U9508 (N_9508,N_9320,N_9324);
or U9509 (N_9509,N_9429,N_9455);
nand U9510 (N_9510,N_9351,N_9414);
or U9511 (N_9511,N_9258,N_9273);
and U9512 (N_9512,N_9452,N_9298);
nand U9513 (N_9513,N_9279,N_9336);
nand U9514 (N_9514,N_9420,N_9494);
and U9515 (N_9515,N_9391,N_9373);
nor U9516 (N_9516,N_9435,N_9255);
and U9517 (N_9517,N_9495,N_9472);
nor U9518 (N_9518,N_9377,N_9422);
or U9519 (N_9519,N_9359,N_9459);
nand U9520 (N_9520,N_9405,N_9441);
nand U9521 (N_9521,N_9306,N_9498);
nor U9522 (N_9522,N_9309,N_9426);
or U9523 (N_9523,N_9382,N_9385);
or U9524 (N_9524,N_9264,N_9434);
or U9525 (N_9525,N_9253,N_9484);
nor U9526 (N_9526,N_9444,N_9406);
and U9527 (N_9527,N_9398,N_9321);
nor U9528 (N_9528,N_9283,N_9346);
and U9529 (N_9529,N_9412,N_9492);
nor U9530 (N_9530,N_9463,N_9311);
nor U9531 (N_9531,N_9278,N_9402);
or U9532 (N_9532,N_9383,N_9421);
nor U9533 (N_9533,N_9487,N_9315);
and U9534 (N_9534,N_9378,N_9295);
and U9535 (N_9535,N_9286,N_9318);
nand U9536 (N_9536,N_9260,N_9267);
or U9537 (N_9537,N_9301,N_9423);
or U9538 (N_9538,N_9416,N_9310);
nand U9539 (N_9539,N_9394,N_9454);
or U9540 (N_9540,N_9296,N_9413);
nor U9541 (N_9541,N_9325,N_9489);
xor U9542 (N_9542,N_9409,N_9331);
nor U9543 (N_9543,N_9375,N_9352);
and U9544 (N_9544,N_9457,N_9330);
or U9545 (N_9545,N_9342,N_9458);
or U9546 (N_9546,N_9427,N_9361);
nor U9547 (N_9547,N_9466,N_9370);
or U9548 (N_9548,N_9282,N_9265);
nor U9549 (N_9549,N_9372,N_9337);
nand U9550 (N_9550,N_9461,N_9460);
and U9551 (N_9551,N_9381,N_9271);
and U9552 (N_9552,N_9432,N_9251);
nand U9553 (N_9553,N_9367,N_9379);
nand U9554 (N_9554,N_9476,N_9479);
and U9555 (N_9555,N_9482,N_9450);
or U9556 (N_9556,N_9308,N_9281);
nand U9557 (N_9557,N_9371,N_9266);
and U9558 (N_9558,N_9274,N_9387);
or U9559 (N_9559,N_9328,N_9467);
and U9560 (N_9560,N_9433,N_9490);
nor U9561 (N_9561,N_9456,N_9488);
or U9562 (N_9562,N_9369,N_9362);
nand U9563 (N_9563,N_9341,N_9288);
nor U9564 (N_9564,N_9477,N_9497);
nor U9565 (N_9565,N_9365,N_9384);
nor U9566 (N_9566,N_9438,N_9289);
nand U9567 (N_9567,N_9478,N_9430);
nor U9568 (N_9568,N_9386,N_9493);
and U9569 (N_9569,N_9410,N_9499);
nand U9570 (N_9570,N_9335,N_9471);
nor U9571 (N_9571,N_9340,N_9483);
and U9572 (N_9572,N_9439,N_9305);
or U9573 (N_9573,N_9350,N_9275);
and U9574 (N_9574,N_9401,N_9332);
nor U9575 (N_9575,N_9411,N_9300);
nand U9576 (N_9576,N_9338,N_9297);
or U9577 (N_9577,N_9408,N_9333);
nor U9578 (N_9578,N_9280,N_9449);
nor U9579 (N_9579,N_9276,N_9363);
nor U9580 (N_9580,N_9451,N_9388);
and U9581 (N_9581,N_9339,N_9272);
and U9582 (N_9582,N_9496,N_9263);
nand U9583 (N_9583,N_9262,N_9254);
or U9584 (N_9584,N_9355,N_9259);
nand U9585 (N_9585,N_9389,N_9436);
nor U9586 (N_9586,N_9291,N_9285);
and U9587 (N_9587,N_9428,N_9474);
or U9588 (N_9588,N_9314,N_9480);
and U9589 (N_9589,N_9293,N_9329);
nor U9590 (N_9590,N_9465,N_9442);
nand U9591 (N_9591,N_9485,N_9304);
nand U9592 (N_9592,N_9425,N_9364);
and U9593 (N_9593,N_9343,N_9415);
xor U9594 (N_9594,N_9307,N_9319);
or U9595 (N_9595,N_9403,N_9270);
xnor U9596 (N_9596,N_9464,N_9395);
and U9597 (N_9597,N_9475,N_9360);
nor U9598 (N_9598,N_9334,N_9349);
and U9599 (N_9599,N_9462,N_9431);
nand U9600 (N_9600,N_9400,N_9473);
nand U9601 (N_9601,N_9322,N_9268);
nor U9602 (N_9602,N_9353,N_9256);
nor U9603 (N_9603,N_9261,N_9368);
or U9604 (N_9604,N_9348,N_9446);
and U9605 (N_9605,N_9404,N_9269);
nor U9606 (N_9606,N_9470,N_9445);
or U9607 (N_9607,N_9417,N_9326);
or U9608 (N_9608,N_9399,N_9486);
nand U9609 (N_9609,N_9380,N_9290);
nor U9610 (N_9610,N_9312,N_9447);
xnor U9611 (N_9611,N_9250,N_9354);
nand U9612 (N_9612,N_9344,N_9376);
nand U9613 (N_9613,N_9468,N_9419);
nor U9614 (N_9614,N_9448,N_9299);
nand U9615 (N_9615,N_9397,N_9347);
nor U9616 (N_9616,N_9453,N_9292);
and U9617 (N_9617,N_9424,N_9303);
or U9618 (N_9618,N_9366,N_9392);
or U9619 (N_9619,N_9302,N_9418);
nand U9620 (N_9620,N_9358,N_9440);
and U9621 (N_9621,N_9469,N_9357);
nand U9622 (N_9622,N_9313,N_9356);
nor U9623 (N_9623,N_9257,N_9491);
nand U9624 (N_9624,N_9287,N_9390);
nor U9625 (N_9625,N_9358,N_9256);
and U9626 (N_9626,N_9290,N_9444);
and U9627 (N_9627,N_9403,N_9320);
and U9628 (N_9628,N_9318,N_9336);
or U9629 (N_9629,N_9434,N_9322);
or U9630 (N_9630,N_9450,N_9435);
nand U9631 (N_9631,N_9259,N_9414);
nand U9632 (N_9632,N_9381,N_9374);
and U9633 (N_9633,N_9448,N_9441);
or U9634 (N_9634,N_9354,N_9302);
nand U9635 (N_9635,N_9336,N_9352);
or U9636 (N_9636,N_9423,N_9436);
nor U9637 (N_9637,N_9312,N_9388);
and U9638 (N_9638,N_9291,N_9404);
and U9639 (N_9639,N_9390,N_9292);
nand U9640 (N_9640,N_9318,N_9472);
nor U9641 (N_9641,N_9467,N_9390);
nor U9642 (N_9642,N_9446,N_9289);
or U9643 (N_9643,N_9276,N_9329);
nor U9644 (N_9644,N_9409,N_9259);
or U9645 (N_9645,N_9495,N_9499);
nand U9646 (N_9646,N_9330,N_9375);
or U9647 (N_9647,N_9478,N_9399);
and U9648 (N_9648,N_9400,N_9258);
or U9649 (N_9649,N_9268,N_9252);
or U9650 (N_9650,N_9413,N_9470);
and U9651 (N_9651,N_9321,N_9311);
nand U9652 (N_9652,N_9475,N_9362);
nor U9653 (N_9653,N_9463,N_9308);
nor U9654 (N_9654,N_9406,N_9437);
and U9655 (N_9655,N_9406,N_9299);
or U9656 (N_9656,N_9453,N_9441);
nand U9657 (N_9657,N_9331,N_9455);
and U9658 (N_9658,N_9364,N_9453);
or U9659 (N_9659,N_9301,N_9325);
nand U9660 (N_9660,N_9437,N_9392);
and U9661 (N_9661,N_9333,N_9309);
and U9662 (N_9662,N_9291,N_9480);
and U9663 (N_9663,N_9252,N_9426);
or U9664 (N_9664,N_9396,N_9303);
nor U9665 (N_9665,N_9490,N_9270);
nand U9666 (N_9666,N_9413,N_9272);
nor U9667 (N_9667,N_9485,N_9411);
nand U9668 (N_9668,N_9387,N_9452);
or U9669 (N_9669,N_9376,N_9369);
nand U9670 (N_9670,N_9363,N_9345);
or U9671 (N_9671,N_9264,N_9383);
xor U9672 (N_9672,N_9270,N_9360);
nand U9673 (N_9673,N_9476,N_9297);
nor U9674 (N_9674,N_9374,N_9373);
or U9675 (N_9675,N_9408,N_9445);
or U9676 (N_9676,N_9328,N_9452);
and U9677 (N_9677,N_9498,N_9463);
or U9678 (N_9678,N_9477,N_9298);
xor U9679 (N_9679,N_9450,N_9365);
or U9680 (N_9680,N_9348,N_9341);
nor U9681 (N_9681,N_9331,N_9373);
and U9682 (N_9682,N_9435,N_9260);
and U9683 (N_9683,N_9462,N_9334);
nor U9684 (N_9684,N_9456,N_9470);
nand U9685 (N_9685,N_9302,N_9355);
or U9686 (N_9686,N_9366,N_9496);
nand U9687 (N_9687,N_9272,N_9286);
xnor U9688 (N_9688,N_9372,N_9475);
nor U9689 (N_9689,N_9355,N_9470);
and U9690 (N_9690,N_9355,N_9337);
nand U9691 (N_9691,N_9336,N_9303);
and U9692 (N_9692,N_9382,N_9273);
and U9693 (N_9693,N_9301,N_9315);
or U9694 (N_9694,N_9357,N_9482);
and U9695 (N_9695,N_9320,N_9441);
nor U9696 (N_9696,N_9363,N_9337);
nor U9697 (N_9697,N_9274,N_9453);
nand U9698 (N_9698,N_9487,N_9428);
nor U9699 (N_9699,N_9364,N_9319);
nand U9700 (N_9700,N_9369,N_9439);
nor U9701 (N_9701,N_9360,N_9332);
nand U9702 (N_9702,N_9337,N_9299);
nand U9703 (N_9703,N_9428,N_9429);
nand U9704 (N_9704,N_9334,N_9481);
or U9705 (N_9705,N_9441,N_9420);
nor U9706 (N_9706,N_9414,N_9427);
or U9707 (N_9707,N_9260,N_9496);
nor U9708 (N_9708,N_9258,N_9283);
nor U9709 (N_9709,N_9386,N_9408);
nand U9710 (N_9710,N_9346,N_9357);
nand U9711 (N_9711,N_9392,N_9453);
nor U9712 (N_9712,N_9292,N_9341);
and U9713 (N_9713,N_9498,N_9403);
nor U9714 (N_9714,N_9417,N_9463);
or U9715 (N_9715,N_9330,N_9380);
nor U9716 (N_9716,N_9397,N_9387);
nand U9717 (N_9717,N_9261,N_9422);
nand U9718 (N_9718,N_9394,N_9391);
nand U9719 (N_9719,N_9431,N_9450);
nor U9720 (N_9720,N_9490,N_9314);
nor U9721 (N_9721,N_9396,N_9310);
nand U9722 (N_9722,N_9325,N_9487);
nor U9723 (N_9723,N_9274,N_9459);
or U9724 (N_9724,N_9337,N_9385);
and U9725 (N_9725,N_9459,N_9418);
and U9726 (N_9726,N_9439,N_9483);
nor U9727 (N_9727,N_9258,N_9344);
xnor U9728 (N_9728,N_9294,N_9349);
and U9729 (N_9729,N_9392,N_9299);
nand U9730 (N_9730,N_9426,N_9382);
and U9731 (N_9731,N_9488,N_9396);
nand U9732 (N_9732,N_9300,N_9277);
and U9733 (N_9733,N_9409,N_9446);
nand U9734 (N_9734,N_9263,N_9346);
nor U9735 (N_9735,N_9398,N_9444);
nor U9736 (N_9736,N_9376,N_9268);
nand U9737 (N_9737,N_9268,N_9484);
and U9738 (N_9738,N_9417,N_9273);
or U9739 (N_9739,N_9396,N_9279);
nor U9740 (N_9740,N_9465,N_9464);
nand U9741 (N_9741,N_9291,N_9490);
and U9742 (N_9742,N_9478,N_9315);
nor U9743 (N_9743,N_9371,N_9478);
and U9744 (N_9744,N_9308,N_9374);
nor U9745 (N_9745,N_9489,N_9338);
or U9746 (N_9746,N_9420,N_9355);
nor U9747 (N_9747,N_9343,N_9441);
nor U9748 (N_9748,N_9339,N_9307);
or U9749 (N_9749,N_9360,N_9463);
and U9750 (N_9750,N_9685,N_9614);
nor U9751 (N_9751,N_9505,N_9747);
nand U9752 (N_9752,N_9524,N_9626);
or U9753 (N_9753,N_9683,N_9735);
xor U9754 (N_9754,N_9669,N_9613);
or U9755 (N_9755,N_9672,N_9511);
nor U9756 (N_9756,N_9595,N_9738);
nand U9757 (N_9757,N_9500,N_9668);
nand U9758 (N_9758,N_9634,N_9562);
or U9759 (N_9759,N_9644,N_9604);
nand U9760 (N_9760,N_9633,N_9717);
nand U9761 (N_9761,N_9729,N_9627);
nor U9762 (N_9762,N_9581,N_9504);
nor U9763 (N_9763,N_9601,N_9661);
and U9764 (N_9764,N_9563,N_9646);
nand U9765 (N_9765,N_9515,N_9682);
or U9766 (N_9766,N_9579,N_9608);
nand U9767 (N_9767,N_9572,N_9700);
nor U9768 (N_9768,N_9609,N_9531);
or U9769 (N_9769,N_9673,N_9691);
and U9770 (N_9770,N_9707,N_9686);
nor U9771 (N_9771,N_9518,N_9720);
nor U9772 (N_9772,N_9605,N_9737);
nand U9773 (N_9773,N_9742,N_9630);
nor U9774 (N_9774,N_9573,N_9592);
or U9775 (N_9775,N_9612,N_9640);
or U9776 (N_9776,N_9526,N_9715);
and U9777 (N_9777,N_9674,N_9525);
nor U9778 (N_9778,N_9652,N_9694);
nand U9779 (N_9779,N_9582,N_9650);
nand U9780 (N_9780,N_9731,N_9701);
nand U9781 (N_9781,N_9624,N_9547);
and U9782 (N_9782,N_9665,N_9522);
nor U9783 (N_9783,N_9734,N_9680);
nand U9784 (N_9784,N_9539,N_9722);
or U9785 (N_9785,N_9559,N_9616);
nor U9786 (N_9786,N_9545,N_9659);
or U9787 (N_9787,N_9546,N_9656);
or U9788 (N_9788,N_9584,N_9567);
and U9789 (N_9789,N_9698,N_9708);
nand U9790 (N_9790,N_9723,N_9745);
nor U9791 (N_9791,N_9536,N_9712);
or U9792 (N_9792,N_9662,N_9615);
nor U9793 (N_9793,N_9543,N_9655);
and U9794 (N_9794,N_9578,N_9570);
and U9795 (N_9795,N_9693,N_9639);
nand U9796 (N_9796,N_9670,N_9599);
or U9797 (N_9797,N_9566,N_9696);
nor U9798 (N_9798,N_9519,N_9533);
nand U9799 (N_9799,N_9657,N_9704);
or U9800 (N_9800,N_9618,N_9689);
and U9801 (N_9801,N_9733,N_9607);
nand U9802 (N_9802,N_9621,N_9564);
nor U9803 (N_9803,N_9516,N_9552);
and U9804 (N_9804,N_9537,N_9663);
or U9805 (N_9805,N_9598,N_9549);
or U9806 (N_9806,N_9502,N_9544);
and U9807 (N_9807,N_9600,N_9538);
or U9808 (N_9808,N_9503,N_9679);
nand U9809 (N_9809,N_9638,N_9588);
nor U9810 (N_9810,N_9619,N_9594);
and U9811 (N_9811,N_9631,N_9535);
and U9812 (N_9812,N_9636,N_9664);
and U9813 (N_9813,N_9517,N_9681);
or U9814 (N_9814,N_9523,N_9643);
and U9815 (N_9815,N_9556,N_9576);
and U9816 (N_9816,N_9706,N_9611);
xnor U9817 (N_9817,N_9530,N_9590);
and U9818 (N_9818,N_9739,N_9645);
and U9819 (N_9819,N_9555,N_9577);
or U9820 (N_9820,N_9695,N_9560);
nor U9821 (N_9821,N_9711,N_9632);
or U9822 (N_9822,N_9724,N_9654);
nand U9823 (N_9823,N_9593,N_9730);
nor U9824 (N_9824,N_9529,N_9603);
or U9825 (N_9825,N_9744,N_9591);
nand U9826 (N_9826,N_9507,N_9716);
nand U9827 (N_9827,N_9623,N_9540);
or U9828 (N_9828,N_9521,N_9649);
or U9829 (N_9829,N_9565,N_9561);
or U9830 (N_9830,N_9727,N_9671);
or U9831 (N_9831,N_9541,N_9574);
or U9832 (N_9832,N_9617,N_9512);
and U9833 (N_9833,N_9667,N_9749);
and U9834 (N_9834,N_9713,N_9666);
and U9835 (N_9835,N_9554,N_9580);
nand U9836 (N_9836,N_9703,N_9575);
or U9837 (N_9837,N_9557,N_9651);
or U9838 (N_9838,N_9597,N_9508);
and U9839 (N_9839,N_9687,N_9709);
or U9840 (N_9840,N_9658,N_9569);
and U9841 (N_9841,N_9520,N_9510);
nand U9842 (N_9842,N_9642,N_9528);
nand U9843 (N_9843,N_9699,N_9660);
nand U9844 (N_9844,N_9558,N_9583);
nand U9845 (N_9845,N_9548,N_9585);
nand U9846 (N_9846,N_9748,N_9676);
and U9847 (N_9847,N_9688,N_9692);
nand U9848 (N_9848,N_9534,N_9736);
nor U9849 (N_9849,N_9506,N_9678);
and U9850 (N_9850,N_9653,N_9501);
nor U9851 (N_9851,N_9635,N_9527);
or U9852 (N_9852,N_9606,N_9718);
nor U9853 (N_9853,N_9714,N_9589);
nor U9854 (N_9854,N_9551,N_9625);
nand U9855 (N_9855,N_9702,N_9550);
or U9856 (N_9856,N_9610,N_9648);
nor U9857 (N_9857,N_9586,N_9628);
and U9858 (N_9858,N_9675,N_9641);
nor U9859 (N_9859,N_9725,N_9684);
and U9860 (N_9860,N_9647,N_9542);
nor U9861 (N_9861,N_9509,N_9553);
xnor U9862 (N_9862,N_9513,N_9602);
and U9863 (N_9863,N_9705,N_9568);
nand U9864 (N_9864,N_9697,N_9677);
and U9865 (N_9865,N_9571,N_9596);
nand U9866 (N_9866,N_9514,N_9629);
and U9867 (N_9867,N_9620,N_9719);
xor U9868 (N_9868,N_9732,N_9637);
or U9869 (N_9869,N_9622,N_9728);
and U9870 (N_9870,N_9721,N_9741);
or U9871 (N_9871,N_9532,N_9740);
nor U9872 (N_9872,N_9746,N_9690);
nor U9873 (N_9873,N_9743,N_9710);
and U9874 (N_9874,N_9726,N_9587);
and U9875 (N_9875,N_9554,N_9685);
and U9876 (N_9876,N_9512,N_9551);
nor U9877 (N_9877,N_9602,N_9564);
and U9878 (N_9878,N_9605,N_9713);
nor U9879 (N_9879,N_9623,N_9700);
and U9880 (N_9880,N_9557,N_9654);
and U9881 (N_9881,N_9689,N_9539);
nor U9882 (N_9882,N_9697,N_9592);
nand U9883 (N_9883,N_9601,N_9749);
nor U9884 (N_9884,N_9729,N_9518);
nand U9885 (N_9885,N_9716,N_9718);
and U9886 (N_9886,N_9657,N_9608);
or U9887 (N_9887,N_9644,N_9537);
and U9888 (N_9888,N_9705,N_9642);
nor U9889 (N_9889,N_9721,N_9529);
or U9890 (N_9890,N_9728,N_9546);
and U9891 (N_9891,N_9637,N_9639);
and U9892 (N_9892,N_9704,N_9748);
and U9893 (N_9893,N_9548,N_9711);
nand U9894 (N_9894,N_9609,N_9634);
or U9895 (N_9895,N_9620,N_9673);
and U9896 (N_9896,N_9740,N_9701);
nor U9897 (N_9897,N_9683,N_9528);
nor U9898 (N_9898,N_9726,N_9714);
or U9899 (N_9899,N_9632,N_9670);
or U9900 (N_9900,N_9667,N_9547);
nand U9901 (N_9901,N_9695,N_9592);
or U9902 (N_9902,N_9634,N_9727);
and U9903 (N_9903,N_9609,N_9543);
nor U9904 (N_9904,N_9626,N_9731);
nand U9905 (N_9905,N_9508,N_9699);
nand U9906 (N_9906,N_9715,N_9717);
xor U9907 (N_9907,N_9625,N_9713);
or U9908 (N_9908,N_9748,N_9652);
and U9909 (N_9909,N_9514,N_9620);
nor U9910 (N_9910,N_9605,N_9530);
and U9911 (N_9911,N_9629,N_9615);
or U9912 (N_9912,N_9584,N_9634);
nor U9913 (N_9913,N_9502,N_9685);
nand U9914 (N_9914,N_9593,N_9501);
or U9915 (N_9915,N_9732,N_9749);
and U9916 (N_9916,N_9564,N_9672);
and U9917 (N_9917,N_9714,N_9666);
and U9918 (N_9918,N_9649,N_9702);
or U9919 (N_9919,N_9716,N_9563);
or U9920 (N_9920,N_9636,N_9705);
or U9921 (N_9921,N_9585,N_9570);
nor U9922 (N_9922,N_9682,N_9542);
nand U9923 (N_9923,N_9616,N_9606);
or U9924 (N_9924,N_9716,N_9506);
nor U9925 (N_9925,N_9695,N_9649);
nor U9926 (N_9926,N_9528,N_9560);
or U9927 (N_9927,N_9587,N_9694);
nand U9928 (N_9928,N_9690,N_9741);
nand U9929 (N_9929,N_9605,N_9645);
nand U9930 (N_9930,N_9516,N_9656);
nor U9931 (N_9931,N_9569,N_9644);
nor U9932 (N_9932,N_9710,N_9602);
nor U9933 (N_9933,N_9541,N_9747);
and U9934 (N_9934,N_9706,N_9652);
nand U9935 (N_9935,N_9669,N_9620);
and U9936 (N_9936,N_9611,N_9538);
and U9937 (N_9937,N_9636,N_9505);
or U9938 (N_9938,N_9623,N_9612);
nand U9939 (N_9939,N_9588,N_9609);
and U9940 (N_9940,N_9706,N_9552);
nor U9941 (N_9941,N_9554,N_9680);
nand U9942 (N_9942,N_9699,N_9709);
nand U9943 (N_9943,N_9724,N_9503);
or U9944 (N_9944,N_9574,N_9620);
or U9945 (N_9945,N_9656,N_9631);
or U9946 (N_9946,N_9609,N_9692);
or U9947 (N_9947,N_9661,N_9551);
xor U9948 (N_9948,N_9730,N_9595);
or U9949 (N_9949,N_9506,N_9638);
or U9950 (N_9950,N_9508,N_9515);
or U9951 (N_9951,N_9653,N_9559);
and U9952 (N_9952,N_9709,N_9715);
nand U9953 (N_9953,N_9748,N_9637);
nor U9954 (N_9954,N_9681,N_9608);
nor U9955 (N_9955,N_9598,N_9632);
and U9956 (N_9956,N_9657,N_9712);
and U9957 (N_9957,N_9633,N_9514);
or U9958 (N_9958,N_9723,N_9743);
or U9959 (N_9959,N_9658,N_9657);
and U9960 (N_9960,N_9621,N_9697);
or U9961 (N_9961,N_9749,N_9619);
xnor U9962 (N_9962,N_9726,N_9524);
and U9963 (N_9963,N_9542,N_9578);
and U9964 (N_9964,N_9717,N_9628);
or U9965 (N_9965,N_9567,N_9588);
or U9966 (N_9966,N_9533,N_9696);
and U9967 (N_9967,N_9598,N_9516);
nor U9968 (N_9968,N_9555,N_9504);
and U9969 (N_9969,N_9552,N_9596);
nand U9970 (N_9970,N_9602,N_9613);
and U9971 (N_9971,N_9674,N_9702);
or U9972 (N_9972,N_9506,N_9670);
or U9973 (N_9973,N_9572,N_9666);
and U9974 (N_9974,N_9501,N_9586);
nand U9975 (N_9975,N_9527,N_9664);
nand U9976 (N_9976,N_9620,N_9613);
nand U9977 (N_9977,N_9526,N_9531);
or U9978 (N_9978,N_9736,N_9564);
or U9979 (N_9979,N_9649,N_9512);
and U9980 (N_9980,N_9566,N_9697);
nor U9981 (N_9981,N_9593,N_9613);
nand U9982 (N_9982,N_9507,N_9683);
nand U9983 (N_9983,N_9509,N_9603);
nand U9984 (N_9984,N_9542,N_9630);
or U9985 (N_9985,N_9696,N_9519);
xor U9986 (N_9986,N_9602,N_9672);
nor U9987 (N_9987,N_9709,N_9707);
nand U9988 (N_9988,N_9576,N_9524);
nor U9989 (N_9989,N_9593,N_9638);
or U9990 (N_9990,N_9668,N_9715);
nor U9991 (N_9991,N_9569,N_9583);
nor U9992 (N_9992,N_9716,N_9586);
nor U9993 (N_9993,N_9656,N_9504);
and U9994 (N_9994,N_9696,N_9647);
nor U9995 (N_9995,N_9738,N_9552);
nor U9996 (N_9996,N_9537,N_9584);
nand U9997 (N_9997,N_9595,N_9681);
or U9998 (N_9998,N_9700,N_9591);
nand U9999 (N_9999,N_9532,N_9584);
or U10000 (N_10000,N_9884,N_9775);
nor U10001 (N_10001,N_9948,N_9906);
or U10002 (N_10002,N_9769,N_9944);
nor U10003 (N_10003,N_9890,N_9964);
nand U10004 (N_10004,N_9959,N_9903);
nor U10005 (N_10005,N_9953,N_9822);
nand U10006 (N_10006,N_9874,N_9770);
or U10007 (N_10007,N_9897,N_9970);
or U10008 (N_10008,N_9788,N_9753);
or U10009 (N_10009,N_9836,N_9973);
and U10010 (N_10010,N_9804,N_9911);
or U10011 (N_10011,N_9875,N_9885);
nand U10012 (N_10012,N_9821,N_9872);
nand U10013 (N_10013,N_9950,N_9998);
nor U10014 (N_10014,N_9812,N_9779);
and U10015 (N_10015,N_9814,N_9777);
nor U10016 (N_10016,N_9895,N_9800);
xnor U10017 (N_10017,N_9947,N_9977);
nor U10018 (N_10018,N_9926,N_9923);
nand U10019 (N_10019,N_9830,N_9837);
xnor U10020 (N_10020,N_9912,N_9939);
or U10021 (N_10021,N_9886,N_9825);
nor U10022 (N_10022,N_9924,N_9856);
or U10023 (N_10023,N_9920,N_9986);
and U10024 (N_10024,N_9867,N_9975);
nor U10025 (N_10025,N_9966,N_9847);
or U10026 (N_10026,N_9853,N_9983);
and U10027 (N_10027,N_9982,N_9971);
and U10028 (N_10028,N_9991,N_9857);
nand U10029 (N_10029,N_9802,N_9962);
nand U10030 (N_10030,N_9976,N_9797);
and U10031 (N_10031,N_9918,N_9900);
or U10032 (N_10032,N_9756,N_9793);
and U10033 (N_10033,N_9784,N_9930);
or U10034 (N_10034,N_9870,N_9901);
xor U10035 (N_10035,N_9844,N_9762);
or U10036 (N_10036,N_9809,N_9915);
or U10037 (N_10037,N_9798,N_9913);
and U10038 (N_10038,N_9969,N_9832);
nand U10039 (N_10039,N_9820,N_9956);
nor U10040 (N_10040,N_9805,N_9979);
nand U10041 (N_10041,N_9851,N_9808);
nand U10042 (N_10042,N_9877,N_9841);
or U10043 (N_10043,N_9878,N_9910);
or U10044 (N_10044,N_9978,N_9790);
xnor U10045 (N_10045,N_9771,N_9985);
and U10046 (N_10046,N_9785,N_9869);
or U10047 (N_10047,N_9866,N_9904);
nand U10048 (N_10048,N_9778,N_9794);
nand U10049 (N_10049,N_9787,N_9846);
nand U10050 (N_10050,N_9834,N_9907);
and U10051 (N_10051,N_9993,N_9781);
and U10052 (N_10052,N_9984,N_9859);
nand U10053 (N_10053,N_9819,N_9765);
or U10054 (N_10054,N_9842,N_9955);
xnor U10055 (N_10055,N_9916,N_9861);
or U10056 (N_10056,N_9854,N_9750);
or U10057 (N_10057,N_9943,N_9908);
or U10058 (N_10058,N_9954,N_9999);
nand U10059 (N_10059,N_9888,N_9782);
nor U10060 (N_10060,N_9925,N_9795);
and U10061 (N_10061,N_9933,N_9806);
nand U10062 (N_10062,N_9965,N_9768);
and U10063 (N_10063,N_9937,N_9810);
nor U10064 (N_10064,N_9772,N_9921);
or U10065 (N_10065,N_9848,N_9989);
nor U10066 (N_10066,N_9791,N_9942);
nand U10067 (N_10067,N_9946,N_9899);
nor U10068 (N_10068,N_9817,N_9862);
or U10069 (N_10069,N_9751,N_9839);
nor U10070 (N_10070,N_9893,N_9776);
or U10071 (N_10071,N_9881,N_9880);
nand U10072 (N_10072,N_9811,N_9882);
and U10073 (N_10073,N_9958,N_9871);
and U10074 (N_10074,N_9868,N_9941);
or U10075 (N_10075,N_9894,N_9818);
nor U10076 (N_10076,N_9988,N_9754);
nor U10077 (N_10077,N_9865,N_9951);
nand U10078 (N_10078,N_9972,N_9849);
xor U10079 (N_10079,N_9758,N_9760);
nor U10080 (N_10080,N_9952,N_9833);
and U10081 (N_10081,N_9914,N_9963);
nand U10082 (N_10082,N_9934,N_9807);
or U10083 (N_10083,N_9783,N_9992);
nand U10084 (N_10084,N_9891,N_9995);
or U10085 (N_10085,N_9902,N_9889);
nor U10086 (N_10086,N_9940,N_9997);
nor U10087 (N_10087,N_9932,N_9845);
or U10088 (N_10088,N_9815,N_9829);
nand U10089 (N_10089,N_9968,N_9835);
or U10090 (N_10090,N_9974,N_9828);
nor U10091 (N_10091,N_9838,N_9858);
nand U10092 (N_10092,N_9766,N_9792);
and U10093 (N_10093,N_9813,N_9987);
nor U10094 (N_10094,N_9981,N_9864);
nor U10095 (N_10095,N_9945,N_9761);
or U10096 (N_10096,N_9764,N_9990);
or U10097 (N_10097,N_9801,N_9831);
nor U10098 (N_10098,N_9892,N_9773);
and U10099 (N_10099,N_9996,N_9850);
nand U10100 (N_10100,N_9759,N_9961);
nor U10101 (N_10101,N_9980,N_9927);
and U10102 (N_10102,N_9757,N_9905);
or U10103 (N_10103,N_9789,N_9938);
nor U10104 (N_10104,N_9898,N_9957);
nor U10105 (N_10105,N_9967,N_9826);
and U10106 (N_10106,N_9823,N_9917);
nand U10107 (N_10107,N_9767,N_9799);
or U10108 (N_10108,N_9879,N_9929);
or U10109 (N_10109,N_9763,N_9824);
nor U10110 (N_10110,N_9896,N_9827);
nor U10111 (N_10111,N_9840,N_9786);
nor U10112 (N_10112,N_9928,N_9873);
and U10113 (N_10113,N_9935,N_9843);
and U10114 (N_10114,N_9816,N_9796);
and U10115 (N_10115,N_9876,N_9855);
nor U10116 (N_10116,N_9919,N_9755);
nor U10117 (N_10117,N_9752,N_9931);
and U10118 (N_10118,N_9803,N_9863);
nand U10119 (N_10119,N_9949,N_9887);
nand U10120 (N_10120,N_9774,N_9994);
and U10121 (N_10121,N_9883,N_9922);
nand U10122 (N_10122,N_9780,N_9909);
xor U10123 (N_10123,N_9860,N_9936);
nand U10124 (N_10124,N_9960,N_9852);
nor U10125 (N_10125,N_9796,N_9787);
nand U10126 (N_10126,N_9878,N_9867);
nand U10127 (N_10127,N_9864,N_9860);
and U10128 (N_10128,N_9962,N_9906);
nand U10129 (N_10129,N_9851,N_9841);
or U10130 (N_10130,N_9753,N_9821);
or U10131 (N_10131,N_9776,N_9977);
and U10132 (N_10132,N_9874,N_9996);
or U10133 (N_10133,N_9930,N_9881);
nand U10134 (N_10134,N_9815,N_9885);
and U10135 (N_10135,N_9873,N_9781);
and U10136 (N_10136,N_9945,N_9934);
and U10137 (N_10137,N_9981,N_9938);
and U10138 (N_10138,N_9779,N_9922);
and U10139 (N_10139,N_9758,N_9792);
and U10140 (N_10140,N_9819,N_9812);
and U10141 (N_10141,N_9839,N_9920);
and U10142 (N_10142,N_9909,N_9914);
and U10143 (N_10143,N_9938,N_9844);
nand U10144 (N_10144,N_9922,N_9795);
nor U10145 (N_10145,N_9863,N_9851);
xor U10146 (N_10146,N_9793,N_9950);
xnor U10147 (N_10147,N_9845,N_9963);
or U10148 (N_10148,N_9851,N_9844);
nand U10149 (N_10149,N_9994,N_9767);
and U10150 (N_10150,N_9987,N_9824);
nand U10151 (N_10151,N_9758,N_9889);
nor U10152 (N_10152,N_9966,N_9956);
and U10153 (N_10153,N_9902,N_9966);
or U10154 (N_10154,N_9898,N_9914);
or U10155 (N_10155,N_9976,N_9954);
and U10156 (N_10156,N_9974,N_9768);
nand U10157 (N_10157,N_9957,N_9839);
or U10158 (N_10158,N_9902,N_9918);
nor U10159 (N_10159,N_9963,N_9850);
nor U10160 (N_10160,N_9880,N_9815);
nor U10161 (N_10161,N_9897,N_9987);
or U10162 (N_10162,N_9764,N_9863);
nor U10163 (N_10163,N_9772,N_9990);
or U10164 (N_10164,N_9945,N_9861);
and U10165 (N_10165,N_9940,N_9927);
nor U10166 (N_10166,N_9827,N_9972);
nor U10167 (N_10167,N_9930,N_9862);
nand U10168 (N_10168,N_9855,N_9830);
nor U10169 (N_10169,N_9900,N_9937);
or U10170 (N_10170,N_9814,N_9771);
nor U10171 (N_10171,N_9955,N_9801);
and U10172 (N_10172,N_9965,N_9860);
and U10173 (N_10173,N_9974,N_9964);
nor U10174 (N_10174,N_9969,N_9903);
nand U10175 (N_10175,N_9885,N_9943);
or U10176 (N_10176,N_9856,N_9797);
nor U10177 (N_10177,N_9935,N_9832);
and U10178 (N_10178,N_9807,N_9865);
nor U10179 (N_10179,N_9766,N_9757);
nand U10180 (N_10180,N_9954,N_9923);
nand U10181 (N_10181,N_9874,N_9969);
nor U10182 (N_10182,N_9910,N_9758);
and U10183 (N_10183,N_9819,N_9807);
and U10184 (N_10184,N_9824,N_9778);
nand U10185 (N_10185,N_9824,N_9837);
nor U10186 (N_10186,N_9956,N_9977);
nand U10187 (N_10187,N_9905,N_9795);
and U10188 (N_10188,N_9961,N_9958);
nor U10189 (N_10189,N_9812,N_9959);
nor U10190 (N_10190,N_9830,N_9854);
nand U10191 (N_10191,N_9936,N_9816);
nor U10192 (N_10192,N_9768,N_9825);
and U10193 (N_10193,N_9876,N_9882);
nand U10194 (N_10194,N_9828,N_9985);
nor U10195 (N_10195,N_9990,N_9906);
and U10196 (N_10196,N_9959,N_9835);
nor U10197 (N_10197,N_9833,N_9770);
nor U10198 (N_10198,N_9822,N_9892);
nor U10199 (N_10199,N_9910,N_9949);
nand U10200 (N_10200,N_9952,N_9797);
nor U10201 (N_10201,N_9835,N_9828);
and U10202 (N_10202,N_9987,N_9819);
and U10203 (N_10203,N_9875,N_9790);
nand U10204 (N_10204,N_9931,N_9847);
and U10205 (N_10205,N_9883,N_9782);
and U10206 (N_10206,N_9967,N_9980);
and U10207 (N_10207,N_9845,N_9906);
xnor U10208 (N_10208,N_9841,N_9902);
or U10209 (N_10209,N_9932,N_9959);
and U10210 (N_10210,N_9831,N_9778);
and U10211 (N_10211,N_9908,N_9882);
and U10212 (N_10212,N_9871,N_9890);
nand U10213 (N_10213,N_9816,N_9904);
nand U10214 (N_10214,N_9823,N_9904);
nor U10215 (N_10215,N_9797,N_9769);
and U10216 (N_10216,N_9898,N_9981);
and U10217 (N_10217,N_9968,N_9847);
and U10218 (N_10218,N_9966,N_9791);
xnor U10219 (N_10219,N_9892,N_9974);
nor U10220 (N_10220,N_9926,N_9765);
nor U10221 (N_10221,N_9789,N_9882);
and U10222 (N_10222,N_9827,N_9757);
or U10223 (N_10223,N_9803,N_9858);
and U10224 (N_10224,N_9859,N_9974);
and U10225 (N_10225,N_9905,N_9915);
and U10226 (N_10226,N_9937,N_9856);
and U10227 (N_10227,N_9876,N_9877);
nand U10228 (N_10228,N_9826,N_9768);
and U10229 (N_10229,N_9953,N_9952);
or U10230 (N_10230,N_9875,N_9841);
nand U10231 (N_10231,N_9779,N_9936);
nand U10232 (N_10232,N_9858,N_9771);
or U10233 (N_10233,N_9993,N_9818);
nor U10234 (N_10234,N_9905,N_9895);
nor U10235 (N_10235,N_9857,N_9898);
and U10236 (N_10236,N_9773,N_9939);
nand U10237 (N_10237,N_9895,N_9919);
nor U10238 (N_10238,N_9929,N_9869);
nor U10239 (N_10239,N_9977,N_9951);
nor U10240 (N_10240,N_9837,N_9816);
and U10241 (N_10241,N_9854,N_9943);
nand U10242 (N_10242,N_9874,N_9784);
or U10243 (N_10243,N_9960,N_9804);
or U10244 (N_10244,N_9899,N_9849);
nor U10245 (N_10245,N_9806,N_9849);
or U10246 (N_10246,N_9944,N_9990);
and U10247 (N_10247,N_9834,N_9883);
or U10248 (N_10248,N_9853,N_9847);
or U10249 (N_10249,N_9751,N_9971);
nand U10250 (N_10250,N_10117,N_10165);
nand U10251 (N_10251,N_10145,N_10043);
nor U10252 (N_10252,N_10130,N_10197);
nor U10253 (N_10253,N_10039,N_10086);
nand U10254 (N_10254,N_10238,N_10021);
nor U10255 (N_10255,N_10074,N_10060);
xor U10256 (N_10256,N_10095,N_10153);
or U10257 (N_10257,N_10027,N_10026);
or U10258 (N_10258,N_10211,N_10169);
and U10259 (N_10259,N_10067,N_10133);
and U10260 (N_10260,N_10141,N_10065);
and U10261 (N_10261,N_10108,N_10122);
and U10262 (N_10262,N_10225,N_10109);
or U10263 (N_10263,N_10177,N_10012);
or U10264 (N_10264,N_10161,N_10030);
xnor U10265 (N_10265,N_10119,N_10000);
or U10266 (N_10266,N_10055,N_10099);
and U10267 (N_10267,N_10227,N_10050);
nor U10268 (N_10268,N_10001,N_10092);
or U10269 (N_10269,N_10113,N_10104);
and U10270 (N_10270,N_10062,N_10068);
nand U10271 (N_10271,N_10129,N_10041);
and U10272 (N_10272,N_10214,N_10193);
nor U10273 (N_10273,N_10066,N_10191);
nand U10274 (N_10274,N_10172,N_10102);
and U10275 (N_10275,N_10024,N_10085);
and U10276 (N_10276,N_10200,N_10002);
nand U10277 (N_10277,N_10090,N_10151);
and U10278 (N_10278,N_10152,N_10166);
nor U10279 (N_10279,N_10233,N_10044);
nor U10280 (N_10280,N_10243,N_10036);
and U10281 (N_10281,N_10244,N_10049);
or U10282 (N_10282,N_10134,N_10140);
nor U10283 (N_10283,N_10196,N_10208);
nand U10284 (N_10284,N_10112,N_10170);
or U10285 (N_10285,N_10031,N_10042);
xor U10286 (N_10286,N_10046,N_10038);
and U10287 (N_10287,N_10162,N_10216);
nor U10288 (N_10288,N_10073,N_10159);
and U10289 (N_10289,N_10123,N_10082);
nand U10290 (N_10290,N_10063,N_10096);
nor U10291 (N_10291,N_10023,N_10246);
nand U10292 (N_10292,N_10081,N_10198);
nand U10293 (N_10293,N_10051,N_10157);
or U10294 (N_10294,N_10004,N_10236);
nand U10295 (N_10295,N_10148,N_10107);
and U10296 (N_10296,N_10127,N_10235);
nor U10297 (N_10297,N_10218,N_10237);
or U10298 (N_10298,N_10014,N_10245);
nand U10299 (N_10299,N_10105,N_10192);
nand U10300 (N_10300,N_10242,N_10158);
and U10301 (N_10301,N_10204,N_10138);
or U10302 (N_10302,N_10248,N_10135);
nand U10303 (N_10303,N_10019,N_10028);
nand U10304 (N_10304,N_10059,N_10173);
and U10305 (N_10305,N_10220,N_10022);
nor U10306 (N_10306,N_10006,N_10229);
nand U10307 (N_10307,N_10056,N_10226);
or U10308 (N_10308,N_10175,N_10201);
and U10309 (N_10309,N_10247,N_10013);
or U10310 (N_10310,N_10185,N_10075);
and U10311 (N_10311,N_10116,N_10215);
nand U10312 (N_10312,N_10020,N_10144);
or U10313 (N_10313,N_10155,N_10132);
or U10314 (N_10314,N_10091,N_10210);
or U10315 (N_10315,N_10111,N_10234);
and U10316 (N_10316,N_10183,N_10047);
or U10317 (N_10317,N_10212,N_10222);
or U10318 (N_10318,N_10121,N_10174);
and U10319 (N_10319,N_10190,N_10205);
nand U10320 (N_10320,N_10057,N_10149);
and U10321 (N_10321,N_10064,N_10098);
or U10322 (N_10322,N_10032,N_10053);
and U10323 (N_10323,N_10194,N_10182);
nand U10324 (N_10324,N_10137,N_10224);
or U10325 (N_10325,N_10131,N_10093);
nand U10326 (N_10326,N_10146,N_10106);
or U10327 (N_10327,N_10156,N_10241);
nor U10328 (N_10328,N_10094,N_10048);
or U10329 (N_10329,N_10180,N_10100);
nor U10330 (N_10330,N_10150,N_10209);
and U10331 (N_10331,N_10163,N_10025);
xnor U10332 (N_10332,N_10097,N_10035);
and U10333 (N_10333,N_10219,N_10178);
nand U10334 (N_10334,N_10018,N_10088);
and U10335 (N_10335,N_10072,N_10167);
or U10336 (N_10336,N_10239,N_10179);
nor U10337 (N_10337,N_10009,N_10213);
and U10338 (N_10338,N_10176,N_10223);
and U10339 (N_10339,N_10003,N_10101);
and U10340 (N_10340,N_10118,N_10083);
and U10341 (N_10341,N_10040,N_10015);
nor U10342 (N_10342,N_10069,N_10171);
nor U10343 (N_10343,N_10240,N_10142);
and U10344 (N_10344,N_10011,N_10115);
nor U10345 (N_10345,N_10079,N_10007);
or U10346 (N_10346,N_10199,N_10168);
nand U10347 (N_10347,N_10249,N_10181);
and U10348 (N_10348,N_10037,N_10184);
or U10349 (N_10349,N_10110,N_10160);
nand U10350 (N_10350,N_10124,N_10207);
and U10351 (N_10351,N_10189,N_10058);
or U10352 (N_10352,N_10232,N_10010);
or U10353 (N_10353,N_10061,N_10080);
and U10354 (N_10354,N_10217,N_10136);
and U10355 (N_10355,N_10008,N_10120);
and U10356 (N_10356,N_10126,N_10078);
or U10357 (N_10357,N_10052,N_10230);
or U10358 (N_10358,N_10231,N_10206);
and U10359 (N_10359,N_10202,N_10164);
nor U10360 (N_10360,N_10071,N_10188);
and U10361 (N_10361,N_10034,N_10045);
and U10362 (N_10362,N_10029,N_10016);
and U10363 (N_10363,N_10070,N_10084);
nand U10364 (N_10364,N_10154,N_10203);
nor U10365 (N_10365,N_10125,N_10076);
or U10366 (N_10366,N_10114,N_10033);
or U10367 (N_10367,N_10054,N_10143);
or U10368 (N_10368,N_10017,N_10128);
nor U10369 (N_10369,N_10005,N_10221);
nand U10370 (N_10370,N_10147,N_10103);
nor U10371 (N_10371,N_10077,N_10195);
xnor U10372 (N_10372,N_10228,N_10087);
nand U10373 (N_10373,N_10187,N_10186);
or U10374 (N_10374,N_10089,N_10139);
nor U10375 (N_10375,N_10159,N_10106);
or U10376 (N_10376,N_10145,N_10079);
and U10377 (N_10377,N_10192,N_10202);
nor U10378 (N_10378,N_10248,N_10106);
nand U10379 (N_10379,N_10057,N_10226);
and U10380 (N_10380,N_10001,N_10004);
nand U10381 (N_10381,N_10103,N_10093);
or U10382 (N_10382,N_10237,N_10178);
or U10383 (N_10383,N_10030,N_10197);
and U10384 (N_10384,N_10000,N_10194);
nand U10385 (N_10385,N_10185,N_10012);
or U10386 (N_10386,N_10218,N_10060);
and U10387 (N_10387,N_10245,N_10019);
and U10388 (N_10388,N_10239,N_10059);
or U10389 (N_10389,N_10113,N_10093);
nor U10390 (N_10390,N_10016,N_10186);
nor U10391 (N_10391,N_10164,N_10100);
nor U10392 (N_10392,N_10248,N_10090);
nor U10393 (N_10393,N_10122,N_10081);
nor U10394 (N_10394,N_10225,N_10124);
or U10395 (N_10395,N_10124,N_10230);
xor U10396 (N_10396,N_10197,N_10163);
and U10397 (N_10397,N_10046,N_10136);
nor U10398 (N_10398,N_10044,N_10199);
nand U10399 (N_10399,N_10124,N_10152);
and U10400 (N_10400,N_10019,N_10007);
and U10401 (N_10401,N_10166,N_10179);
and U10402 (N_10402,N_10107,N_10084);
xnor U10403 (N_10403,N_10207,N_10112);
xnor U10404 (N_10404,N_10112,N_10233);
nor U10405 (N_10405,N_10076,N_10163);
nand U10406 (N_10406,N_10002,N_10179);
and U10407 (N_10407,N_10000,N_10245);
or U10408 (N_10408,N_10226,N_10178);
and U10409 (N_10409,N_10097,N_10176);
and U10410 (N_10410,N_10086,N_10160);
or U10411 (N_10411,N_10023,N_10094);
and U10412 (N_10412,N_10027,N_10210);
nor U10413 (N_10413,N_10167,N_10230);
or U10414 (N_10414,N_10040,N_10201);
and U10415 (N_10415,N_10143,N_10194);
nand U10416 (N_10416,N_10057,N_10064);
nand U10417 (N_10417,N_10177,N_10234);
and U10418 (N_10418,N_10021,N_10154);
nor U10419 (N_10419,N_10091,N_10001);
nand U10420 (N_10420,N_10231,N_10103);
or U10421 (N_10421,N_10170,N_10078);
nor U10422 (N_10422,N_10094,N_10117);
nand U10423 (N_10423,N_10085,N_10206);
or U10424 (N_10424,N_10094,N_10026);
nor U10425 (N_10425,N_10208,N_10214);
and U10426 (N_10426,N_10155,N_10241);
nor U10427 (N_10427,N_10069,N_10191);
nand U10428 (N_10428,N_10112,N_10047);
nor U10429 (N_10429,N_10096,N_10217);
nor U10430 (N_10430,N_10200,N_10180);
or U10431 (N_10431,N_10220,N_10232);
and U10432 (N_10432,N_10170,N_10140);
and U10433 (N_10433,N_10088,N_10236);
nand U10434 (N_10434,N_10122,N_10024);
and U10435 (N_10435,N_10064,N_10013);
nor U10436 (N_10436,N_10004,N_10212);
and U10437 (N_10437,N_10173,N_10236);
nor U10438 (N_10438,N_10035,N_10179);
nor U10439 (N_10439,N_10147,N_10034);
nand U10440 (N_10440,N_10087,N_10120);
or U10441 (N_10441,N_10225,N_10168);
nand U10442 (N_10442,N_10135,N_10147);
nand U10443 (N_10443,N_10055,N_10062);
nor U10444 (N_10444,N_10245,N_10057);
or U10445 (N_10445,N_10035,N_10219);
nor U10446 (N_10446,N_10132,N_10187);
nor U10447 (N_10447,N_10094,N_10200);
or U10448 (N_10448,N_10223,N_10166);
nor U10449 (N_10449,N_10174,N_10041);
or U10450 (N_10450,N_10053,N_10203);
or U10451 (N_10451,N_10075,N_10028);
nor U10452 (N_10452,N_10057,N_10163);
nand U10453 (N_10453,N_10176,N_10065);
and U10454 (N_10454,N_10181,N_10201);
and U10455 (N_10455,N_10022,N_10053);
and U10456 (N_10456,N_10043,N_10183);
and U10457 (N_10457,N_10134,N_10061);
and U10458 (N_10458,N_10170,N_10002);
or U10459 (N_10459,N_10070,N_10035);
nor U10460 (N_10460,N_10218,N_10071);
nor U10461 (N_10461,N_10008,N_10124);
and U10462 (N_10462,N_10081,N_10007);
nand U10463 (N_10463,N_10005,N_10096);
and U10464 (N_10464,N_10237,N_10222);
nand U10465 (N_10465,N_10165,N_10197);
or U10466 (N_10466,N_10095,N_10131);
nand U10467 (N_10467,N_10046,N_10080);
xor U10468 (N_10468,N_10111,N_10045);
nand U10469 (N_10469,N_10022,N_10195);
and U10470 (N_10470,N_10078,N_10014);
and U10471 (N_10471,N_10135,N_10125);
nand U10472 (N_10472,N_10132,N_10177);
and U10473 (N_10473,N_10068,N_10161);
nand U10474 (N_10474,N_10160,N_10007);
xnor U10475 (N_10475,N_10111,N_10196);
or U10476 (N_10476,N_10061,N_10215);
or U10477 (N_10477,N_10025,N_10234);
and U10478 (N_10478,N_10129,N_10211);
nand U10479 (N_10479,N_10067,N_10191);
and U10480 (N_10480,N_10121,N_10215);
nand U10481 (N_10481,N_10128,N_10133);
and U10482 (N_10482,N_10213,N_10206);
nand U10483 (N_10483,N_10035,N_10019);
and U10484 (N_10484,N_10188,N_10091);
nand U10485 (N_10485,N_10031,N_10154);
xnor U10486 (N_10486,N_10001,N_10239);
and U10487 (N_10487,N_10093,N_10158);
or U10488 (N_10488,N_10150,N_10049);
and U10489 (N_10489,N_10071,N_10010);
nor U10490 (N_10490,N_10198,N_10200);
nor U10491 (N_10491,N_10144,N_10071);
nand U10492 (N_10492,N_10155,N_10118);
or U10493 (N_10493,N_10010,N_10208);
or U10494 (N_10494,N_10105,N_10005);
nor U10495 (N_10495,N_10063,N_10169);
or U10496 (N_10496,N_10235,N_10164);
and U10497 (N_10497,N_10132,N_10223);
and U10498 (N_10498,N_10201,N_10187);
nor U10499 (N_10499,N_10154,N_10208);
nor U10500 (N_10500,N_10362,N_10298);
and U10501 (N_10501,N_10251,N_10486);
and U10502 (N_10502,N_10262,N_10358);
or U10503 (N_10503,N_10261,N_10311);
and U10504 (N_10504,N_10332,N_10272);
nand U10505 (N_10505,N_10338,N_10283);
nor U10506 (N_10506,N_10468,N_10340);
or U10507 (N_10507,N_10309,N_10394);
or U10508 (N_10508,N_10315,N_10476);
xor U10509 (N_10509,N_10418,N_10347);
or U10510 (N_10510,N_10491,N_10482);
nor U10511 (N_10511,N_10438,N_10444);
nor U10512 (N_10512,N_10378,N_10307);
nor U10513 (N_10513,N_10286,N_10327);
and U10514 (N_10514,N_10404,N_10429);
or U10515 (N_10515,N_10260,N_10453);
nand U10516 (N_10516,N_10254,N_10289);
nand U10517 (N_10517,N_10353,N_10398);
nor U10518 (N_10518,N_10462,N_10496);
and U10519 (N_10519,N_10250,N_10348);
and U10520 (N_10520,N_10425,N_10379);
nand U10521 (N_10521,N_10451,N_10339);
and U10522 (N_10522,N_10352,N_10382);
and U10523 (N_10523,N_10478,N_10320);
nand U10524 (N_10524,N_10368,N_10492);
nand U10525 (N_10525,N_10393,N_10278);
or U10526 (N_10526,N_10269,N_10414);
and U10527 (N_10527,N_10469,N_10275);
nor U10528 (N_10528,N_10428,N_10480);
nand U10529 (N_10529,N_10433,N_10421);
and U10530 (N_10530,N_10384,N_10360);
nand U10531 (N_10531,N_10460,N_10439);
nand U10532 (N_10532,N_10333,N_10493);
nand U10533 (N_10533,N_10255,N_10411);
nand U10534 (N_10534,N_10291,N_10316);
nor U10535 (N_10535,N_10461,N_10455);
or U10536 (N_10536,N_10489,N_10456);
and U10537 (N_10537,N_10483,N_10390);
and U10538 (N_10538,N_10389,N_10268);
or U10539 (N_10539,N_10424,N_10285);
nor U10540 (N_10540,N_10473,N_10299);
or U10541 (N_10541,N_10446,N_10463);
nand U10542 (N_10542,N_10331,N_10434);
nor U10543 (N_10543,N_10319,N_10498);
nor U10544 (N_10544,N_10426,N_10450);
xor U10545 (N_10545,N_10487,N_10467);
or U10546 (N_10546,N_10263,N_10448);
or U10547 (N_10547,N_10363,N_10313);
xor U10548 (N_10548,N_10397,N_10387);
and U10549 (N_10549,N_10396,N_10284);
nand U10550 (N_10550,N_10335,N_10371);
or U10551 (N_10551,N_10395,N_10290);
and U10552 (N_10552,N_10321,N_10310);
and U10553 (N_10553,N_10343,N_10372);
and U10554 (N_10554,N_10485,N_10256);
or U10555 (N_10555,N_10419,N_10452);
or U10556 (N_10556,N_10258,N_10479);
and U10557 (N_10557,N_10465,N_10477);
nand U10558 (N_10558,N_10364,N_10351);
and U10559 (N_10559,N_10447,N_10361);
xor U10560 (N_10560,N_10430,N_10322);
nand U10561 (N_10561,N_10474,N_10253);
and U10562 (N_10562,N_10345,N_10306);
or U10563 (N_10563,N_10303,N_10296);
nand U10564 (N_10564,N_10427,N_10386);
or U10565 (N_10565,N_10385,N_10472);
or U10566 (N_10566,N_10301,N_10417);
or U10567 (N_10567,N_10350,N_10470);
or U10568 (N_10568,N_10406,N_10399);
xor U10569 (N_10569,N_10449,N_10366);
or U10570 (N_10570,N_10494,N_10317);
and U10571 (N_10571,N_10435,N_10423);
and U10572 (N_10572,N_10356,N_10374);
or U10573 (N_10573,N_10330,N_10266);
nor U10574 (N_10574,N_10293,N_10415);
or U10575 (N_10575,N_10481,N_10369);
nand U10576 (N_10576,N_10323,N_10497);
and U10577 (N_10577,N_10302,N_10308);
nor U10578 (N_10578,N_10341,N_10270);
or U10579 (N_10579,N_10416,N_10454);
and U10580 (N_10580,N_10292,N_10495);
and U10581 (N_10581,N_10388,N_10376);
and U10582 (N_10582,N_10412,N_10324);
nand U10583 (N_10583,N_10377,N_10294);
and U10584 (N_10584,N_10471,N_10466);
or U10585 (N_10585,N_10354,N_10392);
or U10586 (N_10586,N_10304,N_10305);
and U10587 (N_10587,N_10405,N_10484);
nand U10588 (N_10588,N_10349,N_10312);
nand U10589 (N_10589,N_10420,N_10314);
nor U10590 (N_10590,N_10442,N_10445);
or U10591 (N_10591,N_10437,N_10365);
or U10592 (N_10592,N_10432,N_10267);
nand U10593 (N_10593,N_10300,N_10328);
and U10594 (N_10594,N_10464,N_10337);
nand U10595 (N_10595,N_10488,N_10422);
and U10596 (N_10596,N_10401,N_10279);
and U10597 (N_10597,N_10281,N_10499);
or U10598 (N_10598,N_10344,N_10391);
nand U10599 (N_10599,N_10359,N_10274);
and U10600 (N_10600,N_10431,N_10370);
nor U10601 (N_10601,N_10413,N_10402);
and U10602 (N_10602,N_10282,N_10458);
and U10603 (N_10603,N_10409,N_10408);
or U10604 (N_10604,N_10457,N_10297);
and U10605 (N_10605,N_10329,N_10441);
nor U10606 (N_10606,N_10407,N_10273);
nor U10607 (N_10607,N_10295,N_10346);
and U10608 (N_10608,N_10288,N_10318);
and U10609 (N_10609,N_10475,N_10280);
or U10610 (N_10610,N_10334,N_10443);
nor U10611 (N_10611,N_10265,N_10276);
nor U10612 (N_10612,N_10375,N_10325);
or U10613 (N_10613,N_10271,N_10336);
nor U10614 (N_10614,N_10357,N_10367);
nor U10615 (N_10615,N_10380,N_10287);
and U10616 (N_10616,N_10490,N_10400);
and U10617 (N_10617,N_10252,N_10257);
nand U10618 (N_10618,N_10277,N_10326);
nor U10619 (N_10619,N_10381,N_10383);
and U10620 (N_10620,N_10403,N_10259);
nand U10621 (N_10621,N_10342,N_10373);
or U10622 (N_10622,N_10440,N_10264);
nand U10623 (N_10623,N_10459,N_10410);
nor U10624 (N_10624,N_10436,N_10355);
nand U10625 (N_10625,N_10403,N_10361);
nand U10626 (N_10626,N_10405,N_10357);
nor U10627 (N_10627,N_10459,N_10374);
and U10628 (N_10628,N_10430,N_10295);
and U10629 (N_10629,N_10437,N_10399);
nor U10630 (N_10630,N_10497,N_10413);
and U10631 (N_10631,N_10396,N_10373);
nand U10632 (N_10632,N_10420,N_10398);
and U10633 (N_10633,N_10402,N_10265);
or U10634 (N_10634,N_10325,N_10450);
nand U10635 (N_10635,N_10408,N_10434);
nand U10636 (N_10636,N_10325,N_10445);
nand U10637 (N_10637,N_10424,N_10494);
nand U10638 (N_10638,N_10426,N_10457);
nor U10639 (N_10639,N_10413,N_10313);
and U10640 (N_10640,N_10301,N_10360);
or U10641 (N_10641,N_10337,N_10403);
nor U10642 (N_10642,N_10337,N_10447);
or U10643 (N_10643,N_10347,N_10321);
and U10644 (N_10644,N_10417,N_10403);
xnor U10645 (N_10645,N_10310,N_10292);
or U10646 (N_10646,N_10270,N_10370);
or U10647 (N_10647,N_10295,N_10469);
and U10648 (N_10648,N_10349,N_10486);
and U10649 (N_10649,N_10470,N_10372);
and U10650 (N_10650,N_10478,N_10337);
or U10651 (N_10651,N_10413,N_10361);
or U10652 (N_10652,N_10445,N_10485);
nor U10653 (N_10653,N_10363,N_10414);
and U10654 (N_10654,N_10405,N_10350);
nor U10655 (N_10655,N_10337,N_10458);
and U10656 (N_10656,N_10310,N_10485);
nand U10657 (N_10657,N_10437,N_10484);
nand U10658 (N_10658,N_10440,N_10370);
and U10659 (N_10659,N_10259,N_10473);
nand U10660 (N_10660,N_10488,N_10304);
or U10661 (N_10661,N_10419,N_10332);
or U10662 (N_10662,N_10485,N_10386);
nand U10663 (N_10663,N_10366,N_10430);
xor U10664 (N_10664,N_10403,N_10312);
or U10665 (N_10665,N_10385,N_10251);
nor U10666 (N_10666,N_10251,N_10361);
nor U10667 (N_10667,N_10323,N_10472);
or U10668 (N_10668,N_10312,N_10353);
nor U10669 (N_10669,N_10316,N_10447);
or U10670 (N_10670,N_10367,N_10293);
nand U10671 (N_10671,N_10424,N_10293);
or U10672 (N_10672,N_10358,N_10471);
or U10673 (N_10673,N_10437,N_10456);
nand U10674 (N_10674,N_10298,N_10407);
nor U10675 (N_10675,N_10348,N_10309);
and U10676 (N_10676,N_10268,N_10446);
and U10677 (N_10677,N_10378,N_10358);
and U10678 (N_10678,N_10415,N_10348);
nand U10679 (N_10679,N_10312,N_10267);
nand U10680 (N_10680,N_10363,N_10312);
and U10681 (N_10681,N_10326,N_10421);
or U10682 (N_10682,N_10305,N_10443);
or U10683 (N_10683,N_10299,N_10438);
and U10684 (N_10684,N_10280,N_10290);
nand U10685 (N_10685,N_10315,N_10462);
nor U10686 (N_10686,N_10309,N_10294);
and U10687 (N_10687,N_10350,N_10353);
or U10688 (N_10688,N_10354,N_10287);
nor U10689 (N_10689,N_10338,N_10389);
xor U10690 (N_10690,N_10304,N_10463);
and U10691 (N_10691,N_10354,N_10495);
nand U10692 (N_10692,N_10278,N_10285);
nand U10693 (N_10693,N_10378,N_10380);
and U10694 (N_10694,N_10444,N_10469);
nor U10695 (N_10695,N_10405,N_10427);
nand U10696 (N_10696,N_10332,N_10327);
nand U10697 (N_10697,N_10422,N_10307);
and U10698 (N_10698,N_10484,N_10389);
or U10699 (N_10699,N_10352,N_10307);
nor U10700 (N_10700,N_10363,N_10424);
nor U10701 (N_10701,N_10328,N_10413);
or U10702 (N_10702,N_10315,N_10263);
and U10703 (N_10703,N_10412,N_10310);
or U10704 (N_10704,N_10302,N_10330);
or U10705 (N_10705,N_10416,N_10349);
nor U10706 (N_10706,N_10372,N_10495);
or U10707 (N_10707,N_10274,N_10377);
xnor U10708 (N_10708,N_10329,N_10497);
or U10709 (N_10709,N_10307,N_10496);
nor U10710 (N_10710,N_10267,N_10381);
or U10711 (N_10711,N_10458,N_10350);
nand U10712 (N_10712,N_10458,N_10296);
nor U10713 (N_10713,N_10448,N_10316);
nor U10714 (N_10714,N_10370,N_10472);
and U10715 (N_10715,N_10337,N_10476);
nor U10716 (N_10716,N_10425,N_10446);
nand U10717 (N_10717,N_10447,N_10311);
nor U10718 (N_10718,N_10390,N_10318);
nand U10719 (N_10719,N_10315,N_10312);
nor U10720 (N_10720,N_10297,N_10336);
and U10721 (N_10721,N_10411,N_10320);
or U10722 (N_10722,N_10398,N_10445);
nand U10723 (N_10723,N_10406,N_10377);
nor U10724 (N_10724,N_10394,N_10263);
or U10725 (N_10725,N_10429,N_10358);
nand U10726 (N_10726,N_10369,N_10352);
or U10727 (N_10727,N_10312,N_10388);
nor U10728 (N_10728,N_10298,N_10438);
nor U10729 (N_10729,N_10279,N_10371);
or U10730 (N_10730,N_10332,N_10335);
nor U10731 (N_10731,N_10496,N_10423);
or U10732 (N_10732,N_10438,N_10417);
nand U10733 (N_10733,N_10480,N_10289);
nor U10734 (N_10734,N_10323,N_10463);
nor U10735 (N_10735,N_10334,N_10317);
xnor U10736 (N_10736,N_10361,N_10261);
or U10737 (N_10737,N_10413,N_10289);
nor U10738 (N_10738,N_10318,N_10457);
nand U10739 (N_10739,N_10366,N_10450);
nand U10740 (N_10740,N_10398,N_10384);
and U10741 (N_10741,N_10487,N_10451);
or U10742 (N_10742,N_10406,N_10284);
or U10743 (N_10743,N_10390,N_10328);
nor U10744 (N_10744,N_10455,N_10256);
or U10745 (N_10745,N_10276,N_10370);
xnor U10746 (N_10746,N_10294,N_10348);
xor U10747 (N_10747,N_10412,N_10311);
nor U10748 (N_10748,N_10404,N_10299);
or U10749 (N_10749,N_10390,N_10388);
nand U10750 (N_10750,N_10697,N_10536);
or U10751 (N_10751,N_10515,N_10712);
and U10752 (N_10752,N_10699,N_10514);
nor U10753 (N_10753,N_10673,N_10695);
or U10754 (N_10754,N_10669,N_10604);
nand U10755 (N_10755,N_10560,N_10681);
nand U10756 (N_10756,N_10609,N_10539);
or U10757 (N_10757,N_10680,N_10580);
or U10758 (N_10758,N_10607,N_10729);
or U10759 (N_10759,N_10746,N_10717);
nand U10760 (N_10760,N_10525,N_10686);
and U10761 (N_10761,N_10524,N_10508);
or U10762 (N_10762,N_10630,N_10546);
nor U10763 (N_10763,N_10574,N_10690);
and U10764 (N_10764,N_10721,N_10594);
nand U10765 (N_10765,N_10613,N_10572);
nor U10766 (N_10766,N_10521,N_10741);
nor U10767 (N_10767,N_10679,N_10745);
and U10768 (N_10768,N_10675,N_10529);
nand U10769 (N_10769,N_10668,N_10674);
nand U10770 (N_10770,N_10735,N_10502);
xor U10771 (N_10771,N_10715,N_10626);
or U10772 (N_10772,N_10527,N_10654);
or U10773 (N_10773,N_10586,N_10561);
nor U10774 (N_10774,N_10567,N_10710);
nand U10775 (N_10775,N_10621,N_10707);
nand U10776 (N_10776,N_10510,N_10629);
or U10777 (N_10777,N_10584,N_10606);
nor U10778 (N_10778,N_10645,N_10543);
nor U10779 (N_10779,N_10672,N_10661);
nor U10780 (N_10780,N_10598,N_10682);
and U10781 (N_10781,N_10685,N_10605);
nand U10782 (N_10782,N_10612,N_10691);
nor U10783 (N_10783,N_10720,N_10702);
and U10784 (N_10784,N_10727,N_10549);
or U10785 (N_10785,N_10733,N_10581);
or U10786 (N_10786,N_10615,N_10601);
and U10787 (N_10787,N_10706,N_10670);
nor U10788 (N_10788,N_10575,N_10582);
nand U10789 (N_10789,N_10724,N_10624);
nand U10790 (N_10790,N_10657,N_10557);
nor U10791 (N_10791,N_10547,N_10569);
and U10792 (N_10792,N_10718,N_10506);
nor U10793 (N_10793,N_10659,N_10538);
and U10794 (N_10794,N_10507,N_10623);
and U10795 (N_10795,N_10653,N_10590);
and U10796 (N_10796,N_10622,N_10571);
and U10797 (N_10797,N_10503,N_10655);
nand U10798 (N_10798,N_10532,N_10748);
and U10799 (N_10799,N_10520,N_10534);
nand U10800 (N_10800,N_10732,N_10701);
nand U10801 (N_10801,N_10662,N_10704);
nor U10802 (N_10802,N_10716,N_10591);
or U10803 (N_10803,N_10518,N_10652);
and U10804 (N_10804,N_10592,N_10633);
and U10805 (N_10805,N_10738,N_10596);
and U10806 (N_10806,N_10658,N_10648);
or U10807 (N_10807,N_10568,N_10530);
nand U10808 (N_10808,N_10722,N_10696);
and U10809 (N_10809,N_10740,N_10577);
or U10810 (N_10810,N_10641,N_10540);
and U10811 (N_10811,N_10619,N_10734);
or U10812 (N_10812,N_10631,N_10589);
and U10813 (N_10813,N_10643,N_10709);
or U10814 (N_10814,N_10676,N_10666);
and U10815 (N_10815,N_10585,N_10742);
nand U10816 (N_10816,N_10556,N_10684);
nand U10817 (N_10817,N_10531,N_10526);
and U10818 (N_10818,N_10719,N_10550);
or U10819 (N_10819,N_10537,N_10744);
nand U10820 (N_10820,N_10555,N_10583);
nor U10821 (N_10821,N_10687,N_10700);
and U10822 (N_10822,N_10618,N_10714);
and U10823 (N_10823,N_10599,N_10627);
and U10824 (N_10824,N_10677,N_10647);
or U10825 (N_10825,N_10528,N_10671);
nor U10826 (N_10826,N_10642,N_10512);
or U10827 (N_10827,N_10500,N_10665);
nor U10828 (N_10828,N_10708,N_10663);
nor U10829 (N_10829,N_10644,N_10587);
and U10830 (N_10830,N_10638,N_10617);
or U10831 (N_10831,N_10650,N_10737);
nand U10832 (N_10832,N_10646,N_10743);
or U10833 (N_10833,N_10728,N_10573);
nor U10834 (N_10834,N_10632,N_10588);
and U10835 (N_10835,N_10640,N_10637);
nand U10836 (N_10836,N_10639,N_10542);
and U10837 (N_10837,N_10664,N_10552);
nand U10838 (N_10838,N_10509,N_10747);
nor U10839 (N_10839,N_10504,N_10563);
or U10840 (N_10840,N_10603,N_10614);
nor U10841 (N_10841,N_10636,N_10533);
nand U10842 (N_10842,N_10635,N_10656);
nor U10843 (N_10843,N_10620,N_10570);
nand U10844 (N_10844,N_10731,N_10564);
or U10845 (N_10845,N_10689,N_10544);
nor U10846 (N_10846,N_10725,N_10579);
or U10847 (N_10847,N_10595,N_10578);
or U10848 (N_10848,N_10616,N_10535);
nand U10849 (N_10849,N_10693,N_10730);
nor U10850 (N_10850,N_10501,N_10505);
and U10851 (N_10851,N_10694,N_10688);
nor U10852 (N_10852,N_10705,N_10559);
and U10853 (N_10853,N_10593,N_10523);
nand U10854 (N_10854,N_10713,N_10611);
or U10855 (N_10855,N_10522,N_10545);
or U10856 (N_10856,N_10692,N_10548);
nand U10857 (N_10857,N_10634,N_10554);
or U10858 (N_10858,N_10608,N_10565);
and U10859 (N_10859,N_10610,N_10553);
or U10860 (N_10860,N_10541,N_10703);
nand U10861 (N_10861,N_10511,N_10683);
or U10862 (N_10862,N_10516,N_10576);
nor U10863 (N_10863,N_10649,N_10562);
nand U10864 (N_10864,N_10711,N_10566);
nor U10865 (N_10865,N_10726,N_10597);
xnor U10866 (N_10866,N_10628,N_10739);
or U10867 (N_10867,N_10749,N_10517);
nor U10868 (N_10868,N_10736,N_10551);
nor U10869 (N_10869,N_10513,N_10625);
nand U10870 (N_10870,N_10602,N_10723);
nand U10871 (N_10871,N_10667,N_10698);
and U10872 (N_10872,N_10558,N_10678);
nand U10873 (N_10873,N_10660,N_10651);
nor U10874 (N_10874,N_10600,N_10519);
and U10875 (N_10875,N_10557,N_10706);
nand U10876 (N_10876,N_10741,N_10713);
or U10877 (N_10877,N_10621,N_10502);
or U10878 (N_10878,N_10552,N_10687);
nor U10879 (N_10879,N_10645,N_10676);
and U10880 (N_10880,N_10622,N_10505);
and U10881 (N_10881,N_10546,N_10553);
nand U10882 (N_10882,N_10610,N_10674);
or U10883 (N_10883,N_10505,N_10659);
nand U10884 (N_10884,N_10730,N_10739);
and U10885 (N_10885,N_10648,N_10503);
or U10886 (N_10886,N_10718,N_10606);
and U10887 (N_10887,N_10517,N_10608);
or U10888 (N_10888,N_10581,N_10569);
and U10889 (N_10889,N_10703,N_10741);
xnor U10890 (N_10890,N_10577,N_10552);
or U10891 (N_10891,N_10710,N_10680);
or U10892 (N_10892,N_10587,N_10661);
nor U10893 (N_10893,N_10542,N_10667);
nand U10894 (N_10894,N_10668,N_10552);
nand U10895 (N_10895,N_10553,N_10644);
nand U10896 (N_10896,N_10646,N_10533);
nand U10897 (N_10897,N_10638,N_10511);
or U10898 (N_10898,N_10562,N_10746);
nor U10899 (N_10899,N_10510,N_10543);
or U10900 (N_10900,N_10528,N_10644);
nand U10901 (N_10901,N_10716,N_10655);
and U10902 (N_10902,N_10607,N_10664);
nor U10903 (N_10903,N_10580,N_10558);
nor U10904 (N_10904,N_10589,N_10608);
and U10905 (N_10905,N_10670,N_10609);
and U10906 (N_10906,N_10744,N_10602);
nand U10907 (N_10907,N_10689,N_10570);
nor U10908 (N_10908,N_10649,N_10710);
nand U10909 (N_10909,N_10615,N_10504);
or U10910 (N_10910,N_10730,N_10628);
nand U10911 (N_10911,N_10540,N_10661);
or U10912 (N_10912,N_10745,N_10540);
or U10913 (N_10913,N_10621,N_10557);
or U10914 (N_10914,N_10732,N_10531);
nand U10915 (N_10915,N_10562,N_10518);
or U10916 (N_10916,N_10528,N_10533);
or U10917 (N_10917,N_10610,N_10587);
and U10918 (N_10918,N_10610,N_10649);
or U10919 (N_10919,N_10542,N_10676);
nand U10920 (N_10920,N_10633,N_10721);
nor U10921 (N_10921,N_10538,N_10519);
nand U10922 (N_10922,N_10600,N_10724);
or U10923 (N_10923,N_10574,N_10649);
xor U10924 (N_10924,N_10521,N_10616);
and U10925 (N_10925,N_10580,N_10623);
or U10926 (N_10926,N_10609,N_10656);
nor U10927 (N_10927,N_10551,N_10718);
nand U10928 (N_10928,N_10519,N_10691);
nand U10929 (N_10929,N_10679,N_10729);
and U10930 (N_10930,N_10550,N_10539);
or U10931 (N_10931,N_10709,N_10520);
and U10932 (N_10932,N_10620,N_10515);
nand U10933 (N_10933,N_10535,N_10573);
nor U10934 (N_10934,N_10550,N_10628);
and U10935 (N_10935,N_10666,N_10590);
and U10936 (N_10936,N_10575,N_10576);
nor U10937 (N_10937,N_10627,N_10681);
and U10938 (N_10938,N_10634,N_10557);
or U10939 (N_10939,N_10506,N_10542);
nand U10940 (N_10940,N_10567,N_10700);
nand U10941 (N_10941,N_10577,N_10684);
nor U10942 (N_10942,N_10583,N_10524);
nand U10943 (N_10943,N_10671,N_10511);
nand U10944 (N_10944,N_10647,N_10559);
or U10945 (N_10945,N_10568,N_10578);
or U10946 (N_10946,N_10578,N_10681);
or U10947 (N_10947,N_10512,N_10560);
and U10948 (N_10948,N_10567,N_10527);
and U10949 (N_10949,N_10576,N_10669);
or U10950 (N_10950,N_10551,N_10545);
or U10951 (N_10951,N_10590,N_10740);
and U10952 (N_10952,N_10619,N_10666);
or U10953 (N_10953,N_10676,N_10701);
and U10954 (N_10954,N_10500,N_10746);
nand U10955 (N_10955,N_10718,N_10588);
and U10956 (N_10956,N_10699,N_10635);
nor U10957 (N_10957,N_10685,N_10502);
nand U10958 (N_10958,N_10665,N_10686);
nor U10959 (N_10959,N_10526,N_10537);
and U10960 (N_10960,N_10744,N_10502);
nand U10961 (N_10961,N_10743,N_10536);
and U10962 (N_10962,N_10703,N_10567);
and U10963 (N_10963,N_10634,N_10617);
nor U10964 (N_10964,N_10598,N_10748);
or U10965 (N_10965,N_10634,N_10574);
or U10966 (N_10966,N_10717,N_10609);
and U10967 (N_10967,N_10689,N_10733);
or U10968 (N_10968,N_10624,N_10570);
and U10969 (N_10969,N_10628,N_10503);
or U10970 (N_10970,N_10702,N_10506);
nand U10971 (N_10971,N_10540,N_10615);
and U10972 (N_10972,N_10592,N_10730);
nand U10973 (N_10973,N_10579,N_10723);
or U10974 (N_10974,N_10555,N_10541);
or U10975 (N_10975,N_10691,N_10517);
nand U10976 (N_10976,N_10560,N_10735);
nor U10977 (N_10977,N_10647,N_10597);
and U10978 (N_10978,N_10640,N_10592);
nand U10979 (N_10979,N_10561,N_10533);
nor U10980 (N_10980,N_10649,N_10580);
nor U10981 (N_10981,N_10653,N_10655);
nand U10982 (N_10982,N_10685,N_10577);
xnor U10983 (N_10983,N_10652,N_10722);
nand U10984 (N_10984,N_10580,N_10614);
nand U10985 (N_10985,N_10748,N_10546);
nand U10986 (N_10986,N_10659,N_10655);
and U10987 (N_10987,N_10656,N_10555);
or U10988 (N_10988,N_10703,N_10715);
nor U10989 (N_10989,N_10722,N_10593);
nor U10990 (N_10990,N_10653,N_10571);
nand U10991 (N_10991,N_10732,N_10590);
or U10992 (N_10992,N_10745,N_10561);
nor U10993 (N_10993,N_10583,N_10599);
nor U10994 (N_10994,N_10744,N_10545);
nor U10995 (N_10995,N_10615,N_10621);
nand U10996 (N_10996,N_10537,N_10664);
or U10997 (N_10997,N_10619,N_10717);
or U10998 (N_10998,N_10714,N_10691);
nor U10999 (N_10999,N_10564,N_10732);
nor U11000 (N_11000,N_10920,N_10954);
nand U11001 (N_11001,N_10883,N_10816);
nor U11002 (N_11002,N_10995,N_10922);
nand U11003 (N_11003,N_10846,N_10787);
nor U11004 (N_11004,N_10933,N_10869);
and U11005 (N_11005,N_10784,N_10980);
or U11006 (N_11006,N_10976,N_10886);
or U11007 (N_11007,N_10911,N_10835);
and U11008 (N_11008,N_10944,N_10789);
nor U11009 (N_11009,N_10762,N_10998);
nand U11010 (N_11010,N_10760,N_10999);
or U11011 (N_11011,N_10982,N_10884);
nand U11012 (N_11012,N_10751,N_10934);
nand U11013 (N_11013,N_10874,N_10963);
nor U11014 (N_11014,N_10808,N_10904);
nand U11015 (N_11015,N_10773,N_10822);
nand U11016 (N_11016,N_10833,N_10788);
nand U11017 (N_11017,N_10810,N_10850);
nor U11018 (N_11018,N_10771,N_10818);
or U11019 (N_11019,N_10981,N_10813);
nor U11020 (N_11020,N_10928,N_10965);
and U11021 (N_11021,N_10791,N_10907);
or U11022 (N_11022,N_10798,N_10994);
and U11023 (N_11023,N_10848,N_10815);
nor U11024 (N_11024,N_10991,N_10940);
or U11025 (N_11025,N_10840,N_10962);
nand U11026 (N_11026,N_10875,N_10876);
or U11027 (N_11027,N_10975,N_10754);
nor U11028 (N_11028,N_10958,N_10780);
and U11029 (N_11029,N_10839,N_10892);
and U11030 (N_11030,N_10774,N_10864);
nand U11031 (N_11031,N_10782,N_10925);
and U11032 (N_11032,N_10937,N_10896);
and U11033 (N_11033,N_10821,N_10800);
xor U11034 (N_11034,N_10794,N_10842);
or U11035 (N_11035,N_10817,N_10942);
nand U11036 (N_11036,N_10814,N_10752);
and U11037 (N_11037,N_10777,N_10887);
or U11038 (N_11038,N_10870,N_10924);
nand U11039 (N_11039,N_10893,N_10895);
nand U11040 (N_11040,N_10804,N_10832);
xnor U11041 (N_11041,N_10843,N_10889);
nor U11042 (N_11042,N_10974,N_10831);
nand U11043 (N_11043,N_10823,N_10809);
or U11044 (N_11044,N_10903,N_10753);
nor U11045 (N_11045,N_10797,N_10756);
and U11046 (N_11046,N_10918,N_10837);
or U11047 (N_11047,N_10952,N_10897);
nor U11048 (N_11048,N_10939,N_10769);
and U11049 (N_11049,N_10770,N_10917);
or U11050 (N_11050,N_10880,N_10978);
and U11051 (N_11051,N_10992,N_10767);
nand U11052 (N_11052,N_10855,N_10763);
nor U11053 (N_11053,N_10901,N_10865);
or U11054 (N_11054,N_10863,N_10987);
nand U11055 (N_11055,N_10885,N_10970);
nand U11056 (N_11056,N_10931,N_10949);
nor U11057 (N_11057,N_10955,N_10946);
or U11058 (N_11058,N_10882,N_10766);
nand U11059 (N_11059,N_10851,N_10820);
or U11060 (N_11060,N_10775,N_10961);
and U11061 (N_11061,N_10972,N_10881);
and U11062 (N_11062,N_10929,N_10856);
and U11063 (N_11063,N_10902,N_10997);
or U11064 (N_11064,N_10805,N_10894);
nor U11065 (N_11065,N_10964,N_10926);
or U11066 (N_11066,N_10845,N_10802);
nor U11067 (N_11067,N_10830,N_10990);
and U11068 (N_11068,N_10758,N_10825);
nor U11069 (N_11069,N_10793,N_10861);
nor U11070 (N_11070,N_10910,N_10841);
or U11071 (N_11071,N_10913,N_10852);
and U11072 (N_11072,N_10899,N_10916);
and U11073 (N_11073,N_10966,N_10826);
nand U11074 (N_11074,N_10790,N_10945);
nand U11075 (N_11075,N_10948,N_10857);
and U11076 (N_11076,N_10783,N_10768);
xor U11077 (N_11077,N_10898,N_10941);
nand U11078 (N_11078,N_10827,N_10951);
or U11079 (N_11079,N_10776,N_10993);
nor U11080 (N_11080,N_10838,N_10960);
nand U11081 (N_11081,N_10973,N_10986);
nor U11082 (N_11082,N_10866,N_10824);
nand U11083 (N_11083,N_10905,N_10930);
nor U11084 (N_11084,N_10979,N_10750);
nand U11085 (N_11085,N_10936,N_10996);
nor U11086 (N_11086,N_10803,N_10847);
xor U11087 (N_11087,N_10854,N_10950);
nor U11088 (N_11088,N_10812,N_10761);
and U11089 (N_11089,N_10956,N_10877);
nor U11090 (N_11090,N_10988,N_10977);
nor U11091 (N_11091,N_10801,N_10935);
or U11092 (N_11092,N_10957,N_10890);
nand U11093 (N_11093,N_10891,N_10921);
and U11094 (N_11094,N_10836,N_10829);
or U11095 (N_11095,N_10888,N_10859);
nand U11096 (N_11096,N_10938,N_10873);
nand U11097 (N_11097,N_10959,N_10781);
and U11098 (N_11098,N_10858,N_10806);
nor U11099 (N_11099,N_10772,N_10853);
and U11100 (N_11100,N_10906,N_10984);
nand U11101 (N_11101,N_10778,N_10862);
xor U11102 (N_11102,N_10932,N_10878);
nand U11103 (N_11103,N_10755,N_10796);
or U11104 (N_11104,N_10792,N_10900);
and U11105 (N_11105,N_10844,N_10759);
nand U11106 (N_11106,N_10969,N_10968);
or U11107 (N_11107,N_10927,N_10860);
nor U11108 (N_11108,N_10879,N_10834);
and U11109 (N_11109,N_10867,N_10947);
or U11110 (N_11110,N_10908,N_10915);
nand U11111 (N_11111,N_10779,N_10765);
or U11112 (N_11112,N_10872,N_10807);
nand U11113 (N_11113,N_10799,N_10868);
nor U11114 (N_11114,N_10764,N_10811);
and U11115 (N_11115,N_10828,N_10795);
and U11116 (N_11116,N_10757,N_10983);
and U11117 (N_11117,N_10785,N_10914);
nand U11118 (N_11118,N_10871,N_10923);
xor U11119 (N_11119,N_10912,N_10967);
xnor U11120 (N_11120,N_10849,N_10943);
nor U11121 (N_11121,N_10971,N_10909);
and U11122 (N_11122,N_10989,N_10819);
or U11123 (N_11123,N_10985,N_10953);
or U11124 (N_11124,N_10919,N_10786);
and U11125 (N_11125,N_10824,N_10753);
nor U11126 (N_11126,N_10986,N_10808);
nand U11127 (N_11127,N_10923,N_10821);
or U11128 (N_11128,N_10956,N_10808);
or U11129 (N_11129,N_10978,N_10939);
or U11130 (N_11130,N_10875,N_10832);
or U11131 (N_11131,N_10956,N_10918);
or U11132 (N_11132,N_10959,N_10969);
nand U11133 (N_11133,N_10851,N_10843);
nand U11134 (N_11134,N_10962,N_10911);
nor U11135 (N_11135,N_10812,N_10764);
or U11136 (N_11136,N_10771,N_10793);
or U11137 (N_11137,N_10794,N_10880);
nor U11138 (N_11138,N_10957,N_10930);
and U11139 (N_11139,N_10801,N_10823);
nand U11140 (N_11140,N_10818,N_10895);
nor U11141 (N_11141,N_10763,N_10766);
nor U11142 (N_11142,N_10841,N_10925);
and U11143 (N_11143,N_10838,N_10781);
nor U11144 (N_11144,N_10788,N_10995);
nor U11145 (N_11145,N_10864,N_10957);
xor U11146 (N_11146,N_10986,N_10924);
or U11147 (N_11147,N_10840,N_10891);
xor U11148 (N_11148,N_10930,N_10945);
xnor U11149 (N_11149,N_10793,N_10754);
nand U11150 (N_11150,N_10882,N_10914);
or U11151 (N_11151,N_10882,N_10841);
and U11152 (N_11152,N_10834,N_10914);
nand U11153 (N_11153,N_10904,N_10754);
and U11154 (N_11154,N_10925,N_10822);
nand U11155 (N_11155,N_10997,N_10785);
or U11156 (N_11156,N_10926,N_10848);
and U11157 (N_11157,N_10761,N_10908);
nor U11158 (N_11158,N_10805,N_10788);
and U11159 (N_11159,N_10987,N_10865);
and U11160 (N_11160,N_10954,N_10841);
nand U11161 (N_11161,N_10999,N_10990);
or U11162 (N_11162,N_10755,N_10804);
nor U11163 (N_11163,N_10796,N_10957);
nor U11164 (N_11164,N_10896,N_10859);
nand U11165 (N_11165,N_10885,N_10809);
and U11166 (N_11166,N_10879,N_10796);
nand U11167 (N_11167,N_10841,N_10752);
or U11168 (N_11168,N_10860,N_10783);
nand U11169 (N_11169,N_10965,N_10870);
nand U11170 (N_11170,N_10961,N_10907);
nor U11171 (N_11171,N_10967,N_10924);
and U11172 (N_11172,N_10802,N_10864);
nor U11173 (N_11173,N_10756,N_10945);
nand U11174 (N_11174,N_10967,N_10805);
xor U11175 (N_11175,N_10922,N_10889);
and U11176 (N_11176,N_10951,N_10797);
and U11177 (N_11177,N_10994,N_10752);
nand U11178 (N_11178,N_10903,N_10823);
and U11179 (N_11179,N_10781,N_10753);
or U11180 (N_11180,N_10797,N_10900);
or U11181 (N_11181,N_10766,N_10965);
nand U11182 (N_11182,N_10797,N_10891);
nor U11183 (N_11183,N_10859,N_10823);
nand U11184 (N_11184,N_10849,N_10833);
or U11185 (N_11185,N_10938,N_10914);
and U11186 (N_11186,N_10959,N_10867);
or U11187 (N_11187,N_10783,N_10881);
and U11188 (N_11188,N_10804,N_10962);
and U11189 (N_11189,N_10933,N_10781);
nand U11190 (N_11190,N_10873,N_10760);
nand U11191 (N_11191,N_10878,N_10816);
nor U11192 (N_11192,N_10955,N_10962);
nand U11193 (N_11193,N_10756,N_10928);
nand U11194 (N_11194,N_10970,N_10818);
nand U11195 (N_11195,N_10986,N_10773);
nand U11196 (N_11196,N_10940,N_10863);
nand U11197 (N_11197,N_10974,N_10830);
nand U11198 (N_11198,N_10949,N_10789);
or U11199 (N_11199,N_10961,N_10881);
and U11200 (N_11200,N_10886,N_10771);
nor U11201 (N_11201,N_10944,N_10844);
or U11202 (N_11202,N_10802,N_10882);
and U11203 (N_11203,N_10910,N_10813);
and U11204 (N_11204,N_10939,N_10835);
and U11205 (N_11205,N_10852,N_10810);
or U11206 (N_11206,N_10942,N_10859);
and U11207 (N_11207,N_10959,N_10972);
and U11208 (N_11208,N_10759,N_10869);
nand U11209 (N_11209,N_10786,N_10966);
or U11210 (N_11210,N_10936,N_10805);
nor U11211 (N_11211,N_10780,N_10934);
or U11212 (N_11212,N_10892,N_10847);
nor U11213 (N_11213,N_10949,N_10919);
nor U11214 (N_11214,N_10942,N_10833);
and U11215 (N_11215,N_10760,N_10846);
xor U11216 (N_11216,N_10790,N_10924);
and U11217 (N_11217,N_10861,N_10816);
and U11218 (N_11218,N_10954,N_10940);
nor U11219 (N_11219,N_10906,N_10840);
and U11220 (N_11220,N_10919,N_10899);
or U11221 (N_11221,N_10782,N_10879);
nor U11222 (N_11222,N_10767,N_10828);
and U11223 (N_11223,N_10994,N_10933);
nor U11224 (N_11224,N_10890,N_10981);
nand U11225 (N_11225,N_10905,N_10801);
and U11226 (N_11226,N_10894,N_10785);
or U11227 (N_11227,N_10774,N_10798);
nand U11228 (N_11228,N_10801,N_10827);
or U11229 (N_11229,N_10970,N_10776);
nor U11230 (N_11230,N_10952,N_10862);
nor U11231 (N_11231,N_10766,N_10976);
or U11232 (N_11232,N_10905,N_10941);
and U11233 (N_11233,N_10802,N_10953);
nand U11234 (N_11234,N_10852,N_10934);
and U11235 (N_11235,N_10865,N_10859);
nand U11236 (N_11236,N_10836,N_10819);
nand U11237 (N_11237,N_10920,N_10874);
nor U11238 (N_11238,N_10898,N_10823);
and U11239 (N_11239,N_10883,N_10906);
nand U11240 (N_11240,N_10975,N_10962);
or U11241 (N_11241,N_10918,N_10794);
nor U11242 (N_11242,N_10842,N_10896);
nor U11243 (N_11243,N_10881,N_10939);
nor U11244 (N_11244,N_10764,N_10769);
nor U11245 (N_11245,N_10806,N_10928);
nand U11246 (N_11246,N_10874,N_10845);
or U11247 (N_11247,N_10879,N_10982);
nand U11248 (N_11248,N_10784,N_10900);
and U11249 (N_11249,N_10954,N_10893);
or U11250 (N_11250,N_11164,N_11219);
nand U11251 (N_11251,N_11237,N_11109);
nor U11252 (N_11252,N_11134,N_11000);
nor U11253 (N_11253,N_11046,N_11028);
nand U11254 (N_11254,N_11083,N_11146);
or U11255 (N_11255,N_11173,N_11159);
nor U11256 (N_11256,N_11176,N_11067);
and U11257 (N_11257,N_11100,N_11248);
and U11258 (N_11258,N_11025,N_11004);
xnor U11259 (N_11259,N_11145,N_11095);
and U11260 (N_11260,N_11072,N_11027);
nand U11261 (N_11261,N_11189,N_11065);
or U11262 (N_11262,N_11181,N_11130);
or U11263 (N_11263,N_11113,N_11114);
nand U11264 (N_11264,N_11023,N_11018);
or U11265 (N_11265,N_11049,N_11177);
xnor U11266 (N_11266,N_11220,N_11048);
and U11267 (N_11267,N_11239,N_11207);
and U11268 (N_11268,N_11240,N_11168);
and U11269 (N_11269,N_11151,N_11196);
or U11270 (N_11270,N_11226,N_11115);
and U11271 (N_11271,N_11017,N_11092);
nor U11272 (N_11272,N_11011,N_11052);
or U11273 (N_11273,N_11232,N_11241);
nor U11274 (N_11274,N_11131,N_11213);
and U11275 (N_11275,N_11169,N_11055);
nand U11276 (N_11276,N_11247,N_11203);
or U11277 (N_11277,N_11124,N_11099);
or U11278 (N_11278,N_11154,N_11063);
or U11279 (N_11279,N_11127,N_11167);
or U11280 (N_11280,N_11024,N_11102);
nand U11281 (N_11281,N_11197,N_11179);
and U11282 (N_11282,N_11142,N_11101);
nand U11283 (N_11283,N_11078,N_11013);
nand U11284 (N_11284,N_11026,N_11212);
or U11285 (N_11285,N_11079,N_11059);
and U11286 (N_11286,N_11006,N_11244);
or U11287 (N_11287,N_11035,N_11125);
nand U11288 (N_11288,N_11003,N_11221);
nand U11289 (N_11289,N_11193,N_11135);
nand U11290 (N_11290,N_11144,N_11227);
nand U11291 (N_11291,N_11238,N_11082);
or U11292 (N_11292,N_11016,N_11009);
and U11293 (N_11293,N_11061,N_11111);
nand U11294 (N_11294,N_11005,N_11186);
and U11295 (N_11295,N_11107,N_11235);
nand U11296 (N_11296,N_11037,N_11185);
or U11297 (N_11297,N_11056,N_11178);
nand U11298 (N_11298,N_11201,N_11075);
nor U11299 (N_11299,N_11209,N_11128);
and U11300 (N_11300,N_11138,N_11174);
nand U11301 (N_11301,N_11180,N_11084);
or U11302 (N_11302,N_11022,N_11170);
or U11303 (N_11303,N_11204,N_11153);
nor U11304 (N_11304,N_11215,N_11200);
nor U11305 (N_11305,N_11050,N_11105);
nor U11306 (N_11306,N_11042,N_11157);
nand U11307 (N_11307,N_11070,N_11136);
nor U11308 (N_11308,N_11191,N_11007);
or U11309 (N_11309,N_11031,N_11021);
and U11310 (N_11310,N_11195,N_11069);
nor U11311 (N_11311,N_11230,N_11122);
and U11312 (N_11312,N_11071,N_11015);
nor U11313 (N_11313,N_11019,N_11039);
and U11314 (N_11314,N_11162,N_11152);
nor U11315 (N_11315,N_11066,N_11234);
nand U11316 (N_11316,N_11184,N_11097);
and U11317 (N_11317,N_11202,N_11216);
nor U11318 (N_11318,N_11192,N_11121);
or U11319 (N_11319,N_11103,N_11057);
nor U11320 (N_11320,N_11141,N_11058);
nand U11321 (N_11321,N_11077,N_11206);
nand U11322 (N_11322,N_11233,N_11205);
and U11323 (N_11323,N_11047,N_11030);
and U11324 (N_11324,N_11041,N_11093);
or U11325 (N_11325,N_11229,N_11120);
nor U11326 (N_11326,N_11089,N_11171);
nor U11327 (N_11327,N_11053,N_11119);
nor U11328 (N_11328,N_11032,N_11150);
and U11329 (N_11329,N_11002,N_11094);
and U11330 (N_11330,N_11073,N_11236);
nor U11331 (N_11331,N_11137,N_11020);
or U11332 (N_11332,N_11012,N_11222);
nor U11333 (N_11333,N_11117,N_11051);
or U11334 (N_11334,N_11086,N_11108);
nand U11335 (N_11335,N_11225,N_11096);
or U11336 (N_11336,N_11064,N_11231);
nor U11337 (N_11337,N_11228,N_11104);
or U11338 (N_11338,N_11249,N_11029);
nor U11339 (N_11339,N_11098,N_11014);
nand U11340 (N_11340,N_11038,N_11218);
or U11341 (N_11341,N_11034,N_11044);
and U11342 (N_11342,N_11246,N_11198);
or U11343 (N_11343,N_11243,N_11139);
nand U11344 (N_11344,N_11123,N_11210);
nand U11345 (N_11345,N_11001,N_11074);
xor U11346 (N_11346,N_11081,N_11116);
nand U11347 (N_11347,N_11045,N_11126);
and U11348 (N_11348,N_11076,N_11158);
and U11349 (N_11349,N_11187,N_11091);
nor U11350 (N_11350,N_11208,N_11214);
nand U11351 (N_11351,N_11245,N_11165);
or U11352 (N_11352,N_11188,N_11175);
and U11353 (N_11353,N_11080,N_11132);
nor U11354 (N_11354,N_11163,N_11143);
and U11355 (N_11355,N_11043,N_11211);
xnor U11356 (N_11356,N_11161,N_11033);
or U11357 (N_11357,N_11068,N_11224);
and U11358 (N_11358,N_11190,N_11062);
and U11359 (N_11359,N_11112,N_11183);
nor U11360 (N_11360,N_11242,N_11129);
or U11361 (N_11361,N_11085,N_11133);
nor U11362 (N_11362,N_11054,N_11087);
or U11363 (N_11363,N_11155,N_11147);
nor U11364 (N_11364,N_11036,N_11149);
nand U11365 (N_11365,N_11110,N_11140);
and U11366 (N_11366,N_11160,N_11182);
and U11367 (N_11367,N_11156,N_11010);
nor U11368 (N_11368,N_11090,N_11217);
xnor U11369 (N_11369,N_11223,N_11060);
nand U11370 (N_11370,N_11106,N_11166);
nand U11371 (N_11371,N_11148,N_11172);
or U11372 (N_11372,N_11088,N_11199);
nor U11373 (N_11373,N_11194,N_11040);
nand U11374 (N_11374,N_11008,N_11118);
and U11375 (N_11375,N_11233,N_11241);
or U11376 (N_11376,N_11196,N_11180);
nand U11377 (N_11377,N_11005,N_11102);
nor U11378 (N_11378,N_11232,N_11212);
or U11379 (N_11379,N_11157,N_11206);
and U11380 (N_11380,N_11109,N_11039);
and U11381 (N_11381,N_11175,N_11148);
and U11382 (N_11382,N_11123,N_11206);
nand U11383 (N_11383,N_11009,N_11038);
nand U11384 (N_11384,N_11189,N_11164);
and U11385 (N_11385,N_11092,N_11170);
nand U11386 (N_11386,N_11244,N_11247);
nor U11387 (N_11387,N_11246,N_11241);
nand U11388 (N_11388,N_11234,N_11129);
nor U11389 (N_11389,N_11210,N_11060);
nor U11390 (N_11390,N_11086,N_11045);
or U11391 (N_11391,N_11190,N_11067);
and U11392 (N_11392,N_11190,N_11148);
nand U11393 (N_11393,N_11135,N_11112);
nor U11394 (N_11394,N_11242,N_11136);
nor U11395 (N_11395,N_11221,N_11103);
nand U11396 (N_11396,N_11123,N_11108);
nand U11397 (N_11397,N_11016,N_11025);
or U11398 (N_11398,N_11047,N_11143);
and U11399 (N_11399,N_11162,N_11205);
and U11400 (N_11400,N_11160,N_11178);
or U11401 (N_11401,N_11222,N_11153);
nand U11402 (N_11402,N_11167,N_11006);
and U11403 (N_11403,N_11238,N_11186);
nand U11404 (N_11404,N_11246,N_11210);
nand U11405 (N_11405,N_11089,N_11148);
nand U11406 (N_11406,N_11111,N_11190);
nor U11407 (N_11407,N_11211,N_11017);
nor U11408 (N_11408,N_11122,N_11149);
xnor U11409 (N_11409,N_11015,N_11064);
nor U11410 (N_11410,N_11211,N_11183);
or U11411 (N_11411,N_11005,N_11234);
and U11412 (N_11412,N_11070,N_11113);
and U11413 (N_11413,N_11000,N_11204);
nand U11414 (N_11414,N_11244,N_11115);
nand U11415 (N_11415,N_11222,N_11233);
and U11416 (N_11416,N_11244,N_11224);
and U11417 (N_11417,N_11217,N_11038);
and U11418 (N_11418,N_11217,N_11028);
nor U11419 (N_11419,N_11037,N_11076);
or U11420 (N_11420,N_11159,N_11146);
and U11421 (N_11421,N_11127,N_11159);
nor U11422 (N_11422,N_11005,N_11236);
nor U11423 (N_11423,N_11240,N_11178);
xor U11424 (N_11424,N_11128,N_11224);
nor U11425 (N_11425,N_11020,N_11095);
nor U11426 (N_11426,N_11111,N_11183);
nor U11427 (N_11427,N_11051,N_11099);
and U11428 (N_11428,N_11090,N_11197);
nand U11429 (N_11429,N_11219,N_11162);
and U11430 (N_11430,N_11142,N_11158);
nor U11431 (N_11431,N_11065,N_11191);
and U11432 (N_11432,N_11108,N_11187);
or U11433 (N_11433,N_11036,N_11071);
nor U11434 (N_11434,N_11247,N_11124);
nor U11435 (N_11435,N_11143,N_11224);
or U11436 (N_11436,N_11073,N_11150);
nor U11437 (N_11437,N_11131,N_11166);
or U11438 (N_11438,N_11216,N_11061);
nor U11439 (N_11439,N_11073,N_11061);
nand U11440 (N_11440,N_11201,N_11146);
and U11441 (N_11441,N_11203,N_11048);
nand U11442 (N_11442,N_11121,N_11037);
or U11443 (N_11443,N_11111,N_11238);
nor U11444 (N_11444,N_11227,N_11245);
xor U11445 (N_11445,N_11129,N_11211);
nand U11446 (N_11446,N_11113,N_11220);
and U11447 (N_11447,N_11141,N_11132);
nand U11448 (N_11448,N_11009,N_11197);
nor U11449 (N_11449,N_11081,N_11017);
or U11450 (N_11450,N_11211,N_11143);
nand U11451 (N_11451,N_11138,N_11171);
nor U11452 (N_11452,N_11153,N_11106);
or U11453 (N_11453,N_11024,N_11169);
nand U11454 (N_11454,N_11002,N_11013);
and U11455 (N_11455,N_11138,N_11137);
or U11456 (N_11456,N_11145,N_11122);
nor U11457 (N_11457,N_11159,N_11129);
and U11458 (N_11458,N_11108,N_11046);
or U11459 (N_11459,N_11021,N_11199);
or U11460 (N_11460,N_11049,N_11224);
or U11461 (N_11461,N_11022,N_11219);
and U11462 (N_11462,N_11229,N_11083);
and U11463 (N_11463,N_11071,N_11132);
or U11464 (N_11464,N_11090,N_11109);
or U11465 (N_11465,N_11020,N_11207);
and U11466 (N_11466,N_11007,N_11177);
or U11467 (N_11467,N_11059,N_11199);
and U11468 (N_11468,N_11095,N_11038);
nand U11469 (N_11469,N_11102,N_11018);
nor U11470 (N_11470,N_11153,N_11098);
or U11471 (N_11471,N_11117,N_11173);
nand U11472 (N_11472,N_11044,N_11051);
nand U11473 (N_11473,N_11204,N_11176);
xor U11474 (N_11474,N_11092,N_11105);
or U11475 (N_11475,N_11103,N_11211);
nor U11476 (N_11476,N_11046,N_11185);
or U11477 (N_11477,N_11214,N_11081);
xnor U11478 (N_11478,N_11218,N_11141);
nand U11479 (N_11479,N_11072,N_11246);
or U11480 (N_11480,N_11237,N_11162);
nor U11481 (N_11481,N_11121,N_11080);
or U11482 (N_11482,N_11005,N_11231);
nand U11483 (N_11483,N_11064,N_11118);
nor U11484 (N_11484,N_11050,N_11209);
nor U11485 (N_11485,N_11193,N_11147);
nand U11486 (N_11486,N_11107,N_11073);
nand U11487 (N_11487,N_11026,N_11220);
nor U11488 (N_11488,N_11076,N_11150);
nor U11489 (N_11489,N_11092,N_11143);
nor U11490 (N_11490,N_11057,N_11122);
nor U11491 (N_11491,N_11238,N_11061);
and U11492 (N_11492,N_11088,N_11077);
or U11493 (N_11493,N_11197,N_11055);
and U11494 (N_11494,N_11119,N_11246);
nor U11495 (N_11495,N_11070,N_11192);
nand U11496 (N_11496,N_11237,N_11160);
and U11497 (N_11497,N_11196,N_11176);
and U11498 (N_11498,N_11075,N_11241);
xnor U11499 (N_11499,N_11005,N_11043);
nor U11500 (N_11500,N_11463,N_11264);
and U11501 (N_11501,N_11442,N_11353);
or U11502 (N_11502,N_11411,N_11259);
nand U11503 (N_11503,N_11398,N_11298);
nand U11504 (N_11504,N_11446,N_11341);
nor U11505 (N_11505,N_11419,N_11410);
nor U11506 (N_11506,N_11409,N_11344);
or U11507 (N_11507,N_11488,N_11320);
or U11508 (N_11508,N_11273,N_11286);
or U11509 (N_11509,N_11389,N_11303);
nand U11510 (N_11510,N_11433,N_11301);
and U11511 (N_11511,N_11328,N_11417);
nand U11512 (N_11512,N_11289,N_11456);
nand U11513 (N_11513,N_11360,N_11477);
nor U11514 (N_11514,N_11429,N_11279);
and U11515 (N_11515,N_11432,N_11291);
nor U11516 (N_11516,N_11474,N_11428);
nand U11517 (N_11517,N_11375,N_11317);
or U11518 (N_11518,N_11471,N_11497);
nor U11519 (N_11519,N_11380,N_11307);
nand U11520 (N_11520,N_11420,N_11277);
nand U11521 (N_11521,N_11491,N_11422);
or U11522 (N_11522,N_11485,N_11283);
nand U11523 (N_11523,N_11470,N_11454);
xor U11524 (N_11524,N_11413,N_11486);
nand U11525 (N_11525,N_11408,N_11278);
or U11526 (N_11526,N_11430,N_11448);
nor U11527 (N_11527,N_11269,N_11451);
or U11528 (N_11528,N_11476,N_11299);
nand U11529 (N_11529,N_11316,N_11358);
and U11530 (N_11530,N_11350,N_11363);
or U11531 (N_11531,N_11333,N_11272);
nand U11532 (N_11532,N_11346,N_11386);
or U11533 (N_11533,N_11355,N_11250);
nor U11534 (N_11534,N_11458,N_11421);
nor U11535 (N_11535,N_11412,N_11462);
nand U11536 (N_11536,N_11426,N_11468);
nor U11537 (N_11537,N_11449,N_11452);
or U11538 (N_11538,N_11403,N_11295);
nor U11539 (N_11539,N_11304,N_11387);
and U11540 (N_11540,N_11359,N_11349);
and U11541 (N_11541,N_11388,N_11472);
nand U11542 (N_11542,N_11469,N_11483);
and U11543 (N_11543,N_11495,N_11435);
and U11544 (N_11544,N_11345,N_11414);
nor U11545 (N_11545,N_11496,N_11394);
nor U11546 (N_11546,N_11481,N_11268);
and U11547 (N_11547,N_11297,N_11261);
nand U11548 (N_11548,N_11276,N_11484);
nor U11549 (N_11549,N_11423,N_11447);
and U11550 (N_11550,N_11368,N_11364);
nand U11551 (N_11551,N_11251,N_11439);
or U11552 (N_11552,N_11302,N_11257);
nor U11553 (N_11553,N_11332,N_11356);
and U11554 (N_11554,N_11275,N_11313);
nor U11555 (N_11555,N_11370,N_11362);
nor U11556 (N_11556,N_11385,N_11253);
nand U11557 (N_11557,N_11287,N_11311);
nand U11558 (N_11558,N_11280,N_11334);
nand U11559 (N_11559,N_11494,N_11444);
nor U11560 (N_11560,N_11330,N_11336);
and U11561 (N_11561,N_11379,N_11402);
or U11562 (N_11562,N_11323,N_11397);
nand U11563 (N_11563,N_11418,N_11443);
or U11564 (N_11564,N_11445,N_11325);
or U11565 (N_11565,N_11427,N_11267);
nor U11566 (N_11566,N_11489,N_11399);
nor U11567 (N_11567,N_11318,N_11400);
nand U11568 (N_11568,N_11324,N_11347);
and U11569 (N_11569,N_11453,N_11461);
or U11570 (N_11570,N_11367,N_11366);
and U11571 (N_11571,N_11266,N_11331);
nand U11572 (N_11572,N_11436,N_11305);
or U11573 (N_11573,N_11308,N_11256);
nor U11574 (N_11574,N_11343,N_11378);
or U11575 (N_11575,N_11460,N_11450);
or U11576 (N_11576,N_11407,N_11437);
or U11577 (N_11577,N_11282,N_11425);
nand U11578 (N_11578,N_11376,N_11281);
nand U11579 (N_11579,N_11312,N_11296);
and U11580 (N_11580,N_11396,N_11498);
xor U11581 (N_11581,N_11487,N_11338);
nor U11582 (N_11582,N_11404,N_11479);
nand U11583 (N_11583,N_11288,N_11390);
or U11584 (N_11584,N_11357,N_11309);
nor U11585 (N_11585,N_11473,N_11383);
and U11586 (N_11586,N_11274,N_11406);
nand U11587 (N_11587,N_11441,N_11337);
nand U11588 (N_11588,N_11424,N_11361);
or U11589 (N_11589,N_11271,N_11292);
nand U11590 (N_11590,N_11365,N_11369);
and U11591 (N_11591,N_11340,N_11262);
and U11592 (N_11592,N_11265,N_11372);
and U11593 (N_11593,N_11405,N_11490);
or U11594 (N_11594,N_11499,N_11480);
or U11595 (N_11595,N_11381,N_11293);
and U11596 (N_11596,N_11377,N_11254);
nor U11597 (N_11597,N_11310,N_11354);
or U11598 (N_11598,N_11335,N_11457);
or U11599 (N_11599,N_11374,N_11314);
nor U11600 (N_11600,N_11326,N_11392);
nor U11601 (N_11601,N_11270,N_11467);
nor U11602 (N_11602,N_11464,N_11329);
and U11603 (N_11603,N_11416,N_11459);
xor U11604 (N_11604,N_11493,N_11351);
and U11605 (N_11605,N_11290,N_11255);
or U11606 (N_11606,N_11391,N_11492);
or U11607 (N_11607,N_11348,N_11306);
xnor U11608 (N_11608,N_11440,N_11319);
nor U11609 (N_11609,N_11401,N_11327);
and U11610 (N_11610,N_11322,N_11252);
and U11611 (N_11611,N_11434,N_11315);
and U11612 (N_11612,N_11258,N_11285);
nor U11613 (N_11613,N_11352,N_11339);
and U11614 (N_11614,N_11284,N_11415);
or U11615 (N_11615,N_11382,N_11300);
or U11616 (N_11616,N_11384,N_11431);
nand U11617 (N_11617,N_11466,N_11321);
nand U11618 (N_11618,N_11263,N_11455);
and U11619 (N_11619,N_11260,N_11482);
or U11620 (N_11620,N_11294,N_11393);
or U11621 (N_11621,N_11465,N_11373);
nor U11622 (N_11622,N_11438,N_11478);
or U11623 (N_11623,N_11371,N_11475);
nand U11624 (N_11624,N_11342,N_11395);
and U11625 (N_11625,N_11425,N_11350);
nor U11626 (N_11626,N_11464,N_11332);
nand U11627 (N_11627,N_11287,N_11345);
and U11628 (N_11628,N_11372,N_11301);
and U11629 (N_11629,N_11365,N_11286);
xnor U11630 (N_11630,N_11305,N_11402);
nor U11631 (N_11631,N_11425,N_11375);
and U11632 (N_11632,N_11446,N_11357);
and U11633 (N_11633,N_11493,N_11469);
nand U11634 (N_11634,N_11316,N_11267);
nor U11635 (N_11635,N_11274,N_11288);
nand U11636 (N_11636,N_11428,N_11253);
and U11637 (N_11637,N_11287,N_11423);
and U11638 (N_11638,N_11331,N_11258);
nor U11639 (N_11639,N_11363,N_11314);
or U11640 (N_11640,N_11431,N_11427);
nand U11641 (N_11641,N_11373,N_11420);
or U11642 (N_11642,N_11461,N_11437);
or U11643 (N_11643,N_11454,N_11469);
nor U11644 (N_11644,N_11255,N_11284);
and U11645 (N_11645,N_11454,N_11265);
or U11646 (N_11646,N_11283,N_11486);
or U11647 (N_11647,N_11363,N_11481);
or U11648 (N_11648,N_11316,N_11356);
or U11649 (N_11649,N_11383,N_11390);
nor U11650 (N_11650,N_11350,N_11354);
or U11651 (N_11651,N_11488,N_11468);
or U11652 (N_11652,N_11382,N_11444);
and U11653 (N_11653,N_11328,N_11299);
nand U11654 (N_11654,N_11353,N_11440);
nand U11655 (N_11655,N_11327,N_11488);
or U11656 (N_11656,N_11337,N_11335);
or U11657 (N_11657,N_11329,N_11375);
xor U11658 (N_11658,N_11395,N_11453);
and U11659 (N_11659,N_11429,N_11341);
nand U11660 (N_11660,N_11368,N_11270);
nand U11661 (N_11661,N_11429,N_11347);
nand U11662 (N_11662,N_11497,N_11359);
nor U11663 (N_11663,N_11391,N_11441);
xnor U11664 (N_11664,N_11360,N_11421);
or U11665 (N_11665,N_11418,N_11460);
and U11666 (N_11666,N_11311,N_11389);
nand U11667 (N_11667,N_11383,N_11259);
nand U11668 (N_11668,N_11443,N_11398);
nand U11669 (N_11669,N_11368,N_11414);
nor U11670 (N_11670,N_11443,N_11309);
nor U11671 (N_11671,N_11291,N_11498);
and U11672 (N_11672,N_11352,N_11488);
nand U11673 (N_11673,N_11410,N_11378);
or U11674 (N_11674,N_11485,N_11310);
nor U11675 (N_11675,N_11362,N_11347);
nand U11676 (N_11676,N_11318,N_11443);
and U11677 (N_11677,N_11256,N_11381);
or U11678 (N_11678,N_11457,N_11325);
or U11679 (N_11679,N_11289,N_11461);
nor U11680 (N_11680,N_11285,N_11292);
nor U11681 (N_11681,N_11373,N_11330);
nor U11682 (N_11682,N_11348,N_11290);
and U11683 (N_11683,N_11332,N_11486);
or U11684 (N_11684,N_11269,N_11323);
or U11685 (N_11685,N_11488,N_11370);
nor U11686 (N_11686,N_11353,N_11411);
nand U11687 (N_11687,N_11430,N_11369);
nor U11688 (N_11688,N_11414,N_11297);
or U11689 (N_11689,N_11399,N_11413);
xor U11690 (N_11690,N_11418,N_11424);
nor U11691 (N_11691,N_11315,N_11357);
and U11692 (N_11692,N_11369,N_11438);
nand U11693 (N_11693,N_11408,N_11272);
or U11694 (N_11694,N_11328,N_11289);
and U11695 (N_11695,N_11439,N_11457);
nand U11696 (N_11696,N_11448,N_11283);
nor U11697 (N_11697,N_11364,N_11328);
nor U11698 (N_11698,N_11432,N_11482);
xnor U11699 (N_11699,N_11432,N_11481);
or U11700 (N_11700,N_11419,N_11460);
and U11701 (N_11701,N_11497,N_11339);
nor U11702 (N_11702,N_11400,N_11275);
nand U11703 (N_11703,N_11465,N_11335);
and U11704 (N_11704,N_11360,N_11480);
nand U11705 (N_11705,N_11428,N_11490);
nor U11706 (N_11706,N_11460,N_11360);
nand U11707 (N_11707,N_11496,N_11303);
or U11708 (N_11708,N_11370,N_11394);
nor U11709 (N_11709,N_11427,N_11480);
and U11710 (N_11710,N_11273,N_11343);
or U11711 (N_11711,N_11332,N_11256);
nand U11712 (N_11712,N_11487,N_11493);
nand U11713 (N_11713,N_11418,N_11328);
and U11714 (N_11714,N_11447,N_11424);
nand U11715 (N_11715,N_11271,N_11354);
nor U11716 (N_11716,N_11323,N_11479);
nand U11717 (N_11717,N_11438,N_11263);
and U11718 (N_11718,N_11346,N_11319);
and U11719 (N_11719,N_11453,N_11427);
nand U11720 (N_11720,N_11498,N_11265);
nor U11721 (N_11721,N_11404,N_11326);
nand U11722 (N_11722,N_11293,N_11325);
nand U11723 (N_11723,N_11446,N_11494);
or U11724 (N_11724,N_11338,N_11495);
nand U11725 (N_11725,N_11252,N_11352);
nor U11726 (N_11726,N_11284,N_11346);
and U11727 (N_11727,N_11432,N_11333);
nand U11728 (N_11728,N_11425,N_11462);
nand U11729 (N_11729,N_11440,N_11410);
nand U11730 (N_11730,N_11274,N_11429);
or U11731 (N_11731,N_11317,N_11499);
nand U11732 (N_11732,N_11308,N_11464);
nor U11733 (N_11733,N_11250,N_11325);
nor U11734 (N_11734,N_11410,N_11358);
and U11735 (N_11735,N_11426,N_11278);
nand U11736 (N_11736,N_11475,N_11418);
and U11737 (N_11737,N_11275,N_11300);
nor U11738 (N_11738,N_11402,N_11324);
nand U11739 (N_11739,N_11465,N_11485);
or U11740 (N_11740,N_11382,N_11436);
nor U11741 (N_11741,N_11420,N_11425);
or U11742 (N_11742,N_11468,N_11342);
xor U11743 (N_11743,N_11472,N_11267);
nor U11744 (N_11744,N_11447,N_11279);
nand U11745 (N_11745,N_11421,N_11348);
or U11746 (N_11746,N_11408,N_11387);
or U11747 (N_11747,N_11357,N_11367);
nor U11748 (N_11748,N_11449,N_11318);
nand U11749 (N_11749,N_11333,N_11404);
and U11750 (N_11750,N_11669,N_11597);
xor U11751 (N_11751,N_11589,N_11728);
nand U11752 (N_11752,N_11749,N_11501);
and U11753 (N_11753,N_11559,N_11659);
or U11754 (N_11754,N_11718,N_11660);
xor U11755 (N_11755,N_11699,N_11617);
xnor U11756 (N_11756,N_11746,N_11735);
or U11757 (N_11757,N_11541,N_11712);
nand U11758 (N_11758,N_11637,N_11619);
and U11759 (N_11759,N_11590,N_11640);
or U11760 (N_11760,N_11638,N_11647);
and U11761 (N_11761,N_11503,N_11561);
nor U11762 (N_11762,N_11730,N_11719);
or U11763 (N_11763,N_11681,N_11573);
and U11764 (N_11764,N_11729,N_11510);
and U11765 (N_11765,N_11511,N_11635);
nand U11766 (N_11766,N_11701,N_11671);
nor U11767 (N_11767,N_11738,N_11650);
nor U11768 (N_11768,N_11717,N_11508);
or U11769 (N_11769,N_11734,N_11513);
and U11770 (N_11770,N_11506,N_11620);
and U11771 (N_11771,N_11535,N_11727);
or U11772 (N_11772,N_11581,N_11525);
nor U11773 (N_11773,N_11693,N_11615);
xnor U11774 (N_11774,N_11526,N_11556);
nor U11775 (N_11775,N_11592,N_11580);
or U11776 (N_11776,N_11545,N_11611);
nand U11777 (N_11777,N_11588,N_11628);
nand U11778 (N_11778,N_11532,N_11540);
and U11779 (N_11779,N_11686,N_11572);
or U11780 (N_11780,N_11586,N_11537);
nand U11781 (N_11781,N_11654,N_11582);
nand U11782 (N_11782,N_11575,N_11697);
nand U11783 (N_11783,N_11632,N_11737);
or U11784 (N_11784,N_11704,N_11722);
nor U11785 (N_11785,N_11715,N_11695);
nor U11786 (N_11786,N_11577,N_11550);
nor U11787 (N_11787,N_11595,N_11713);
or U11788 (N_11788,N_11744,N_11566);
and U11789 (N_11789,N_11736,N_11666);
or U11790 (N_11790,N_11564,N_11594);
nand U11791 (N_11791,N_11538,N_11684);
and U11792 (N_11792,N_11583,N_11683);
nor U11793 (N_11793,N_11720,N_11601);
nor U11794 (N_11794,N_11558,N_11618);
or U11795 (N_11795,N_11642,N_11740);
and U11796 (N_11796,N_11552,N_11731);
xnor U11797 (N_11797,N_11646,N_11672);
nor U11798 (N_11798,N_11578,N_11527);
or U11799 (N_11799,N_11544,N_11610);
nand U11800 (N_11800,N_11587,N_11733);
or U11801 (N_11801,N_11514,N_11613);
xnor U11802 (N_11802,N_11531,N_11745);
nand U11803 (N_11803,N_11591,N_11626);
or U11804 (N_11804,N_11534,N_11546);
or U11805 (N_11805,N_11656,N_11612);
or U11806 (N_11806,N_11702,N_11658);
and U11807 (N_11807,N_11533,N_11563);
nand U11808 (N_11808,N_11677,N_11609);
or U11809 (N_11809,N_11748,N_11623);
xnor U11810 (N_11810,N_11554,N_11521);
nor U11811 (N_11811,N_11690,N_11604);
or U11812 (N_11812,N_11674,N_11673);
and U11813 (N_11813,N_11689,N_11747);
nand U11814 (N_11814,N_11696,N_11543);
xnor U11815 (N_11815,N_11648,N_11668);
nor U11816 (N_11816,N_11678,N_11644);
and U11817 (N_11817,N_11553,N_11523);
nand U11818 (N_11818,N_11643,N_11520);
xor U11819 (N_11819,N_11622,N_11529);
nor U11820 (N_11820,N_11542,N_11562);
and U11821 (N_11821,N_11555,N_11725);
or U11822 (N_11822,N_11692,N_11518);
and U11823 (N_11823,N_11739,N_11710);
and U11824 (N_11824,N_11516,N_11680);
and U11825 (N_11825,N_11625,N_11574);
xor U11826 (N_11826,N_11726,N_11688);
nand U11827 (N_11827,N_11706,N_11585);
nor U11828 (N_11828,N_11652,N_11636);
nand U11829 (N_11829,N_11641,N_11627);
nand U11830 (N_11830,N_11530,N_11724);
and U11831 (N_11831,N_11662,N_11711);
and U11832 (N_11832,N_11676,N_11528);
or U11833 (N_11833,N_11603,N_11560);
nand U11834 (N_11834,N_11605,N_11505);
xor U11835 (N_11835,N_11682,N_11567);
or U11836 (N_11836,N_11517,N_11570);
nand U11837 (N_11837,N_11512,N_11721);
or U11838 (N_11838,N_11569,N_11741);
or U11839 (N_11839,N_11519,N_11515);
nor U11840 (N_11840,N_11700,N_11703);
nand U11841 (N_11841,N_11624,N_11629);
nand U11842 (N_11842,N_11565,N_11698);
or U11843 (N_11843,N_11548,N_11708);
and U11844 (N_11844,N_11653,N_11507);
and U11845 (N_11845,N_11657,N_11547);
nor U11846 (N_11846,N_11522,N_11716);
or U11847 (N_11847,N_11714,N_11705);
nor U11848 (N_11848,N_11549,N_11551);
and U11849 (N_11849,N_11502,N_11630);
nand U11850 (N_11850,N_11500,N_11707);
and U11851 (N_11851,N_11539,N_11557);
nand U11852 (N_11852,N_11599,N_11593);
or U11853 (N_11853,N_11742,N_11743);
and U11854 (N_11854,N_11723,N_11621);
nand U11855 (N_11855,N_11584,N_11649);
and U11856 (N_11856,N_11687,N_11600);
nor U11857 (N_11857,N_11607,N_11631);
and U11858 (N_11858,N_11651,N_11606);
or U11859 (N_11859,N_11655,N_11694);
nand U11860 (N_11860,N_11639,N_11670);
and U11861 (N_11861,N_11576,N_11664);
and U11862 (N_11862,N_11579,N_11633);
nor U11863 (N_11863,N_11602,N_11685);
and U11864 (N_11864,N_11504,N_11571);
or U11865 (N_11865,N_11661,N_11645);
and U11866 (N_11866,N_11524,N_11509);
or U11867 (N_11867,N_11536,N_11691);
nand U11868 (N_11868,N_11614,N_11665);
nor U11869 (N_11869,N_11634,N_11596);
nor U11870 (N_11870,N_11616,N_11732);
and U11871 (N_11871,N_11667,N_11709);
nand U11872 (N_11872,N_11663,N_11568);
or U11873 (N_11873,N_11598,N_11608);
nor U11874 (N_11874,N_11679,N_11675);
and U11875 (N_11875,N_11564,N_11537);
and U11876 (N_11876,N_11724,N_11615);
xor U11877 (N_11877,N_11539,N_11581);
and U11878 (N_11878,N_11605,N_11534);
and U11879 (N_11879,N_11726,N_11592);
or U11880 (N_11880,N_11581,N_11659);
nor U11881 (N_11881,N_11599,N_11509);
nor U11882 (N_11882,N_11516,N_11730);
and U11883 (N_11883,N_11746,N_11546);
and U11884 (N_11884,N_11622,N_11615);
nand U11885 (N_11885,N_11598,N_11678);
nand U11886 (N_11886,N_11621,N_11633);
or U11887 (N_11887,N_11547,N_11665);
nand U11888 (N_11888,N_11691,N_11697);
or U11889 (N_11889,N_11596,N_11707);
and U11890 (N_11890,N_11592,N_11568);
nand U11891 (N_11891,N_11637,N_11677);
or U11892 (N_11892,N_11523,N_11694);
nor U11893 (N_11893,N_11573,N_11571);
and U11894 (N_11894,N_11546,N_11701);
nand U11895 (N_11895,N_11618,N_11678);
or U11896 (N_11896,N_11523,N_11607);
or U11897 (N_11897,N_11609,N_11604);
or U11898 (N_11898,N_11714,N_11603);
and U11899 (N_11899,N_11575,N_11528);
and U11900 (N_11900,N_11725,N_11611);
or U11901 (N_11901,N_11714,N_11667);
nand U11902 (N_11902,N_11612,N_11565);
nand U11903 (N_11903,N_11679,N_11637);
and U11904 (N_11904,N_11657,N_11532);
nor U11905 (N_11905,N_11636,N_11539);
or U11906 (N_11906,N_11525,N_11600);
nor U11907 (N_11907,N_11534,N_11700);
and U11908 (N_11908,N_11621,N_11678);
or U11909 (N_11909,N_11540,N_11561);
and U11910 (N_11910,N_11725,N_11642);
nor U11911 (N_11911,N_11607,N_11656);
nor U11912 (N_11912,N_11711,N_11606);
nor U11913 (N_11913,N_11549,N_11662);
nor U11914 (N_11914,N_11609,N_11647);
nor U11915 (N_11915,N_11739,N_11565);
nor U11916 (N_11916,N_11713,N_11627);
nand U11917 (N_11917,N_11521,N_11705);
and U11918 (N_11918,N_11694,N_11699);
nand U11919 (N_11919,N_11683,N_11682);
nand U11920 (N_11920,N_11565,N_11509);
or U11921 (N_11921,N_11709,N_11572);
or U11922 (N_11922,N_11501,N_11643);
nand U11923 (N_11923,N_11693,N_11675);
nor U11924 (N_11924,N_11522,N_11642);
and U11925 (N_11925,N_11572,N_11714);
nor U11926 (N_11926,N_11658,N_11577);
nand U11927 (N_11927,N_11556,N_11638);
and U11928 (N_11928,N_11718,N_11720);
and U11929 (N_11929,N_11527,N_11688);
and U11930 (N_11930,N_11540,N_11718);
and U11931 (N_11931,N_11689,N_11502);
or U11932 (N_11932,N_11654,N_11509);
nor U11933 (N_11933,N_11737,N_11590);
and U11934 (N_11934,N_11732,N_11739);
or U11935 (N_11935,N_11742,N_11611);
and U11936 (N_11936,N_11578,N_11652);
and U11937 (N_11937,N_11724,N_11741);
and U11938 (N_11938,N_11743,N_11651);
nor U11939 (N_11939,N_11650,N_11529);
nand U11940 (N_11940,N_11528,N_11631);
and U11941 (N_11941,N_11525,N_11602);
nand U11942 (N_11942,N_11649,N_11736);
nand U11943 (N_11943,N_11588,N_11735);
and U11944 (N_11944,N_11536,N_11582);
nand U11945 (N_11945,N_11705,N_11533);
nor U11946 (N_11946,N_11530,N_11622);
nor U11947 (N_11947,N_11651,N_11608);
nand U11948 (N_11948,N_11684,N_11521);
xnor U11949 (N_11949,N_11560,N_11561);
and U11950 (N_11950,N_11553,N_11544);
nand U11951 (N_11951,N_11637,N_11564);
nand U11952 (N_11952,N_11565,N_11660);
nor U11953 (N_11953,N_11669,N_11706);
nor U11954 (N_11954,N_11731,N_11668);
and U11955 (N_11955,N_11574,N_11627);
nand U11956 (N_11956,N_11697,N_11627);
and U11957 (N_11957,N_11663,N_11545);
nor U11958 (N_11958,N_11626,N_11562);
nor U11959 (N_11959,N_11657,N_11631);
nand U11960 (N_11960,N_11724,N_11561);
nand U11961 (N_11961,N_11681,N_11519);
or U11962 (N_11962,N_11735,N_11601);
nor U11963 (N_11963,N_11567,N_11683);
and U11964 (N_11964,N_11644,N_11614);
xnor U11965 (N_11965,N_11727,N_11651);
or U11966 (N_11966,N_11518,N_11661);
or U11967 (N_11967,N_11509,N_11608);
xnor U11968 (N_11968,N_11587,N_11623);
and U11969 (N_11969,N_11683,N_11680);
and U11970 (N_11970,N_11720,N_11612);
and U11971 (N_11971,N_11583,N_11601);
and U11972 (N_11972,N_11586,N_11557);
nand U11973 (N_11973,N_11525,N_11509);
nor U11974 (N_11974,N_11679,N_11749);
nand U11975 (N_11975,N_11558,N_11641);
nand U11976 (N_11976,N_11655,N_11711);
nand U11977 (N_11977,N_11747,N_11589);
or U11978 (N_11978,N_11723,N_11609);
nor U11979 (N_11979,N_11589,N_11554);
and U11980 (N_11980,N_11690,N_11529);
and U11981 (N_11981,N_11745,N_11654);
or U11982 (N_11982,N_11715,N_11699);
and U11983 (N_11983,N_11739,N_11579);
nor U11984 (N_11984,N_11555,N_11500);
or U11985 (N_11985,N_11741,N_11559);
or U11986 (N_11986,N_11540,N_11557);
nor U11987 (N_11987,N_11593,N_11748);
nand U11988 (N_11988,N_11632,N_11661);
nor U11989 (N_11989,N_11668,N_11551);
nand U11990 (N_11990,N_11520,N_11521);
or U11991 (N_11991,N_11539,N_11524);
nor U11992 (N_11992,N_11620,N_11656);
nor U11993 (N_11993,N_11749,N_11618);
nor U11994 (N_11994,N_11530,N_11730);
and U11995 (N_11995,N_11615,N_11711);
or U11996 (N_11996,N_11644,N_11734);
or U11997 (N_11997,N_11677,N_11700);
nand U11998 (N_11998,N_11514,N_11645);
nand U11999 (N_11999,N_11687,N_11534);
nand U12000 (N_12000,N_11882,N_11889);
and U12001 (N_12001,N_11850,N_11910);
and U12002 (N_12002,N_11833,N_11950);
or U12003 (N_12003,N_11841,N_11798);
nor U12004 (N_12004,N_11951,N_11771);
nor U12005 (N_12005,N_11872,N_11812);
and U12006 (N_12006,N_11875,N_11917);
nand U12007 (N_12007,N_11813,N_11896);
and U12008 (N_12008,N_11905,N_11801);
xor U12009 (N_12009,N_11919,N_11756);
nor U12010 (N_12010,N_11851,N_11909);
or U12011 (N_12011,N_11804,N_11774);
nand U12012 (N_12012,N_11932,N_11878);
nor U12013 (N_12013,N_11754,N_11811);
nor U12014 (N_12014,N_11862,N_11855);
nor U12015 (N_12015,N_11758,N_11794);
nor U12016 (N_12016,N_11874,N_11877);
nor U12017 (N_12017,N_11777,N_11791);
or U12018 (N_12018,N_11834,N_11900);
and U12019 (N_12019,N_11803,N_11986);
and U12020 (N_12020,N_11787,N_11757);
and U12021 (N_12021,N_11987,N_11821);
nor U12022 (N_12022,N_11946,N_11890);
and U12023 (N_12023,N_11881,N_11956);
and U12024 (N_12024,N_11892,N_11810);
nor U12025 (N_12025,N_11886,N_11969);
and U12026 (N_12026,N_11891,N_11764);
nand U12027 (N_12027,N_11869,N_11830);
nand U12028 (N_12028,N_11785,N_11782);
or U12029 (N_12029,N_11924,N_11795);
and U12030 (N_12030,N_11867,N_11947);
nand U12031 (N_12031,N_11957,N_11888);
xor U12032 (N_12032,N_11752,N_11999);
and U12033 (N_12033,N_11974,N_11768);
nor U12034 (N_12034,N_11822,N_11995);
nand U12035 (N_12035,N_11854,N_11818);
nor U12036 (N_12036,N_11817,N_11927);
nor U12037 (N_12037,N_11808,N_11898);
nor U12038 (N_12038,N_11981,N_11860);
and U12039 (N_12039,N_11793,N_11997);
nand U12040 (N_12040,N_11998,N_11922);
nor U12041 (N_12041,N_11823,N_11784);
nand U12042 (N_12042,N_11959,N_11903);
and U12043 (N_12043,N_11937,N_11870);
or U12044 (N_12044,N_11883,N_11994);
xnor U12045 (N_12045,N_11968,N_11766);
nor U12046 (N_12046,N_11879,N_11781);
or U12047 (N_12047,N_11980,N_11966);
nand U12048 (N_12048,N_11928,N_11926);
nand U12049 (N_12049,N_11753,N_11831);
nor U12050 (N_12050,N_11836,N_11983);
nor U12051 (N_12051,N_11780,N_11972);
nor U12052 (N_12052,N_11975,N_11887);
nor U12053 (N_12053,N_11936,N_11770);
and U12054 (N_12054,N_11920,N_11802);
xor U12055 (N_12055,N_11827,N_11837);
or U12056 (N_12056,N_11824,N_11835);
or U12057 (N_12057,N_11904,N_11933);
nand U12058 (N_12058,N_11982,N_11943);
nand U12059 (N_12059,N_11805,N_11897);
nand U12060 (N_12060,N_11977,N_11952);
or U12061 (N_12061,N_11992,N_11846);
nor U12062 (N_12062,N_11852,N_11988);
nand U12063 (N_12063,N_11944,N_11884);
and U12064 (N_12064,N_11991,N_11894);
and U12065 (N_12065,N_11779,N_11790);
xnor U12066 (N_12066,N_11778,N_11913);
nor U12067 (N_12067,N_11847,N_11865);
nand U12068 (N_12068,N_11807,N_11767);
and U12069 (N_12069,N_11985,N_11989);
nor U12070 (N_12070,N_11792,N_11755);
nand U12071 (N_12071,N_11765,N_11921);
or U12072 (N_12072,N_11858,N_11799);
and U12073 (N_12073,N_11839,N_11819);
and U12074 (N_12074,N_11762,N_11911);
and U12075 (N_12075,N_11964,N_11930);
nor U12076 (N_12076,N_11857,N_11963);
nand U12077 (N_12077,N_11976,N_11797);
xor U12078 (N_12078,N_11861,N_11916);
nand U12079 (N_12079,N_11751,N_11843);
nand U12080 (N_12080,N_11901,N_11949);
nand U12081 (N_12081,N_11978,N_11816);
nand U12082 (N_12082,N_11825,N_11939);
nor U12083 (N_12083,N_11907,N_11772);
nor U12084 (N_12084,N_11853,N_11965);
or U12085 (N_12085,N_11942,N_11856);
or U12086 (N_12086,N_11828,N_11842);
and U12087 (N_12087,N_11786,N_11925);
nor U12088 (N_12088,N_11996,N_11938);
nor U12089 (N_12089,N_11769,N_11954);
nand U12090 (N_12090,N_11970,N_11893);
nor U12091 (N_12091,N_11962,N_11826);
nor U12092 (N_12092,N_11973,N_11960);
nor U12093 (N_12093,N_11760,N_11815);
or U12094 (N_12094,N_11908,N_11961);
nand U12095 (N_12095,N_11773,N_11829);
nor U12096 (N_12096,N_11871,N_11820);
nand U12097 (N_12097,N_11923,N_11906);
nand U12098 (N_12098,N_11912,N_11895);
nor U12099 (N_12099,N_11914,N_11832);
nand U12100 (N_12100,N_11955,N_11776);
and U12101 (N_12101,N_11848,N_11750);
nand U12102 (N_12102,N_11940,N_11806);
nand U12103 (N_12103,N_11880,N_11967);
and U12104 (N_12104,N_11866,N_11971);
or U12105 (N_12105,N_11931,N_11979);
or U12106 (N_12106,N_11761,N_11885);
nor U12107 (N_12107,N_11934,N_11876);
and U12108 (N_12108,N_11849,N_11941);
nor U12109 (N_12109,N_11800,N_11990);
and U12110 (N_12110,N_11873,N_11948);
nand U12111 (N_12111,N_11935,N_11863);
nor U12112 (N_12112,N_11840,N_11788);
nand U12113 (N_12113,N_11945,N_11868);
nand U12114 (N_12114,N_11789,N_11953);
or U12115 (N_12115,N_11864,N_11899);
nand U12116 (N_12116,N_11929,N_11775);
nor U12117 (N_12117,N_11838,N_11759);
or U12118 (N_12118,N_11918,N_11958);
or U12119 (N_12119,N_11915,N_11796);
nor U12120 (N_12120,N_11814,N_11809);
nand U12121 (N_12121,N_11859,N_11844);
or U12122 (N_12122,N_11763,N_11984);
and U12123 (N_12123,N_11783,N_11993);
and U12124 (N_12124,N_11902,N_11845);
nor U12125 (N_12125,N_11758,N_11754);
nand U12126 (N_12126,N_11793,N_11811);
and U12127 (N_12127,N_11851,N_11797);
nor U12128 (N_12128,N_11960,N_11783);
or U12129 (N_12129,N_11781,N_11932);
or U12130 (N_12130,N_11751,N_11787);
and U12131 (N_12131,N_11912,N_11836);
nand U12132 (N_12132,N_11918,N_11768);
nand U12133 (N_12133,N_11763,N_11791);
nand U12134 (N_12134,N_11856,N_11777);
nand U12135 (N_12135,N_11835,N_11750);
nand U12136 (N_12136,N_11878,N_11820);
or U12137 (N_12137,N_11867,N_11765);
nand U12138 (N_12138,N_11938,N_11861);
nor U12139 (N_12139,N_11961,N_11886);
or U12140 (N_12140,N_11941,N_11858);
nor U12141 (N_12141,N_11895,N_11816);
nand U12142 (N_12142,N_11808,N_11927);
nor U12143 (N_12143,N_11917,N_11979);
and U12144 (N_12144,N_11919,N_11957);
nor U12145 (N_12145,N_11935,N_11956);
nand U12146 (N_12146,N_11845,N_11888);
xor U12147 (N_12147,N_11799,N_11771);
and U12148 (N_12148,N_11976,N_11987);
nor U12149 (N_12149,N_11837,N_11903);
and U12150 (N_12150,N_11876,N_11955);
nand U12151 (N_12151,N_11756,N_11790);
nor U12152 (N_12152,N_11907,N_11828);
or U12153 (N_12153,N_11807,N_11859);
nand U12154 (N_12154,N_11960,N_11941);
and U12155 (N_12155,N_11942,N_11908);
nand U12156 (N_12156,N_11995,N_11867);
nor U12157 (N_12157,N_11992,N_11963);
and U12158 (N_12158,N_11881,N_11931);
and U12159 (N_12159,N_11971,N_11921);
or U12160 (N_12160,N_11877,N_11997);
or U12161 (N_12161,N_11840,N_11924);
nand U12162 (N_12162,N_11876,N_11907);
nand U12163 (N_12163,N_11860,N_11946);
nand U12164 (N_12164,N_11770,N_11872);
and U12165 (N_12165,N_11819,N_11939);
nor U12166 (N_12166,N_11859,N_11796);
or U12167 (N_12167,N_11881,N_11894);
or U12168 (N_12168,N_11806,N_11879);
nor U12169 (N_12169,N_11925,N_11843);
and U12170 (N_12170,N_11953,N_11753);
nand U12171 (N_12171,N_11987,N_11839);
nand U12172 (N_12172,N_11948,N_11766);
nor U12173 (N_12173,N_11987,N_11757);
and U12174 (N_12174,N_11842,N_11935);
and U12175 (N_12175,N_11765,N_11818);
and U12176 (N_12176,N_11846,N_11756);
or U12177 (N_12177,N_11937,N_11885);
nand U12178 (N_12178,N_11894,N_11846);
nand U12179 (N_12179,N_11911,N_11761);
or U12180 (N_12180,N_11888,N_11981);
nor U12181 (N_12181,N_11966,N_11772);
or U12182 (N_12182,N_11992,N_11943);
nand U12183 (N_12183,N_11809,N_11928);
or U12184 (N_12184,N_11960,N_11838);
and U12185 (N_12185,N_11901,N_11798);
nand U12186 (N_12186,N_11902,N_11936);
nor U12187 (N_12187,N_11912,N_11932);
nand U12188 (N_12188,N_11932,N_11977);
nor U12189 (N_12189,N_11873,N_11811);
or U12190 (N_12190,N_11886,N_11846);
nor U12191 (N_12191,N_11910,N_11774);
nor U12192 (N_12192,N_11811,N_11843);
and U12193 (N_12193,N_11784,N_11814);
or U12194 (N_12194,N_11815,N_11843);
nor U12195 (N_12195,N_11984,N_11831);
nand U12196 (N_12196,N_11876,N_11847);
or U12197 (N_12197,N_11964,N_11903);
or U12198 (N_12198,N_11764,N_11931);
nand U12199 (N_12199,N_11887,N_11967);
and U12200 (N_12200,N_11966,N_11890);
nand U12201 (N_12201,N_11994,N_11935);
and U12202 (N_12202,N_11955,N_11977);
and U12203 (N_12203,N_11991,N_11958);
nor U12204 (N_12204,N_11861,N_11885);
or U12205 (N_12205,N_11851,N_11940);
nor U12206 (N_12206,N_11873,N_11878);
xnor U12207 (N_12207,N_11910,N_11803);
or U12208 (N_12208,N_11848,N_11767);
and U12209 (N_12209,N_11831,N_11833);
nand U12210 (N_12210,N_11765,N_11770);
or U12211 (N_12211,N_11946,N_11789);
and U12212 (N_12212,N_11822,N_11823);
xor U12213 (N_12213,N_11861,N_11978);
and U12214 (N_12214,N_11961,N_11956);
and U12215 (N_12215,N_11894,N_11921);
nor U12216 (N_12216,N_11812,N_11927);
and U12217 (N_12217,N_11860,N_11877);
nor U12218 (N_12218,N_11919,N_11939);
and U12219 (N_12219,N_11750,N_11975);
and U12220 (N_12220,N_11897,N_11970);
nor U12221 (N_12221,N_11835,N_11931);
and U12222 (N_12222,N_11938,N_11869);
nor U12223 (N_12223,N_11833,N_11864);
xnor U12224 (N_12224,N_11763,N_11817);
xnor U12225 (N_12225,N_11756,N_11840);
or U12226 (N_12226,N_11994,N_11982);
nand U12227 (N_12227,N_11936,N_11764);
or U12228 (N_12228,N_11787,N_11777);
or U12229 (N_12229,N_11930,N_11801);
nor U12230 (N_12230,N_11964,N_11763);
and U12231 (N_12231,N_11944,N_11989);
or U12232 (N_12232,N_11812,N_11811);
and U12233 (N_12233,N_11852,N_11935);
and U12234 (N_12234,N_11971,N_11958);
nand U12235 (N_12235,N_11961,N_11968);
or U12236 (N_12236,N_11998,N_11971);
nand U12237 (N_12237,N_11923,N_11812);
nand U12238 (N_12238,N_11935,N_11907);
or U12239 (N_12239,N_11898,N_11995);
xor U12240 (N_12240,N_11751,N_11857);
nand U12241 (N_12241,N_11819,N_11856);
nor U12242 (N_12242,N_11914,N_11880);
and U12243 (N_12243,N_11832,N_11805);
nand U12244 (N_12244,N_11905,N_11815);
and U12245 (N_12245,N_11883,N_11904);
nand U12246 (N_12246,N_11782,N_11948);
and U12247 (N_12247,N_11942,N_11819);
or U12248 (N_12248,N_11908,N_11769);
nor U12249 (N_12249,N_11801,N_11781);
nand U12250 (N_12250,N_12015,N_12205);
and U12251 (N_12251,N_12013,N_12114);
nand U12252 (N_12252,N_12041,N_12115);
nor U12253 (N_12253,N_12188,N_12062);
xnor U12254 (N_12254,N_12142,N_12216);
nand U12255 (N_12255,N_12137,N_12133);
and U12256 (N_12256,N_12206,N_12161);
or U12257 (N_12257,N_12171,N_12162);
nor U12258 (N_12258,N_12042,N_12049);
nor U12259 (N_12259,N_12058,N_12066);
or U12260 (N_12260,N_12122,N_12201);
nor U12261 (N_12261,N_12138,N_12094);
and U12262 (N_12262,N_12127,N_12144);
or U12263 (N_12263,N_12173,N_12241);
nor U12264 (N_12264,N_12123,N_12223);
or U12265 (N_12265,N_12139,N_12184);
and U12266 (N_12266,N_12008,N_12072);
or U12267 (N_12267,N_12151,N_12101);
nor U12268 (N_12268,N_12028,N_12134);
nand U12269 (N_12269,N_12167,N_12045);
nor U12270 (N_12270,N_12048,N_12249);
nor U12271 (N_12271,N_12116,N_12248);
nand U12272 (N_12272,N_12197,N_12016);
and U12273 (N_12273,N_12177,N_12172);
and U12274 (N_12274,N_12017,N_12095);
nand U12275 (N_12275,N_12104,N_12176);
and U12276 (N_12276,N_12007,N_12166);
nand U12277 (N_12277,N_12090,N_12189);
or U12278 (N_12278,N_12237,N_12180);
nor U12279 (N_12279,N_12185,N_12059);
or U12280 (N_12280,N_12235,N_12165);
and U12281 (N_12281,N_12211,N_12202);
nor U12282 (N_12282,N_12034,N_12093);
and U12283 (N_12283,N_12074,N_12033);
or U12284 (N_12284,N_12175,N_12023);
or U12285 (N_12285,N_12082,N_12196);
or U12286 (N_12286,N_12024,N_12030);
nor U12287 (N_12287,N_12061,N_12052);
nand U12288 (N_12288,N_12010,N_12021);
and U12289 (N_12289,N_12079,N_12147);
nand U12290 (N_12290,N_12232,N_12131);
nand U12291 (N_12291,N_12207,N_12210);
nand U12292 (N_12292,N_12136,N_12113);
and U12293 (N_12293,N_12003,N_12157);
nor U12294 (N_12294,N_12190,N_12227);
or U12295 (N_12295,N_12078,N_12213);
or U12296 (N_12296,N_12009,N_12174);
and U12297 (N_12297,N_12056,N_12168);
nand U12298 (N_12298,N_12195,N_12199);
nor U12299 (N_12299,N_12051,N_12239);
or U12300 (N_12300,N_12043,N_12158);
nor U12301 (N_12301,N_12191,N_12014);
and U12302 (N_12302,N_12244,N_12055);
or U12303 (N_12303,N_12225,N_12182);
or U12304 (N_12304,N_12106,N_12245);
nor U12305 (N_12305,N_12057,N_12129);
nor U12306 (N_12306,N_12198,N_12154);
nor U12307 (N_12307,N_12040,N_12192);
or U12308 (N_12308,N_12083,N_12109);
and U12309 (N_12309,N_12152,N_12145);
nand U12310 (N_12310,N_12100,N_12118);
and U12311 (N_12311,N_12170,N_12080);
nand U12312 (N_12312,N_12230,N_12220);
nor U12313 (N_12313,N_12012,N_12046);
and U12314 (N_12314,N_12099,N_12200);
or U12315 (N_12315,N_12027,N_12037);
and U12316 (N_12316,N_12053,N_12224);
nor U12317 (N_12317,N_12087,N_12036);
nor U12318 (N_12318,N_12153,N_12086);
and U12319 (N_12319,N_12209,N_12143);
nor U12320 (N_12320,N_12039,N_12077);
nor U12321 (N_12321,N_12092,N_12035);
nor U12322 (N_12322,N_12060,N_12215);
or U12323 (N_12323,N_12005,N_12018);
nand U12324 (N_12324,N_12096,N_12064);
nand U12325 (N_12325,N_12219,N_12164);
or U12326 (N_12326,N_12070,N_12000);
nor U12327 (N_12327,N_12121,N_12022);
nor U12328 (N_12328,N_12098,N_12050);
nand U12329 (N_12329,N_12063,N_12125);
nand U12330 (N_12330,N_12214,N_12246);
or U12331 (N_12331,N_12120,N_12038);
or U12332 (N_12332,N_12044,N_12084);
nand U12333 (N_12333,N_12111,N_12004);
or U12334 (N_12334,N_12065,N_12132);
nor U12335 (N_12335,N_12141,N_12085);
nand U12336 (N_12336,N_12026,N_12054);
and U12337 (N_12337,N_12135,N_12238);
or U12338 (N_12338,N_12081,N_12217);
nand U12339 (N_12339,N_12240,N_12140);
or U12340 (N_12340,N_12218,N_12163);
nand U12341 (N_12341,N_12073,N_12148);
or U12342 (N_12342,N_12047,N_12117);
nor U12343 (N_12343,N_12102,N_12242);
or U12344 (N_12344,N_12181,N_12075);
or U12345 (N_12345,N_12108,N_12193);
nand U12346 (N_12346,N_12146,N_12029);
or U12347 (N_12347,N_12222,N_12091);
and U12348 (N_12348,N_12088,N_12001);
nand U12349 (N_12349,N_12179,N_12247);
and U12350 (N_12350,N_12208,N_12203);
and U12351 (N_12351,N_12126,N_12089);
nand U12352 (N_12352,N_12243,N_12149);
nor U12353 (N_12353,N_12226,N_12069);
nor U12354 (N_12354,N_12124,N_12032);
nor U12355 (N_12355,N_12020,N_12128);
nand U12356 (N_12356,N_12234,N_12186);
nor U12357 (N_12357,N_12228,N_12006);
nor U12358 (N_12358,N_12233,N_12105);
and U12359 (N_12359,N_12025,N_12130);
and U12360 (N_12360,N_12150,N_12221);
or U12361 (N_12361,N_12229,N_12067);
xnor U12362 (N_12362,N_12011,N_12236);
nand U12363 (N_12363,N_12160,N_12155);
nor U12364 (N_12364,N_12071,N_12169);
nor U12365 (N_12365,N_12194,N_12107);
nor U12366 (N_12366,N_12204,N_12002);
nand U12367 (N_12367,N_12231,N_12019);
and U12368 (N_12368,N_12119,N_12159);
and U12369 (N_12369,N_12076,N_12183);
and U12370 (N_12370,N_12112,N_12110);
or U12371 (N_12371,N_12178,N_12156);
nor U12372 (N_12372,N_12031,N_12097);
or U12373 (N_12373,N_12103,N_12187);
nand U12374 (N_12374,N_12212,N_12068);
nor U12375 (N_12375,N_12061,N_12100);
nor U12376 (N_12376,N_12110,N_12145);
and U12377 (N_12377,N_12068,N_12009);
or U12378 (N_12378,N_12205,N_12199);
nor U12379 (N_12379,N_12171,N_12161);
nand U12380 (N_12380,N_12146,N_12166);
nand U12381 (N_12381,N_12239,N_12123);
and U12382 (N_12382,N_12087,N_12181);
nand U12383 (N_12383,N_12083,N_12024);
nand U12384 (N_12384,N_12121,N_12224);
xor U12385 (N_12385,N_12249,N_12234);
or U12386 (N_12386,N_12003,N_12041);
or U12387 (N_12387,N_12181,N_12100);
and U12388 (N_12388,N_12132,N_12232);
nand U12389 (N_12389,N_12172,N_12144);
nand U12390 (N_12390,N_12027,N_12182);
nor U12391 (N_12391,N_12113,N_12092);
nor U12392 (N_12392,N_12155,N_12091);
nor U12393 (N_12393,N_12003,N_12113);
nor U12394 (N_12394,N_12080,N_12237);
xnor U12395 (N_12395,N_12186,N_12166);
and U12396 (N_12396,N_12058,N_12215);
or U12397 (N_12397,N_12084,N_12141);
and U12398 (N_12398,N_12177,N_12070);
nor U12399 (N_12399,N_12085,N_12144);
and U12400 (N_12400,N_12172,N_12233);
nor U12401 (N_12401,N_12019,N_12132);
and U12402 (N_12402,N_12189,N_12110);
nand U12403 (N_12403,N_12205,N_12125);
nand U12404 (N_12404,N_12128,N_12023);
and U12405 (N_12405,N_12069,N_12159);
nand U12406 (N_12406,N_12182,N_12099);
nand U12407 (N_12407,N_12187,N_12145);
xor U12408 (N_12408,N_12087,N_12219);
or U12409 (N_12409,N_12193,N_12117);
xnor U12410 (N_12410,N_12195,N_12158);
nand U12411 (N_12411,N_12132,N_12195);
or U12412 (N_12412,N_12023,N_12143);
nor U12413 (N_12413,N_12219,N_12055);
nor U12414 (N_12414,N_12140,N_12045);
nor U12415 (N_12415,N_12096,N_12137);
or U12416 (N_12416,N_12237,N_12000);
nand U12417 (N_12417,N_12006,N_12108);
nand U12418 (N_12418,N_12139,N_12213);
nand U12419 (N_12419,N_12208,N_12073);
or U12420 (N_12420,N_12164,N_12130);
nor U12421 (N_12421,N_12048,N_12164);
xnor U12422 (N_12422,N_12196,N_12038);
and U12423 (N_12423,N_12050,N_12007);
or U12424 (N_12424,N_12143,N_12211);
or U12425 (N_12425,N_12150,N_12068);
nand U12426 (N_12426,N_12008,N_12205);
and U12427 (N_12427,N_12020,N_12169);
nand U12428 (N_12428,N_12101,N_12210);
nor U12429 (N_12429,N_12015,N_12088);
or U12430 (N_12430,N_12042,N_12075);
or U12431 (N_12431,N_12222,N_12181);
xnor U12432 (N_12432,N_12117,N_12079);
or U12433 (N_12433,N_12123,N_12061);
and U12434 (N_12434,N_12088,N_12183);
nor U12435 (N_12435,N_12179,N_12229);
nor U12436 (N_12436,N_12228,N_12087);
xor U12437 (N_12437,N_12116,N_12182);
or U12438 (N_12438,N_12006,N_12038);
nor U12439 (N_12439,N_12017,N_12222);
or U12440 (N_12440,N_12088,N_12083);
nand U12441 (N_12441,N_12117,N_12054);
xor U12442 (N_12442,N_12238,N_12249);
nand U12443 (N_12443,N_12240,N_12234);
nor U12444 (N_12444,N_12101,N_12117);
and U12445 (N_12445,N_12002,N_12109);
nor U12446 (N_12446,N_12018,N_12155);
or U12447 (N_12447,N_12115,N_12121);
xor U12448 (N_12448,N_12082,N_12102);
or U12449 (N_12449,N_12111,N_12131);
nor U12450 (N_12450,N_12240,N_12243);
nand U12451 (N_12451,N_12014,N_12156);
nand U12452 (N_12452,N_12210,N_12238);
nand U12453 (N_12453,N_12158,N_12038);
and U12454 (N_12454,N_12071,N_12127);
nor U12455 (N_12455,N_12197,N_12022);
nand U12456 (N_12456,N_12247,N_12103);
nand U12457 (N_12457,N_12022,N_12072);
and U12458 (N_12458,N_12222,N_12225);
nor U12459 (N_12459,N_12158,N_12125);
nand U12460 (N_12460,N_12247,N_12052);
nand U12461 (N_12461,N_12232,N_12236);
and U12462 (N_12462,N_12104,N_12102);
nand U12463 (N_12463,N_12128,N_12150);
and U12464 (N_12464,N_12010,N_12055);
nand U12465 (N_12465,N_12239,N_12135);
and U12466 (N_12466,N_12153,N_12155);
or U12467 (N_12467,N_12100,N_12136);
nor U12468 (N_12468,N_12058,N_12232);
and U12469 (N_12469,N_12177,N_12065);
and U12470 (N_12470,N_12033,N_12067);
nor U12471 (N_12471,N_12123,N_12115);
or U12472 (N_12472,N_12220,N_12153);
nor U12473 (N_12473,N_12187,N_12000);
nor U12474 (N_12474,N_12087,N_12009);
or U12475 (N_12475,N_12140,N_12138);
and U12476 (N_12476,N_12081,N_12164);
nor U12477 (N_12477,N_12140,N_12113);
xnor U12478 (N_12478,N_12208,N_12011);
or U12479 (N_12479,N_12094,N_12092);
and U12480 (N_12480,N_12028,N_12205);
or U12481 (N_12481,N_12203,N_12108);
and U12482 (N_12482,N_12167,N_12015);
nand U12483 (N_12483,N_12198,N_12241);
and U12484 (N_12484,N_12018,N_12147);
nand U12485 (N_12485,N_12231,N_12217);
and U12486 (N_12486,N_12060,N_12167);
nand U12487 (N_12487,N_12034,N_12248);
nand U12488 (N_12488,N_12087,N_12224);
nor U12489 (N_12489,N_12094,N_12235);
nand U12490 (N_12490,N_12077,N_12081);
nand U12491 (N_12491,N_12249,N_12017);
nand U12492 (N_12492,N_12134,N_12196);
xnor U12493 (N_12493,N_12011,N_12104);
and U12494 (N_12494,N_12060,N_12242);
nand U12495 (N_12495,N_12063,N_12009);
or U12496 (N_12496,N_12136,N_12029);
nor U12497 (N_12497,N_12112,N_12070);
or U12498 (N_12498,N_12070,N_12037);
or U12499 (N_12499,N_12149,N_12086);
nand U12500 (N_12500,N_12276,N_12288);
nor U12501 (N_12501,N_12309,N_12263);
and U12502 (N_12502,N_12357,N_12268);
and U12503 (N_12503,N_12476,N_12397);
nor U12504 (N_12504,N_12256,N_12337);
nor U12505 (N_12505,N_12376,N_12449);
or U12506 (N_12506,N_12467,N_12374);
nand U12507 (N_12507,N_12336,N_12365);
nand U12508 (N_12508,N_12287,N_12345);
nand U12509 (N_12509,N_12342,N_12458);
and U12510 (N_12510,N_12391,N_12463);
nor U12511 (N_12511,N_12270,N_12335);
nor U12512 (N_12512,N_12412,N_12411);
or U12513 (N_12513,N_12447,N_12278);
nor U12514 (N_12514,N_12304,N_12427);
or U12515 (N_12515,N_12290,N_12407);
or U12516 (N_12516,N_12460,N_12487);
nand U12517 (N_12517,N_12349,N_12462);
nor U12518 (N_12518,N_12338,N_12355);
or U12519 (N_12519,N_12395,N_12421);
or U12520 (N_12520,N_12348,N_12334);
nor U12521 (N_12521,N_12394,N_12445);
nor U12522 (N_12522,N_12428,N_12405);
xor U12523 (N_12523,N_12398,N_12381);
nor U12524 (N_12524,N_12383,N_12451);
or U12525 (N_12525,N_12389,N_12300);
and U12526 (N_12526,N_12497,N_12436);
nor U12527 (N_12527,N_12302,N_12306);
and U12528 (N_12528,N_12344,N_12253);
or U12529 (N_12529,N_12354,N_12340);
nand U12530 (N_12530,N_12311,N_12316);
and U12531 (N_12531,N_12377,N_12274);
and U12532 (N_12532,N_12258,N_12281);
nor U12533 (N_12533,N_12275,N_12386);
nand U12534 (N_12534,N_12385,N_12390);
or U12535 (N_12535,N_12308,N_12474);
nor U12536 (N_12536,N_12489,N_12439);
xnor U12537 (N_12537,N_12272,N_12319);
nor U12538 (N_12538,N_12322,N_12314);
and U12539 (N_12539,N_12343,N_12438);
nor U12540 (N_12540,N_12452,N_12495);
nand U12541 (N_12541,N_12372,N_12317);
nor U12542 (N_12542,N_12339,N_12468);
or U12543 (N_12543,N_12415,N_12356);
nor U12544 (N_12544,N_12271,N_12273);
and U12545 (N_12545,N_12424,N_12472);
nand U12546 (N_12546,N_12291,N_12283);
or U12547 (N_12547,N_12353,N_12456);
nor U12548 (N_12548,N_12453,N_12384);
nand U12549 (N_12549,N_12437,N_12293);
and U12550 (N_12550,N_12418,N_12406);
and U12551 (N_12551,N_12260,N_12396);
nor U12552 (N_12552,N_12423,N_12368);
nor U12553 (N_12553,N_12426,N_12471);
or U12554 (N_12554,N_12446,N_12461);
and U12555 (N_12555,N_12475,N_12366);
nor U12556 (N_12556,N_12265,N_12433);
nand U12557 (N_12557,N_12465,N_12257);
nor U12558 (N_12558,N_12499,N_12332);
or U12559 (N_12559,N_12483,N_12251);
and U12560 (N_12560,N_12402,N_12358);
or U12561 (N_12561,N_12488,N_12303);
nor U12562 (N_12562,N_12417,N_12359);
and U12563 (N_12563,N_12444,N_12387);
or U12564 (N_12564,N_12413,N_12295);
nand U12565 (N_12565,N_12410,N_12482);
or U12566 (N_12566,N_12312,N_12364);
nand U12567 (N_12567,N_12380,N_12481);
or U12568 (N_12568,N_12261,N_12455);
and U12569 (N_12569,N_12414,N_12379);
xnor U12570 (N_12570,N_12297,N_12484);
and U12571 (N_12571,N_12425,N_12360);
nor U12572 (N_12572,N_12370,N_12315);
and U12573 (N_12573,N_12459,N_12473);
nand U12574 (N_12574,N_12255,N_12400);
nor U12575 (N_12575,N_12301,N_12313);
nand U12576 (N_12576,N_12352,N_12375);
and U12577 (N_12577,N_12250,N_12448);
and U12578 (N_12578,N_12430,N_12404);
or U12579 (N_12579,N_12254,N_12470);
nand U12580 (N_12580,N_12399,N_12477);
nand U12581 (N_12581,N_12422,N_12442);
xor U12582 (N_12582,N_12351,N_12259);
or U12583 (N_12583,N_12331,N_12333);
nor U12584 (N_12584,N_12420,N_12269);
nand U12585 (N_12585,N_12371,N_12419);
or U12586 (N_12586,N_12267,N_12443);
nand U12587 (N_12587,N_12491,N_12252);
nor U12588 (N_12588,N_12327,N_12494);
or U12589 (N_12589,N_12480,N_12431);
and U12590 (N_12590,N_12279,N_12321);
or U12591 (N_12591,N_12378,N_12266);
or U12592 (N_12592,N_12289,N_12329);
nand U12593 (N_12593,N_12429,N_12496);
nor U12594 (N_12594,N_12292,N_12296);
nand U12595 (N_12595,N_12490,N_12294);
nand U12596 (N_12596,N_12485,N_12280);
xnor U12597 (N_12597,N_12416,N_12388);
and U12598 (N_12598,N_12284,N_12367);
and U12599 (N_12599,N_12305,N_12408);
nand U12600 (N_12600,N_12454,N_12307);
nand U12601 (N_12601,N_12493,N_12285);
or U12602 (N_12602,N_12324,N_12286);
and U12603 (N_12603,N_12298,N_12326);
or U12604 (N_12604,N_12478,N_12403);
nor U12605 (N_12605,N_12361,N_12435);
or U12606 (N_12606,N_12457,N_12264);
and U12607 (N_12607,N_12369,N_12393);
nor U12608 (N_12608,N_12320,N_12401);
and U12609 (N_12609,N_12347,N_12362);
or U12610 (N_12610,N_12450,N_12310);
nand U12611 (N_12611,N_12299,N_12328);
nand U12612 (N_12612,N_12277,N_12486);
xor U12613 (N_12613,N_12492,N_12382);
or U12614 (N_12614,N_12441,N_12469);
or U12615 (N_12615,N_12330,N_12464);
xnor U12616 (N_12616,N_12440,N_12346);
or U12617 (N_12617,N_12498,N_12341);
nand U12618 (N_12618,N_12282,N_12350);
or U12619 (N_12619,N_12262,N_12373);
nor U12620 (N_12620,N_12434,N_12479);
or U12621 (N_12621,N_12466,N_12318);
or U12622 (N_12622,N_12325,N_12392);
nand U12623 (N_12623,N_12409,N_12363);
or U12624 (N_12624,N_12432,N_12323);
and U12625 (N_12625,N_12443,N_12379);
nand U12626 (N_12626,N_12413,N_12372);
and U12627 (N_12627,N_12279,N_12319);
or U12628 (N_12628,N_12318,N_12341);
nor U12629 (N_12629,N_12257,N_12390);
nor U12630 (N_12630,N_12378,N_12260);
nand U12631 (N_12631,N_12364,N_12264);
or U12632 (N_12632,N_12435,N_12307);
nor U12633 (N_12633,N_12372,N_12442);
nor U12634 (N_12634,N_12430,N_12379);
and U12635 (N_12635,N_12321,N_12317);
nor U12636 (N_12636,N_12326,N_12478);
and U12637 (N_12637,N_12320,N_12455);
and U12638 (N_12638,N_12324,N_12461);
or U12639 (N_12639,N_12478,N_12459);
nor U12640 (N_12640,N_12373,N_12293);
nand U12641 (N_12641,N_12275,N_12313);
or U12642 (N_12642,N_12298,N_12478);
and U12643 (N_12643,N_12316,N_12487);
nor U12644 (N_12644,N_12268,N_12499);
or U12645 (N_12645,N_12492,N_12298);
or U12646 (N_12646,N_12373,N_12362);
nand U12647 (N_12647,N_12278,N_12412);
nand U12648 (N_12648,N_12286,N_12276);
and U12649 (N_12649,N_12273,N_12384);
or U12650 (N_12650,N_12457,N_12383);
nand U12651 (N_12651,N_12350,N_12354);
and U12652 (N_12652,N_12394,N_12482);
nor U12653 (N_12653,N_12334,N_12343);
xnor U12654 (N_12654,N_12403,N_12291);
nand U12655 (N_12655,N_12476,N_12329);
or U12656 (N_12656,N_12392,N_12472);
nor U12657 (N_12657,N_12425,N_12460);
and U12658 (N_12658,N_12481,N_12334);
or U12659 (N_12659,N_12384,N_12361);
and U12660 (N_12660,N_12356,N_12464);
nand U12661 (N_12661,N_12263,N_12267);
nor U12662 (N_12662,N_12448,N_12479);
nor U12663 (N_12663,N_12428,N_12415);
nor U12664 (N_12664,N_12415,N_12388);
nor U12665 (N_12665,N_12281,N_12392);
xnor U12666 (N_12666,N_12429,N_12370);
and U12667 (N_12667,N_12434,N_12395);
or U12668 (N_12668,N_12446,N_12327);
or U12669 (N_12669,N_12296,N_12415);
nor U12670 (N_12670,N_12453,N_12444);
nand U12671 (N_12671,N_12414,N_12428);
or U12672 (N_12672,N_12459,N_12335);
or U12673 (N_12673,N_12308,N_12303);
nand U12674 (N_12674,N_12392,N_12380);
or U12675 (N_12675,N_12267,N_12353);
nand U12676 (N_12676,N_12448,N_12441);
nor U12677 (N_12677,N_12439,N_12267);
and U12678 (N_12678,N_12452,N_12387);
nor U12679 (N_12679,N_12364,N_12347);
nand U12680 (N_12680,N_12404,N_12282);
or U12681 (N_12681,N_12316,N_12321);
or U12682 (N_12682,N_12272,N_12424);
and U12683 (N_12683,N_12416,N_12404);
or U12684 (N_12684,N_12263,N_12460);
nor U12685 (N_12685,N_12348,N_12338);
or U12686 (N_12686,N_12405,N_12488);
or U12687 (N_12687,N_12269,N_12377);
nor U12688 (N_12688,N_12471,N_12372);
nor U12689 (N_12689,N_12317,N_12363);
and U12690 (N_12690,N_12266,N_12398);
and U12691 (N_12691,N_12363,N_12353);
and U12692 (N_12692,N_12416,N_12413);
nor U12693 (N_12693,N_12331,N_12261);
xor U12694 (N_12694,N_12400,N_12468);
nor U12695 (N_12695,N_12257,N_12400);
nand U12696 (N_12696,N_12343,N_12313);
or U12697 (N_12697,N_12471,N_12368);
nor U12698 (N_12698,N_12286,N_12291);
nand U12699 (N_12699,N_12251,N_12484);
or U12700 (N_12700,N_12388,N_12490);
and U12701 (N_12701,N_12308,N_12371);
nand U12702 (N_12702,N_12403,N_12445);
nor U12703 (N_12703,N_12359,N_12406);
and U12704 (N_12704,N_12323,N_12322);
and U12705 (N_12705,N_12407,N_12402);
nand U12706 (N_12706,N_12316,N_12484);
or U12707 (N_12707,N_12485,N_12302);
and U12708 (N_12708,N_12386,N_12321);
xor U12709 (N_12709,N_12436,N_12320);
or U12710 (N_12710,N_12335,N_12287);
and U12711 (N_12711,N_12261,N_12430);
nor U12712 (N_12712,N_12281,N_12453);
nor U12713 (N_12713,N_12278,N_12259);
and U12714 (N_12714,N_12340,N_12473);
nand U12715 (N_12715,N_12328,N_12349);
nand U12716 (N_12716,N_12454,N_12475);
nor U12717 (N_12717,N_12369,N_12485);
xor U12718 (N_12718,N_12477,N_12359);
or U12719 (N_12719,N_12396,N_12410);
and U12720 (N_12720,N_12432,N_12393);
or U12721 (N_12721,N_12403,N_12298);
xor U12722 (N_12722,N_12452,N_12476);
nor U12723 (N_12723,N_12399,N_12346);
nor U12724 (N_12724,N_12290,N_12392);
nand U12725 (N_12725,N_12497,N_12336);
nor U12726 (N_12726,N_12342,N_12373);
nor U12727 (N_12727,N_12448,N_12415);
nand U12728 (N_12728,N_12388,N_12484);
nor U12729 (N_12729,N_12458,N_12422);
or U12730 (N_12730,N_12399,N_12374);
nor U12731 (N_12731,N_12406,N_12379);
and U12732 (N_12732,N_12396,N_12493);
or U12733 (N_12733,N_12363,N_12300);
nor U12734 (N_12734,N_12467,N_12379);
nand U12735 (N_12735,N_12252,N_12447);
nand U12736 (N_12736,N_12284,N_12307);
nand U12737 (N_12737,N_12459,N_12451);
nand U12738 (N_12738,N_12489,N_12393);
nand U12739 (N_12739,N_12328,N_12309);
or U12740 (N_12740,N_12276,N_12492);
or U12741 (N_12741,N_12490,N_12352);
nor U12742 (N_12742,N_12277,N_12396);
nand U12743 (N_12743,N_12436,N_12348);
nand U12744 (N_12744,N_12389,N_12283);
or U12745 (N_12745,N_12258,N_12429);
nand U12746 (N_12746,N_12358,N_12332);
nor U12747 (N_12747,N_12353,N_12498);
nor U12748 (N_12748,N_12391,N_12322);
and U12749 (N_12749,N_12321,N_12270);
nand U12750 (N_12750,N_12536,N_12507);
nor U12751 (N_12751,N_12623,N_12561);
and U12752 (N_12752,N_12527,N_12668);
or U12753 (N_12753,N_12639,N_12608);
nand U12754 (N_12754,N_12506,N_12731);
or U12755 (N_12755,N_12620,N_12563);
or U12756 (N_12756,N_12571,N_12710);
or U12757 (N_12757,N_12733,N_12663);
and U12758 (N_12758,N_12607,N_12677);
xnor U12759 (N_12759,N_12640,N_12535);
and U12760 (N_12760,N_12554,N_12503);
and U12761 (N_12761,N_12655,N_12558);
nand U12762 (N_12762,N_12517,N_12728);
and U12763 (N_12763,N_12635,N_12642);
nor U12764 (N_12764,N_12701,N_12675);
nand U12765 (N_12765,N_12511,N_12567);
nand U12766 (N_12766,N_12590,N_12665);
and U12767 (N_12767,N_12593,N_12707);
and U12768 (N_12768,N_12589,N_12723);
nand U12769 (N_12769,N_12541,N_12621);
and U12770 (N_12770,N_12553,N_12513);
nor U12771 (N_12771,N_12574,N_12572);
or U12772 (N_12772,N_12534,N_12587);
and U12773 (N_12773,N_12697,N_12520);
and U12774 (N_12774,N_12595,N_12573);
nor U12775 (N_12775,N_12652,N_12649);
and U12776 (N_12776,N_12727,N_12551);
or U12777 (N_12777,N_12521,N_12526);
or U12778 (N_12778,N_12687,N_12606);
nand U12779 (N_12779,N_12648,N_12523);
or U12780 (N_12780,N_12748,N_12596);
and U12781 (N_12781,N_12634,N_12700);
and U12782 (N_12782,N_12709,N_12694);
nand U12783 (N_12783,N_12721,N_12614);
or U12784 (N_12784,N_12547,N_12657);
nand U12785 (N_12785,N_12539,N_12550);
and U12786 (N_12786,N_12653,N_12586);
or U12787 (N_12787,N_12680,N_12722);
or U12788 (N_12788,N_12669,N_12712);
and U12789 (N_12789,N_12603,N_12515);
nand U12790 (N_12790,N_12670,N_12662);
nand U12791 (N_12791,N_12568,N_12514);
nand U12792 (N_12792,N_12556,N_12601);
and U12793 (N_12793,N_12602,N_12691);
nor U12794 (N_12794,N_12674,N_12559);
or U12795 (N_12795,N_12647,N_12509);
nand U12796 (N_12796,N_12616,N_12717);
and U12797 (N_12797,N_12718,N_12693);
or U12798 (N_12798,N_12531,N_12549);
and U12799 (N_12799,N_12598,N_12711);
and U12800 (N_12800,N_12505,N_12622);
nor U12801 (N_12801,N_12726,N_12583);
nor U12802 (N_12802,N_12530,N_12502);
nand U12803 (N_12803,N_12724,N_12729);
nor U12804 (N_12804,N_12540,N_12599);
nor U12805 (N_12805,N_12747,N_12638);
nor U12806 (N_12806,N_12678,N_12538);
nand U12807 (N_12807,N_12736,N_12546);
and U12808 (N_12808,N_12562,N_12570);
or U12809 (N_12809,N_12588,N_12661);
nor U12810 (N_12810,N_12676,N_12544);
nor U12811 (N_12811,N_12664,N_12508);
nand U12812 (N_12812,N_12725,N_12730);
or U12813 (N_12813,N_12633,N_12519);
nor U12814 (N_12814,N_12537,N_12630);
nand U12815 (N_12815,N_12720,N_12636);
nand U12816 (N_12816,N_12529,N_12582);
or U12817 (N_12817,N_12518,N_12658);
nor U12818 (N_12818,N_12631,N_12714);
and U12819 (N_12819,N_12719,N_12594);
nor U12820 (N_12820,N_12743,N_12597);
or U12821 (N_12821,N_12600,N_12651);
or U12822 (N_12822,N_12738,N_12692);
nand U12823 (N_12823,N_12681,N_12643);
and U12824 (N_12824,N_12525,N_12592);
nor U12825 (N_12825,N_12627,N_12732);
or U12826 (N_12826,N_12552,N_12581);
or U12827 (N_12827,N_12659,N_12500);
nand U12828 (N_12828,N_12579,N_12690);
or U12829 (N_12829,N_12613,N_12685);
nand U12830 (N_12830,N_12737,N_12605);
and U12831 (N_12831,N_12686,N_12695);
nor U12832 (N_12832,N_12637,N_12713);
and U12833 (N_12833,N_12501,N_12628);
or U12834 (N_12834,N_12580,N_12645);
nor U12835 (N_12835,N_12734,N_12688);
nor U12836 (N_12836,N_12611,N_12584);
nor U12837 (N_12837,N_12504,N_12735);
or U12838 (N_12838,N_12644,N_12566);
or U12839 (N_12839,N_12660,N_12545);
nand U12840 (N_12840,N_12656,N_12749);
or U12841 (N_12841,N_12512,N_12560);
nand U12842 (N_12842,N_12650,N_12705);
and U12843 (N_12843,N_12524,N_12673);
and U12844 (N_12844,N_12682,N_12683);
nor U12845 (N_12845,N_12578,N_12702);
or U12846 (N_12846,N_12585,N_12565);
and U12847 (N_12847,N_12667,N_12615);
nand U12848 (N_12848,N_12604,N_12569);
nand U12849 (N_12849,N_12679,N_12609);
nor U12850 (N_12850,N_12575,N_12703);
nand U12851 (N_12851,N_12704,N_12699);
and U12852 (N_12852,N_12624,N_12542);
and U12853 (N_12853,N_12744,N_12618);
or U12854 (N_12854,N_12740,N_12557);
nor U12855 (N_12855,N_12619,N_12666);
nand U12856 (N_12856,N_12510,N_12742);
nor U12857 (N_12857,N_12646,N_12543);
nand U12858 (N_12858,N_12591,N_12739);
or U12859 (N_12859,N_12532,N_12629);
and U12860 (N_12860,N_12672,N_12625);
or U12861 (N_12861,N_12632,N_12564);
nor U12862 (N_12862,N_12610,N_12522);
and U12863 (N_12863,N_12576,N_12626);
nand U12864 (N_12864,N_12555,N_12741);
nand U12865 (N_12865,N_12696,N_12528);
nand U12866 (N_12866,N_12617,N_12698);
or U12867 (N_12867,N_12654,N_12689);
and U12868 (N_12868,N_12746,N_12671);
and U12869 (N_12869,N_12684,N_12577);
or U12870 (N_12870,N_12706,N_12745);
and U12871 (N_12871,N_12716,N_12533);
and U12872 (N_12872,N_12516,N_12708);
and U12873 (N_12873,N_12548,N_12715);
nor U12874 (N_12874,N_12641,N_12612);
nor U12875 (N_12875,N_12522,N_12727);
nor U12876 (N_12876,N_12535,N_12714);
or U12877 (N_12877,N_12735,N_12616);
and U12878 (N_12878,N_12571,N_12690);
nor U12879 (N_12879,N_12635,N_12526);
nor U12880 (N_12880,N_12662,N_12635);
nor U12881 (N_12881,N_12503,N_12645);
or U12882 (N_12882,N_12501,N_12553);
and U12883 (N_12883,N_12657,N_12664);
and U12884 (N_12884,N_12704,N_12695);
or U12885 (N_12885,N_12588,N_12580);
or U12886 (N_12886,N_12674,N_12624);
or U12887 (N_12887,N_12595,N_12607);
and U12888 (N_12888,N_12685,N_12748);
nor U12889 (N_12889,N_12539,N_12537);
or U12890 (N_12890,N_12542,N_12744);
nor U12891 (N_12891,N_12737,N_12537);
or U12892 (N_12892,N_12660,N_12687);
or U12893 (N_12893,N_12722,N_12578);
nand U12894 (N_12894,N_12553,N_12601);
and U12895 (N_12895,N_12666,N_12736);
nand U12896 (N_12896,N_12601,N_12520);
nor U12897 (N_12897,N_12645,N_12536);
or U12898 (N_12898,N_12630,N_12627);
or U12899 (N_12899,N_12572,N_12570);
nand U12900 (N_12900,N_12659,N_12618);
or U12901 (N_12901,N_12567,N_12669);
nor U12902 (N_12902,N_12562,N_12531);
nand U12903 (N_12903,N_12664,N_12527);
nor U12904 (N_12904,N_12724,N_12659);
and U12905 (N_12905,N_12741,N_12719);
and U12906 (N_12906,N_12725,N_12712);
nand U12907 (N_12907,N_12514,N_12692);
xnor U12908 (N_12908,N_12719,N_12570);
nor U12909 (N_12909,N_12583,N_12569);
nor U12910 (N_12910,N_12630,N_12631);
nor U12911 (N_12911,N_12725,N_12649);
nand U12912 (N_12912,N_12530,N_12748);
nand U12913 (N_12913,N_12737,N_12713);
and U12914 (N_12914,N_12559,N_12564);
and U12915 (N_12915,N_12606,N_12655);
nor U12916 (N_12916,N_12615,N_12671);
nand U12917 (N_12917,N_12507,N_12629);
nand U12918 (N_12918,N_12552,N_12523);
nand U12919 (N_12919,N_12633,N_12682);
or U12920 (N_12920,N_12648,N_12701);
nand U12921 (N_12921,N_12540,N_12577);
nand U12922 (N_12922,N_12721,N_12653);
nand U12923 (N_12923,N_12542,N_12698);
nor U12924 (N_12924,N_12694,N_12625);
and U12925 (N_12925,N_12669,N_12621);
nand U12926 (N_12926,N_12671,N_12714);
nor U12927 (N_12927,N_12521,N_12500);
nor U12928 (N_12928,N_12602,N_12549);
nand U12929 (N_12929,N_12662,N_12673);
and U12930 (N_12930,N_12650,N_12679);
nand U12931 (N_12931,N_12742,N_12709);
nand U12932 (N_12932,N_12718,N_12593);
and U12933 (N_12933,N_12676,N_12514);
nor U12934 (N_12934,N_12609,N_12639);
nand U12935 (N_12935,N_12632,N_12748);
nor U12936 (N_12936,N_12716,N_12619);
or U12937 (N_12937,N_12577,N_12641);
or U12938 (N_12938,N_12748,N_12649);
or U12939 (N_12939,N_12623,N_12721);
nor U12940 (N_12940,N_12500,N_12701);
and U12941 (N_12941,N_12650,N_12504);
nor U12942 (N_12942,N_12700,N_12619);
nor U12943 (N_12943,N_12628,N_12670);
nor U12944 (N_12944,N_12710,N_12512);
nor U12945 (N_12945,N_12669,N_12640);
and U12946 (N_12946,N_12677,N_12642);
and U12947 (N_12947,N_12686,N_12517);
nor U12948 (N_12948,N_12720,N_12651);
and U12949 (N_12949,N_12540,N_12632);
nor U12950 (N_12950,N_12595,N_12725);
and U12951 (N_12951,N_12585,N_12559);
or U12952 (N_12952,N_12540,N_12677);
and U12953 (N_12953,N_12612,N_12741);
and U12954 (N_12954,N_12655,N_12527);
nand U12955 (N_12955,N_12545,N_12714);
or U12956 (N_12956,N_12682,N_12694);
nand U12957 (N_12957,N_12551,N_12701);
nand U12958 (N_12958,N_12502,N_12583);
nand U12959 (N_12959,N_12680,N_12562);
nor U12960 (N_12960,N_12691,N_12720);
or U12961 (N_12961,N_12728,N_12654);
and U12962 (N_12962,N_12663,N_12677);
xor U12963 (N_12963,N_12509,N_12579);
or U12964 (N_12964,N_12561,N_12681);
nor U12965 (N_12965,N_12652,N_12615);
nor U12966 (N_12966,N_12682,N_12595);
xnor U12967 (N_12967,N_12521,N_12640);
nand U12968 (N_12968,N_12581,N_12567);
and U12969 (N_12969,N_12540,N_12669);
nor U12970 (N_12970,N_12706,N_12550);
nor U12971 (N_12971,N_12660,N_12544);
nand U12972 (N_12972,N_12559,N_12649);
nand U12973 (N_12973,N_12500,N_12566);
or U12974 (N_12974,N_12614,N_12720);
or U12975 (N_12975,N_12681,N_12540);
or U12976 (N_12976,N_12739,N_12703);
or U12977 (N_12977,N_12722,N_12503);
or U12978 (N_12978,N_12718,N_12699);
nor U12979 (N_12979,N_12738,N_12633);
nand U12980 (N_12980,N_12654,N_12665);
and U12981 (N_12981,N_12630,N_12502);
and U12982 (N_12982,N_12680,N_12691);
nor U12983 (N_12983,N_12628,N_12547);
and U12984 (N_12984,N_12690,N_12600);
nand U12985 (N_12985,N_12672,N_12567);
nor U12986 (N_12986,N_12670,N_12701);
and U12987 (N_12987,N_12655,N_12626);
nor U12988 (N_12988,N_12746,N_12739);
or U12989 (N_12989,N_12689,N_12565);
or U12990 (N_12990,N_12627,N_12504);
nor U12991 (N_12991,N_12525,N_12608);
nor U12992 (N_12992,N_12637,N_12572);
and U12993 (N_12993,N_12517,N_12639);
nand U12994 (N_12994,N_12582,N_12689);
or U12995 (N_12995,N_12577,N_12648);
nor U12996 (N_12996,N_12640,N_12658);
or U12997 (N_12997,N_12505,N_12661);
or U12998 (N_12998,N_12502,N_12693);
nor U12999 (N_12999,N_12722,N_12698);
nor U13000 (N_13000,N_12821,N_12801);
or U13001 (N_13001,N_12756,N_12762);
nand U13002 (N_13002,N_12933,N_12826);
nand U13003 (N_13003,N_12780,N_12992);
nor U13004 (N_13004,N_12943,N_12911);
or U13005 (N_13005,N_12881,N_12897);
nor U13006 (N_13006,N_12833,N_12787);
and U13007 (N_13007,N_12949,N_12925);
nand U13008 (N_13008,N_12868,N_12975);
or U13009 (N_13009,N_12853,N_12812);
xor U13010 (N_13010,N_12841,N_12888);
and U13011 (N_13011,N_12993,N_12931);
nor U13012 (N_13012,N_12921,N_12919);
nor U13013 (N_13013,N_12983,N_12770);
nor U13014 (N_13014,N_12832,N_12773);
nand U13015 (N_13015,N_12968,N_12816);
or U13016 (N_13016,N_12935,N_12909);
and U13017 (N_13017,N_12761,N_12807);
nor U13018 (N_13018,N_12959,N_12858);
nand U13019 (N_13019,N_12910,N_12890);
or U13020 (N_13020,N_12808,N_12784);
or U13021 (N_13021,N_12991,N_12914);
nor U13022 (N_13022,N_12994,N_12779);
nor U13023 (N_13023,N_12940,N_12892);
or U13024 (N_13024,N_12789,N_12901);
nand U13025 (N_13025,N_12978,N_12945);
and U13026 (N_13026,N_12989,N_12844);
nand U13027 (N_13027,N_12995,N_12848);
nand U13028 (N_13028,N_12946,N_12786);
nor U13029 (N_13029,N_12857,N_12750);
nand U13030 (N_13030,N_12781,N_12842);
and U13031 (N_13031,N_12904,N_12818);
or U13032 (N_13032,N_12755,N_12934);
xor U13033 (N_13033,N_12976,N_12837);
nor U13034 (N_13034,N_12898,N_12856);
or U13035 (N_13035,N_12954,N_12894);
or U13036 (N_13036,N_12906,N_12889);
xnor U13037 (N_13037,N_12777,N_12916);
nand U13038 (N_13038,N_12928,N_12969);
or U13039 (N_13039,N_12938,N_12822);
and U13040 (N_13040,N_12918,N_12964);
or U13041 (N_13041,N_12942,N_12776);
and U13042 (N_13042,N_12820,N_12893);
nor U13043 (N_13043,N_12852,N_12758);
nand U13044 (N_13044,N_12955,N_12751);
nand U13045 (N_13045,N_12797,N_12865);
nand U13046 (N_13046,N_12835,N_12800);
and U13047 (N_13047,N_12956,N_12887);
nor U13048 (N_13048,N_12971,N_12917);
and U13049 (N_13049,N_12802,N_12859);
and U13050 (N_13050,N_12899,N_12782);
or U13051 (N_13051,N_12951,N_12783);
nor U13052 (N_13052,N_12900,N_12847);
nor U13053 (N_13053,N_12774,N_12997);
and U13054 (N_13054,N_12882,N_12813);
and U13055 (N_13055,N_12923,N_12905);
nand U13056 (N_13056,N_12984,N_12757);
nand U13057 (N_13057,N_12752,N_12966);
or U13058 (N_13058,N_12869,N_12759);
or U13059 (N_13059,N_12815,N_12877);
or U13060 (N_13060,N_12788,N_12936);
nor U13061 (N_13061,N_12962,N_12965);
nor U13062 (N_13062,N_12861,N_12769);
or U13063 (N_13063,N_12768,N_12947);
and U13064 (N_13064,N_12885,N_12793);
nor U13065 (N_13065,N_12834,N_12760);
nor U13066 (N_13066,N_12957,N_12778);
nand U13067 (N_13067,N_12825,N_12836);
nor U13068 (N_13068,N_12948,N_12950);
nor U13069 (N_13069,N_12952,N_12831);
nand U13070 (N_13070,N_12884,N_12765);
and U13071 (N_13071,N_12796,N_12990);
and U13072 (N_13072,N_12871,N_12985);
and U13073 (N_13073,N_12932,N_12794);
nor U13074 (N_13074,N_12875,N_12874);
or U13075 (N_13075,N_12754,N_12790);
or U13076 (N_13076,N_12915,N_12814);
nand U13077 (N_13077,N_12799,N_12850);
nand U13078 (N_13078,N_12840,N_12939);
nor U13079 (N_13079,N_12903,N_12772);
nand U13080 (N_13080,N_12974,N_12902);
and U13081 (N_13081,N_12977,N_12827);
nor U13082 (N_13082,N_12810,N_12920);
and U13083 (N_13083,N_12843,N_12960);
nand U13084 (N_13084,N_12876,N_12922);
nor U13085 (N_13085,N_12880,N_12879);
nand U13086 (N_13086,N_12775,N_12980);
nor U13087 (N_13087,N_12883,N_12866);
and U13088 (N_13088,N_12766,N_12873);
nand U13089 (N_13089,N_12926,N_12792);
nand U13090 (N_13090,N_12771,N_12927);
nand U13091 (N_13091,N_12806,N_12849);
or U13092 (N_13092,N_12941,N_12864);
or U13093 (N_13093,N_12838,N_12981);
or U13094 (N_13094,N_12970,N_12798);
nand U13095 (N_13095,N_12785,N_12886);
and U13096 (N_13096,N_12867,N_12828);
and U13097 (N_13097,N_12830,N_12958);
nand U13098 (N_13098,N_12988,N_12863);
nand U13099 (N_13099,N_12961,N_12823);
nor U13100 (N_13100,N_12817,N_12862);
nor U13101 (N_13101,N_12953,N_12896);
nor U13102 (N_13102,N_12982,N_12963);
nand U13103 (N_13103,N_12764,N_12753);
and U13104 (N_13104,N_12908,N_12891);
nor U13105 (N_13105,N_12986,N_12973);
nand U13106 (N_13106,N_12845,N_12913);
or U13107 (N_13107,N_12929,N_12854);
and U13108 (N_13108,N_12878,N_12972);
nand U13109 (N_13109,N_12907,N_12924);
nor U13110 (N_13110,N_12860,N_12805);
nand U13111 (N_13111,N_12839,N_12944);
and U13112 (N_13112,N_12795,N_12809);
and U13113 (N_13113,N_12979,N_12937);
nor U13114 (N_13114,N_12791,N_12846);
nor U13115 (N_13115,N_12851,N_12895);
or U13116 (N_13116,N_12763,N_12811);
or U13117 (N_13117,N_12872,N_12804);
nand U13118 (N_13118,N_12870,N_12767);
and U13119 (N_13119,N_12819,N_12987);
or U13120 (N_13120,N_12829,N_12930);
and U13121 (N_13121,N_12998,N_12967);
nand U13122 (N_13122,N_12999,N_12855);
and U13123 (N_13123,N_12803,N_12912);
and U13124 (N_13124,N_12824,N_12996);
nand U13125 (N_13125,N_12872,N_12966);
nor U13126 (N_13126,N_12818,N_12821);
nor U13127 (N_13127,N_12938,N_12919);
nor U13128 (N_13128,N_12758,N_12783);
nor U13129 (N_13129,N_12864,N_12784);
nand U13130 (N_13130,N_12934,N_12858);
nor U13131 (N_13131,N_12791,N_12944);
or U13132 (N_13132,N_12940,N_12877);
and U13133 (N_13133,N_12928,N_12943);
and U13134 (N_13134,N_12926,N_12973);
or U13135 (N_13135,N_12967,N_12950);
and U13136 (N_13136,N_12871,N_12816);
nand U13137 (N_13137,N_12790,N_12765);
and U13138 (N_13138,N_12798,N_12911);
nor U13139 (N_13139,N_12892,N_12866);
or U13140 (N_13140,N_12948,N_12794);
nand U13141 (N_13141,N_12962,N_12834);
nor U13142 (N_13142,N_12782,N_12758);
nand U13143 (N_13143,N_12978,N_12898);
nor U13144 (N_13144,N_12783,N_12821);
nand U13145 (N_13145,N_12998,N_12798);
nand U13146 (N_13146,N_12898,N_12792);
and U13147 (N_13147,N_12846,N_12924);
nand U13148 (N_13148,N_12995,N_12871);
nand U13149 (N_13149,N_12797,N_12774);
and U13150 (N_13150,N_12963,N_12847);
or U13151 (N_13151,N_12940,N_12867);
nand U13152 (N_13152,N_12801,N_12996);
nor U13153 (N_13153,N_12976,N_12953);
nand U13154 (N_13154,N_12963,N_12825);
or U13155 (N_13155,N_12986,N_12772);
and U13156 (N_13156,N_12821,N_12836);
xnor U13157 (N_13157,N_12760,N_12860);
nor U13158 (N_13158,N_12810,N_12932);
nand U13159 (N_13159,N_12914,N_12865);
or U13160 (N_13160,N_12984,N_12910);
nor U13161 (N_13161,N_12855,N_12932);
nand U13162 (N_13162,N_12900,N_12778);
nor U13163 (N_13163,N_12873,N_12987);
or U13164 (N_13164,N_12812,N_12898);
nand U13165 (N_13165,N_12860,N_12802);
nand U13166 (N_13166,N_12797,N_12884);
nor U13167 (N_13167,N_12835,N_12833);
nor U13168 (N_13168,N_12936,N_12844);
or U13169 (N_13169,N_12785,N_12880);
or U13170 (N_13170,N_12949,N_12821);
nor U13171 (N_13171,N_12891,N_12948);
and U13172 (N_13172,N_12787,N_12868);
nor U13173 (N_13173,N_12952,N_12860);
or U13174 (N_13174,N_12879,N_12888);
nor U13175 (N_13175,N_12936,N_12945);
nor U13176 (N_13176,N_12763,N_12768);
or U13177 (N_13177,N_12943,N_12827);
xor U13178 (N_13178,N_12758,N_12908);
or U13179 (N_13179,N_12876,N_12786);
nor U13180 (N_13180,N_12954,N_12836);
nand U13181 (N_13181,N_12832,N_12902);
nand U13182 (N_13182,N_12906,N_12854);
nor U13183 (N_13183,N_12951,N_12977);
xnor U13184 (N_13184,N_12866,N_12837);
and U13185 (N_13185,N_12843,N_12847);
nand U13186 (N_13186,N_12881,N_12990);
or U13187 (N_13187,N_12956,N_12761);
or U13188 (N_13188,N_12873,N_12979);
nor U13189 (N_13189,N_12990,N_12955);
nand U13190 (N_13190,N_12856,N_12953);
nand U13191 (N_13191,N_12903,N_12916);
and U13192 (N_13192,N_12949,N_12863);
nor U13193 (N_13193,N_12963,N_12846);
xor U13194 (N_13194,N_12915,N_12768);
nand U13195 (N_13195,N_12887,N_12997);
nor U13196 (N_13196,N_12852,N_12815);
nor U13197 (N_13197,N_12921,N_12984);
and U13198 (N_13198,N_12963,N_12969);
and U13199 (N_13199,N_12945,N_12909);
or U13200 (N_13200,N_12941,N_12847);
or U13201 (N_13201,N_12788,N_12954);
or U13202 (N_13202,N_12942,N_12956);
and U13203 (N_13203,N_12904,N_12826);
nand U13204 (N_13204,N_12858,N_12936);
nor U13205 (N_13205,N_12957,N_12886);
nor U13206 (N_13206,N_12899,N_12840);
nor U13207 (N_13207,N_12775,N_12977);
nand U13208 (N_13208,N_12868,N_12933);
nor U13209 (N_13209,N_12861,N_12934);
nor U13210 (N_13210,N_12814,N_12831);
nand U13211 (N_13211,N_12801,N_12948);
nand U13212 (N_13212,N_12750,N_12894);
or U13213 (N_13213,N_12946,N_12811);
or U13214 (N_13214,N_12904,N_12780);
or U13215 (N_13215,N_12801,N_12795);
or U13216 (N_13216,N_12945,N_12905);
and U13217 (N_13217,N_12946,N_12890);
nand U13218 (N_13218,N_12935,N_12762);
and U13219 (N_13219,N_12854,N_12771);
and U13220 (N_13220,N_12797,N_12821);
or U13221 (N_13221,N_12901,N_12842);
nand U13222 (N_13222,N_12824,N_12780);
nor U13223 (N_13223,N_12791,N_12773);
and U13224 (N_13224,N_12855,N_12891);
nor U13225 (N_13225,N_12764,N_12992);
or U13226 (N_13226,N_12954,N_12759);
or U13227 (N_13227,N_12854,N_12894);
or U13228 (N_13228,N_12968,N_12845);
nor U13229 (N_13229,N_12846,N_12888);
or U13230 (N_13230,N_12764,N_12766);
nand U13231 (N_13231,N_12830,N_12954);
or U13232 (N_13232,N_12866,N_12869);
nand U13233 (N_13233,N_12798,N_12997);
nand U13234 (N_13234,N_12995,N_12852);
nor U13235 (N_13235,N_12935,N_12971);
nand U13236 (N_13236,N_12814,N_12871);
and U13237 (N_13237,N_12886,N_12768);
or U13238 (N_13238,N_12822,N_12751);
and U13239 (N_13239,N_12915,N_12992);
or U13240 (N_13240,N_12802,N_12805);
and U13241 (N_13241,N_12782,N_12965);
nor U13242 (N_13242,N_12912,N_12835);
nor U13243 (N_13243,N_12990,N_12982);
nand U13244 (N_13244,N_12806,N_12757);
nor U13245 (N_13245,N_12861,N_12772);
xor U13246 (N_13246,N_12924,N_12760);
and U13247 (N_13247,N_12972,N_12877);
or U13248 (N_13248,N_12808,N_12792);
nor U13249 (N_13249,N_12847,N_12948);
nor U13250 (N_13250,N_13222,N_13084);
and U13251 (N_13251,N_13154,N_13020);
xnor U13252 (N_13252,N_13002,N_13055);
nand U13253 (N_13253,N_13120,N_13219);
nor U13254 (N_13254,N_13122,N_13177);
nand U13255 (N_13255,N_13054,N_13212);
xnor U13256 (N_13256,N_13062,N_13076);
nor U13257 (N_13257,N_13053,N_13081);
nand U13258 (N_13258,N_13206,N_13153);
or U13259 (N_13259,N_13190,N_13136);
nand U13260 (N_13260,N_13021,N_13189);
or U13261 (N_13261,N_13051,N_13188);
nand U13262 (N_13262,N_13080,N_13075);
or U13263 (N_13263,N_13155,N_13126);
or U13264 (N_13264,N_13235,N_13152);
nand U13265 (N_13265,N_13245,N_13224);
nor U13266 (N_13266,N_13160,N_13073);
nand U13267 (N_13267,N_13181,N_13230);
nand U13268 (N_13268,N_13040,N_13172);
or U13269 (N_13269,N_13241,N_13010);
nand U13270 (N_13270,N_13159,N_13134);
nor U13271 (N_13271,N_13066,N_13028);
and U13272 (N_13272,N_13201,N_13070);
nand U13273 (N_13273,N_13069,N_13146);
nand U13274 (N_13274,N_13128,N_13005);
or U13275 (N_13275,N_13068,N_13242);
and U13276 (N_13276,N_13141,N_13077);
nor U13277 (N_13277,N_13197,N_13063);
nand U13278 (N_13278,N_13047,N_13158);
nor U13279 (N_13279,N_13100,N_13228);
nand U13280 (N_13280,N_13096,N_13173);
and U13281 (N_13281,N_13044,N_13238);
nand U13282 (N_13282,N_13210,N_13031);
xor U13283 (N_13283,N_13208,N_13161);
and U13284 (N_13284,N_13101,N_13150);
nand U13285 (N_13285,N_13112,N_13137);
nor U13286 (N_13286,N_13102,N_13038);
nor U13287 (N_13287,N_13168,N_13133);
nand U13288 (N_13288,N_13016,N_13200);
xor U13289 (N_13289,N_13113,N_13083);
nor U13290 (N_13290,N_13111,N_13012);
nor U13291 (N_13291,N_13204,N_13139);
or U13292 (N_13292,N_13087,N_13032);
or U13293 (N_13293,N_13202,N_13024);
and U13294 (N_13294,N_13240,N_13116);
nor U13295 (N_13295,N_13013,N_13034);
and U13296 (N_13296,N_13018,N_13037);
and U13297 (N_13297,N_13079,N_13050);
nor U13298 (N_13298,N_13019,N_13138);
and U13299 (N_13299,N_13052,N_13184);
nor U13300 (N_13300,N_13004,N_13125);
nor U13301 (N_13301,N_13108,N_13085);
or U13302 (N_13302,N_13180,N_13022);
and U13303 (N_13303,N_13223,N_13175);
and U13304 (N_13304,N_13178,N_13135);
nor U13305 (N_13305,N_13248,N_13000);
nor U13306 (N_13306,N_13213,N_13114);
and U13307 (N_13307,N_13218,N_13104);
nor U13308 (N_13308,N_13029,N_13234);
and U13309 (N_13309,N_13232,N_13151);
nand U13310 (N_13310,N_13209,N_13045);
nor U13311 (N_13311,N_13086,N_13140);
and U13312 (N_13312,N_13127,N_13131);
nor U13313 (N_13313,N_13095,N_13191);
or U13314 (N_13314,N_13129,N_13064);
or U13315 (N_13315,N_13119,N_13014);
and U13316 (N_13316,N_13030,N_13237);
nand U13317 (N_13317,N_13067,N_13233);
nand U13318 (N_13318,N_13121,N_13078);
or U13319 (N_13319,N_13124,N_13166);
nor U13320 (N_13320,N_13174,N_13149);
or U13321 (N_13321,N_13229,N_13183);
nand U13322 (N_13322,N_13198,N_13033);
nand U13323 (N_13323,N_13236,N_13249);
nor U13324 (N_13324,N_13221,N_13061);
nand U13325 (N_13325,N_13057,N_13042);
nor U13326 (N_13326,N_13003,N_13093);
nor U13327 (N_13327,N_13110,N_13176);
or U13328 (N_13328,N_13058,N_13049);
or U13329 (N_13329,N_13098,N_13006);
nand U13330 (N_13330,N_13106,N_13107);
and U13331 (N_13331,N_13001,N_13071);
and U13332 (N_13332,N_13036,N_13059);
and U13333 (N_13333,N_13041,N_13163);
and U13334 (N_13334,N_13142,N_13164);
nor U13335 (N_13335,N_13105,N_13089);
nor U13336 (N_13336,N_13148,N_13231);
nand U13337 (N_13337,N_13097,N_13060);
and U13338 (N_13338,N_13090,N_13074);
and U13339 (N_13339,N_13072,N_13179);
and U13340 (N_13340,N_13220,N_13169);
or U13341 (N_13341,N_13167,N_13196);
or U13342 (N_13342,N_13046,N_13007);
and U13343 (N_13343,N_13216,N_13192);
and U13344 (N_13344,N_13117,N_13011);
and U13345 (N_13345,N_13094,N_13227);
nor U13346 (N_13346,N_13182,N_13144);
nor U13347 (N_13347,N_13043,N_13185);
nand U13348 (N_13348,N_13145,N_13156);
or U13349 (N_13349,N_13143,N_13027);
and U13350 (N_13350,N_13091,N_13203);
nor U13351 (N_13351,N_13195,N_13035);
or U13352 (N_13352,N_13115,N_13170);
and U13353 (N_13353,N_13205,N_13048);
nor U13354 (N_13354,N_13244,N_13065);
and U13355 (N_13355,N_13039,N_13109);
or U13356 (N_13356,N_13023,N_13132);
and U13357 (N_13357,N_13194,N_13088);
nor U13358 (N_13358,N_13243,N_13092);
or U13359 (N_13359,N_13186,N_13193);
and U13360 (N_13360,N_13015,N_13225);
or U13361 (N_13361,N_13017,N_13118);
and U13362 (N_13362,N_13214,N_13025);
nand U13363 (N_13363,N_13239,N_13171);
nor U13364 (N_13364,N_13103,N_13207);
nand U13365 (N_13365,N_13215,N_13026);
nand U13366 (N_13366,N_13226,N_13217);
nand U13367 (N_13367,N_13247,N_13246);
or U13368 (N_13368,N_13199,N_13157);
nor U13369 (N_13369,N_13082,N_13056);
or U13370 (N_13370,N_13130,N_13147);
or U13371 (N_13371,N_13009,N_13187);
nand U13372 (N_13372,N_13123,N_13008);
or U13373 (N_13373,N_13211,N_13162);
nor U13374 (N_13374,N_13099,N_13165);
and U13375 (N_13375,N_13012,N_13211);
nor U13376 (N_13376,N_13038,N_13242);
or U13377 (N_13377,N_13050,N_13188);
nand U13378 (N_13378,N_13249,N_13038);
and U13379 (N_13379,N_13140,N_13191);
and U13380 (N_13380,N_13182,N_13139);
nor U13381 (N_13381,N_13145,N_13118);
or U13382 (N_13382,N_13123,N_13022);
or U13383 (N_13383,N_13169,N_13219);
and U13384 (N_13384,N_13007,N_13094);
nor U13385 (N_13385,N_13058,N_13080);
nand U13386 (N_13386,N_13193,N_13175);
and U13387 (N_13387,N_13247,N_13209);
and U13388 (N_13388,N_13169,N_13183);
xor U13389 (N_13389,N_13037,N_13199);
nor U13390 (N_13390,N_13073,N_13223);
nand U13391 (N_13391,N_13188,N_13002);
nand U13392 (N_13392,N_13248,N_13180);
and U13393 (N_13393,N_13129,N_13178);
nand U13394 (N_13394,N_13171,N_13183);
nor U13395 (N_13395,N_13128,N_13165);
or U13396 (N_13396,N_13187,N_13159);
and U13397 (N_13397,N_13128,N_13131);
nor U13398 (N_13398,N_13212,N_13174);
nand U13399 (N_13399,N_13037,N_13106);
nor U13400 (N_13400,N_13120,N_13071);
or U13401 (N_13401,N_13185,N_13044);
nor U13402 (N_13402,N_13225,N_13186);
nand U13403 (N_13403,N_13211,N_13226);
or U13404 (N_13404,N_13032,N_13223);
nor U13405 (N_13405,N_13168,N_13039);
and U13406 (N_13406,N_13154,N_13141);
nor U13407 (N_13407,N_13076,N_13221);
or U13408 (N_13408,N_13024,N_13196);
or U13409 (N_13409,N_13061,N_13231);
or U13410 (N_13410,N_13015,N_13243);
and U13411 (N_13411,N_13121,N_13144);
nand U13412 (N_13412,N_13040,N_13118);
nand U13413 (N_13413,N_13037,N_13225);
and U13414 (N_13414,N_13038,N_13091);
or U13415 (N_13415,N_13241,N_13073);
and U13416 (N_13416,N_13210,N_13006);
nor U13417 (N_13417,N_13226,N_13012);
and U13418 (N_13418,N_13071,N_13007);
or U13419 (N_13419,N_13230,N_13190);
nor U13420 (N_13420,N_13236,N_13238);
nand U13421 (N_13421,N_13132,N_13078);
or U13422 (N_13422,N_13232,N_13025);
nand U13423 (N_13423,N_13190,N_13210);
and U13424 (N_13424,N_13168,N_13190);
nand U13425 (N_13425,N_13081,N_13133);
nand U13426 (N_13426,N_13104,N_13186);
or U13427 (N_13427,N_13007,N_13114);
or U13428 (N_13428,N_13034,N_13078);
nand U13429 (N_13429,N_13151,N_13072);
nor U13430 (N_13430,N_13034,N_13072);
and U13431 (N_13431,N_13188,N_13046);
nor U13432 (N_13432,N_13233,N_13244);
nand U13433 (N_13433,N_13207,N_13109);
nand U13434 (N_13434,N_13159,N_13092);
and U13435 (N_13435,N_13120,N_13231);
nand U13436 (N_13436,N_13018,N_13097);
or U13437 (N_13437,N_13197,N_13244);
nand U13438 (N_13438,N_13091,N_13103);
or U13439 (N_13439,N_13047,N_13009);
nor U13440 (N_13440,N_13080,N_13026);
or U13441 (N_13441,N_13108,N_13107);
nor U13442 (N_13442,N_13131,N_13203);
xor U13443 (N_13443,N_13123,N_13172);
and U13444 (N_13444,N_13215,N_13237);
or U13445 (N_13445,N_13210,N_13046);
or U13446 (N_13446,N_13158,N_13071);
or U13447 (N_13447,N_13148,N_13136);
nor U13448 (N_13448,N_13009,N_13050);
or U13449 (N_13449,N_13098,N_13242);
nor U13450 (N_13450,N_13036,N_13089);
or U13451 (N_13451,N_13245,N_13074);
or U13452 (N_13452,N_13244,N_13194);
and U13453 (N_13453,N_13108,N_13062);
nand U13454 (N_13454,N_13081,N_13097);
nor U13455 (N_13455,N_13027,N_13197);
nor U13456 (N_13456,N_13133,N_13118);
nand U13457 (N_13457,N_13129,N_13132);
and U13458 (N_13458,N_13075,N_13158);
nor U13459 (N_13459,N_13147,N_13050);
nand U13460 (N_13460,N_13089,N_13169);
nand U13461 (N_13461,N_13190,N_13148);
and U13462 (N_13462,N_13152,N_13063);
nand U13463 (N_13463,N_13232,N_13019);
xor U13464 (N_13464,N_13152,N_13189);
nor U13465 (N_13465,N_13242,N_13214);
nor U13466 (N_13466,N_13000,N_13236);
nor U13467 (N_13467,N_13061,N_13148);
or U13468 (N_13468,N_13184,N_13059);
xnor U13469 (N_13469,N_13208,N_13024);
or U13470 (N_13470,N_13086,N_13176);
nand U13471 (N_13471,N_13133,N_13146);
nor U13472 (N_13472,N_13205,N_13149);
and U13473 (N_13473,N_13135,N_13189);
or U13474 (N_13474,N_13246,N_13147);
xnor U13475 (N_13475,N_13162,N_13102);
nand U13476 (N_13476,N_13008,N_13159);
nor U13477 (N_13477,N_13098,N_13115);
or U13478 (N_13478,N_13114,N_13049);
or U13479 (N_13479,N_13120,N_13149);
nor U13480 (N_13480,N_13085,N_13056);
or U13481 (N_13481,N_13134,N_13093);
and U13482 (N_13482,N_13192,N_13021);
or U13483 (N_13483,N_13037,N_13197);
nor U13484 (N_13484,N_13130,N_13142);
or U13485 (N_13485,N_13022,N_13202);
or U13486 (N_13486,N_13031,N_13183);
and U13487 (N_13487,N_13145,N_13191);
or U13488 (N_13488,N_13130,N_13222);
and U13489 (N_13489,N_13244,N_13243);
nand U13490 (N_13490,N_13120,N_13131);
nand U13491 (N_13491,N_13027,N_13044);
and U13492 (N_13492,N_13196,N_13044);
nor U13493 (N_13493,N_13132,N_13053);
or U13494 (N_13494,N_13206,N_13017);
xor U13495 (N_13495,N_13214,N_13102);
nor U13496 (N_13496,N_13200,N_13008);
nand U13497 (N_13497,N_13042,N_13098);
and U13498 (N_13498,N_13062,N_13126);
nor U13499 (N_13499,N_13223,N_13068);
nor U13500 (N_13500,N_13459,N_13294);
nor U13501 (N_13501,N_13277,N_13349);
or U13502 (N_13502,N_13333,N_13412);
nor U13503 (N_13503,N_13490,N_13324);
or U13504 (N_13504,N_13458,N_13291);
and U13505 (N_13505,N_13356,N_13382);
nand U13506 (N_13506,N_13334,N_13481);
nand U13507 (N_13507,N_13306,N_13394);
and U13508 (N_13508,N_13397,N_13275);
and U13509 (N_13509,N_13494,N_13474);
and U13510 (N_13510,N_13461,N_13423);
nand U13511 (N_13511,N_13337,N_13331);
nor U13512 (N_13512,N_13477,N_13390);
or U13513 (N_13513,N_13319,N_13431);
nand U13514 (N_13514,N_13419,N_13372);
and U13515 (N_13515,N_13491,N_13395);
and U13516 (N_13516,N_13411,N_13449);
nand U13517 (N_13517,N_13311,N_13376);
nor U13518 (N_13518,N_13389,N_13295);
nand U13519 (N_13519,N_13385,N_13377);
and U13520 (N_13520,N_13262,N_13417);
or U13521 (N_13521,N_13384,N_13393);
or U13522 (N_13522,N_13413,N_13342);
xor U13523 (N_13523,N_13332,N_13261);
nand U13524 (N_13524,N_13454,N_13338);
nor U13525 (N_13525,N_13369,N_13478);
nor U13526 (N_13526,N_13355,N_13406);
nor U13527 (N_13527,N_13433,N_13467);
or U13528 (N_13528,N_13399,N_13301);
and U13529 (N_13529,N_13391,N_13363);
and U13530 (N_13530,N_13466,N_13407);
nand U13531 (N_13531,N_13316,N_13489);
and U13532 (N_13532,N_13348,N_13401);
nand U13533 (N_13533,N_13396,N_13498);
nor U13534 (N_13534,N_13476,N_13297);
and U13535 (N_13535,N_13367,N_13444);
nand U13536 (N_13536,N_13254,N_13317);
nor U13537 (N_13537,N_13462,N_13463);
nor U13538 (N_13538,N_13480,N_13373);
nand U13539 (N_13539,N_13264,N_13460);
xor U13540 (N_13540,N_13361,N_13370);
xnor U13541 (N_13541,N_13434,N_13487);
nor U13542 (N_13542,N_13256,N_13479);
or U13543 (N_13543,N_13260,N_13402);
and U13544 (N_13544,N_13299,N_13421);
or U13545 (N_13545,N_13440,N_13410);
nor U13546 (N_13546,N_13329,N_13308);
or U13547 (N_13547,N_13379,N_13496);
nand U13548 (N_13548,N_13469,N_13427);
or U13549 (N_13549,N_13259,N_13403);
nand U13550 (N_13550,N_13252,N_13271);
or U13551 (N_13551,N_13457,N_13298);
or U13552 (N_13552,N_13300,N_13339);
nand U13553 (N_13553,N_13255,N_13253);
nand U13554 (N_13554,N_13442,N_13352);
or U13555 (N_13555,N_13430,N_13375);
or U13556 (N_13556,N_13280,N_13320);
xnor U13557 (N_13557,N_13428,N_13350);
or U13558 (N_13558,N_13282,N_13445);
nor U13559 (N_13559,N_13269,N_13371);
xnor U13560 (N_13560,N_13270,N_13327);
nor U13561 (N_13561,N_13416,N_13482);
nor U13562 (N_13562,N_13472,N_13485);
and U13563 (N_13563,N_13447,N_13383);
nand U13564 (N_13564,N_13415,N_13464);
and U13565 (N_13565,N_13388,N_13404);
nand U13566 (N_13566,N_13314,N_13340);
nand U13567 (N_13567,N_13307,N_13368);
nand U13568 (N_13568,N_13330,N_13343);
nor U13569 (N_13569,N_13336,N_13290);
and U13570 (N_13570,N_13360,N_13437);
and U13571 (N_13571,N_13288,N_13344);
nor U13572 (N_13572,N_13499,N_13456);
nor U13573 (N_13573,N_13424,N_13303);
nor U13574 (N_13574,N_13465,N_13283);
and U13575 (N_13575,N_13439,N_13436);
or U13576 (N_13576,N_13276,N_13287);
nand U13577 (N_13577,N_13279,N_13258);
nand U13578 (N_13578,N_13273,N_13351);
nand U13579 (N_13579,N_13378,N_13400);
nand U13580 (N_13580,N_13446,N_13278);
nor U13581 (N_13581,N_13274,N_13451);
nand U13582 (N_13582,N_13285,N_13492);
nand U13583 (N_13583,N_13328,N_13268);
or U13584 (N_13584,N_13321,N_13289);
nand U13585 (N_13585,N_13263,N_13475);
nor U13586 (N_13586,N_13380,N_13325);
or U13587 (N_13587,N_13470,N_13432);
nor U13588 (N_13588,N_13408,N_13364);
or U13589 (N_13589,N_13353,N_13405);
and U13590 (N_13590,N_13358,N_13296);
nand U13591 (N_13591,N_13292,N_13335);
nor U13592 (N_13592,N_13251,N_13354);
nand U13593 (N_13593,N_13323,N_13315);
nand U13594 (N_13594,N_13365,N_13293);
nand U13595 (N_13595,N_13266,N_13429);
nand U13596 (N_13596,N_13357,N_13386);
or U13597 (N_13597,N_13359,N_13302);
nor U13598 (N_13598,N_13435,N_13473);
and U13599 (N_13599,N_13448,N_13450);
and U13600 (N_13600,N_13486,N_13366);
nor U13601 (N_13601,N_13286,N_13326);
or U13602 (N_13602,N_13272,N_13322);
or U13603 (N_13603,N_13452,N_13443);
nor U13604 (N_13604,N_13284,N_13312);
and U13605 (N_13605,N_13398,N_13414);
nor U13606 (N_13606,N_13392,N_13471);
nand U13607 (N_13607,N_13310,N_13438);
nor U13608 (N_13608,N_13453,N_13346);
nor U13609 (N_13609,N_13257,N_13265);
and U13610 (N_13610,N_13409,N_13250);
and U13611 (N_13611,N_13455,N_13493);
or U13612 (N_13612,N_13483,N_13425);
and U13613 (N_13613,N_13387,N_13305);
nand U13614 (N_13614,N_13345,N_13341);
and U13615 (N_13615,N_13267,N_13441);
nand U13616 (N_13616,N_13313,N_13495);
nand U13617 (N_13617,N_13426,N_13420);
nor U13618 (N_13618,N_13347,N_13381);
nand U13619 (N_13619,N_13484,N_13281);
xnor U13620 (N_13620,N_13418,N_13488);
or U13621 (N_13621,N_13374,N_13362);
nor U13622 (N_13622,N_13304,N_13318);
nand U13623 (N_13623,N_13497,N_13309);
and U13624 (N_13624,N_13422,N_13468);
nor U13625 (N_13625,N_13279,N_13308);
nor U13626 (N_13626,N_13346,N_13403);
and U13627 (N_13627,N_13302,N_13399);
nor U13628 (N_13628,N_13293,N_13348);
and U13629 (N_13629,N_13480,N_13485);
nor U13630 (N_13630,N_13396,N_13333);
nand U13631 (N_13631,N_13452,N_13466);
or U13632 (N_13632,N_13288,N_13498);
nor U13633 (N_13633,N_13369,N_13469);
and U13634 (N_13634,N_13431,N_13377);
or U13635 (N_13635,N_13483,N_13265);
and U13636 (N_13636,N_13430,N_13373);
or U13637 (N_13637,N_13339,N_13492);
or U13638 (N_13638,N_13331,N_13441);
nor U13639 (N_13639,N_13268,N_13424);
nand U13640 (N_13640,N_13368,N_13440);
or U13641 (N_13641,N_13286,N_13481);
nand U13642 (N_13642,N_13362,N_13414);
nor U13643 (N_13643,N_13465,N_13433);
nor U13644 (N_13644,N_13294,N_13471);
or U13645 (N_13645,N_13368,N_13430);
or U13646 (N_13646,N_13454,N_13335);
and U13647 (N_13647,N_13441,N_13302);
or U13648 (N_13648,N_13460,N_13308);
or U13649 (N_13649,N_13492,N_13461);
nand U13650 (N_13650,N_13450,N_13277);
and U13651 (N_13651,N_13467,N_13344);
xor U13652 (N_13652,N_13254,N_13272);
nor U13653 (N_13653,N_13456,N_13275);
and U13654 (N_13654,N_13400,N_13401);
nor U13655 (N_13655,N_13496,N_13399);
xnor U13656 (N_13656,N_13399,N_13298);
or U13657 (N_13657,N_13484,N_13362);
and U13658 (N_13658,N_13377,N_13346);
nor U13659 (N_13659,N_13275,N_13457);
nand U13660 (N_13660,N_13483,N_13496);
or U13661 (N_13661,N_13487,N_13459);
nor U13662 (N_13662,N_13449,N_13414);
nand U13663 (N_13663,N_13268,N_13430);
and U13664 (N_13664,N_13464,N_13250);
and U13665 (N_13665,N_13287,N_13337);
nor U13666 (N_13666,N_13340,N_13453);
nand U13667 (N_13667,N_13345,N_13312);
or U13668 (N_13668,N_13301,N_13376);
or U13669 (N_13669,N_13431,N_13461);
and U13670 (N_13670,N_13277,N_13446);
nand U13671 (N_13671,N_13476,N_13428);
nand U13672 (N_13672,N_13351,N_13338);
or U13673 (N_13673,N_13333,N_13257);
or U13674 (N_13674,N_13369,N_13318);
or U13675 (N_13675,N_13342,N_13440);
nor U13676 (N_13676,N_13382,N_13369);
and U13677 (N_13677,N_13254,N_13352);
or U13678 (N_13678,N_13381,N_13360);
and U13679 (N_13679,N_13473,N_13280);
and U13680 (N_13680,N_13431,N_13282);
or U13681 (N_13681,N_13390,N_13453);
nor U13682 (N_13682,N_13298,N_13252);
nor U13683 (N_13683,N_13305,N_13494);
nand U13684 (N_13684,N_13398,N_13303);
or U13685 (N_13685,N_13338,N_13266);
nand U13686 (N_13686,N_13461,N_13416);
nor U13687 (N_13687,N_13489,N_13296);
nor U13688 (N_13688,N_13409,N_13394);
nor U13689 (N_13689,N_13333,N_13384);
nor U13690 (N_13690,N_13308,N_13491);
and U13691 (N_13691,N_13333,N_13450);
or U13692 (N_13692,N_13369,N_13485);
and U13693 (N_13693,N_13286,N_13437);
nor U13694 (N_13694,N_13345,N_13410);
nor U13695 (N_13695,N_13363,N_13473);
nor U13696 (N_13696,N_13464,N_13313);
nand U13697 (N_13697,N_13310,N_13421);
and U13698 (N_13698,N_13369,N_13268);
nand U13699 (N_13699,N_13410,N_13295);
nand U13700 (N_13700,N_13407,N_13388);
nor U13701 (N_13701,N_13290,N_13489);
or U13702 (N_13702,N_13275,N_13289);
nand U13703 (N_13703,N_13336,N_13388);
or U13704 (N_13704,N_13354,N_13305);
and U13705 (N_13705,N_13380,N_13406);
or U13706 (N_13706,N_13363,N_13353);
and U13707 (N_13707,N_13276,N_13497);
nand U13708 (N_13708,N_13385,N_13303);
or U13709 (N_13709,N_13403,N_13491);
nor U13710 (N_13710,N_13401,N_13462);
and U13711 (N_13711,N_13472,N_13454);
and U13712 (N_13712,N_13358,N_13405);
nor U13713 (N_13713,N_13337,N_13453);
and U13714 (N_13714,N_13276,N_13298);
xnor U13715 (N_13715,N_13357,N_13305);
and U13716 (N_13716,N_13258,N_13497);
nand U13717 (N_13717,N_13455,N_13394);
nand U13718 (N_13718,N_13372,N_13417);
and U13719 (N_13719,N_13498,N_13251);
or U13720 (N_13720,N_13318,N_13475);
nand U13721 (N_13721,N_13350,N_13474);
nor U13722 (N_13722,N_13403,N_13454);
nand U13723 (N_13723,N_13394,N_13463);
nand U13724 (N_13724,N_13328,N_13396);
and U13725 (N_13725,N_13447,N_13420);
nor U13726 (N_13726,N_13434,N_13407);
nor U13727 (N_13727,N_13356,N_13279);
and U13728 (N_13728,N_13270,N_13484);
or U13729 (N_13729,N_13367,N_13393);
nand U13730 (N_13730,N_13372,N_13311);
nor U13731 (N_13731,N_13297,N_13323);
or U13732 (N_13732,N_13319,N_13330);
or U13733 (N_13733,N_13435,N_13468);
nor U13734 (N_13734,N_13252,N_13344);
nor U13735 (N_13735,N_13283,N_13282);
and U13736 (N_13736,N_13458,N_13470);
nand U13737 (N_13737,N_13482,N_13454);
or U13738 (N_13738,N_13297,N_13332);
nor U13739 (N_13739,N_13465,N_13497);
nor U13740 (N_13740,N_13285,N_13287);
or U13741 (N_13741,N_13433,N_13332);
nand U13742 (N_13742,N_13351,N_13413);
and U13743 (N_13743,N_13390,N_13263);
nand U13744 (N_13744,N_13267,N_13352);
nand U13745 (N_13745,N_13432,N_13465);
nand U13746 (N_13746,N_13403,N_13411);
nor U13747 (N_13747,N_13264,N_13259);
and U13748 (N_13748,N_13297,N_13400);
and U13749 (N_13749,N_13263,N_13456);
nor U13750 (N_13750,N_13517,N_13562);
or U13751 (N_13751,N_13534,N_13577);
xnor U13752 (N_13752,N_13741,N_13656);
and U13753 (N_13753,N_13550,N_13711);
nand U13754 (N_13754,N_13669,N_13571);
nor U13755 (N_13755,N_13526,N_13692);
and U13756 (N_13756,N_13608,N_13716);
nor U13757 (N_13757,N_13717,N_13603);
nand U13758 (N_13758,N_13681,N_13593);
nor U13759 (N_13759,N_13589,N_13732);
nor U13760 (N_13760,N_13743,N_13582);
or U13761 (N_13761,N_13502,N_13702);
nand U13762 (N_13762,N_13590,N_13715);
or U13763 (N_13763,N_13504,N_13503);
nor U13764 (N_13764,N_13720,N_13726);
nand U13765 (N_13765,N_13630,N_13733);
nand U13766 (N_13766,N_13606,N_13611);
or U13767 (N_13767,N_13700,N_13668);
nor U13768 (N_13768,N_13614,N_13609);
nand U13769 (N_13769,N_13632,N_13535);
nand U13770 (N_13770,N_13547,N_13557);
nor U13771 (N_13771,N_13687,N_13554);
nor U13772 (N_13772,N_13588,N_13610);
nor U13773 (N_13773,N_13706,N_13636);
or U13774 (N_13774,N_13500,N_13725);
nand U13775 (N_13775,N_13604,N_13602);
nand U13776 (N_13776,N_13713,N_13703);
nor U13777 (N_13777,N_13727,N_13506);
or U13778 (N_13778,N_13701,N_13651);
nand U13779 (N_13779,N_13634,N_13528);
or U13780 (N_13780,N_13661,N_13573);
nor U13781 (N_13781,N_13745,N_13530);
nand U13782 (N_13782,N_13657,N_13537);
or U13783 (N_13783,N_13637,N_13655);
or U13784 (N_13784,N_13639,N_13540);
nand U13785 (N_13785,N_13561,N_13564);
and U13786 (N_13786,N_13719,N_13551);
or U13787 (N_13787,N_13680,N_13635);
nand U13788 (N_13788,N_13516,N_13621);
or U13789 (N_13789,N_13677,N_13746);
or U13790 (N_13790,N_13568,N_13638);
and U13791 (N_13791,N_13524,N_13660);
nor U13792 (N_13792,N_13599,N_13652);
nor U13793 (N_13793,N_13605,N_13553);
nor U13794 (N_13794,N_13645,N_13539);
nand U13795 (N_13795,N_13744,N_13617);
or U13796 (N_13796,N_13514,N_13714);
or U13797 (N_13797,N_13730,N_13559);
or U13798 (N_13798,N_13649,N_13616);
nand U13799 (N_13799,N_13710,N_13529);
nand U13800 (N_13800,N_13523,N_13722);
and U13801 (N_13801,N_13654,N_13736);
nand U13802 (N_13802,N_13664,N_13576);
or U13803 (N_13803,N_13674,N_13709);
or U13804 (N_13804,N_13629,N_13527);
nor U13805 (N_13805,N_13563,N_13574);
or U13806 (N_13806,N_13671,N_13558);
and U13807 (N_13807,N_13676,N_13545);
nor U13808 (N_13808,N_13643,N_13749);
or U13809 (N_13809,N_13640,N_13572);
nor U13810 (N_13810,N_13531,N_13625);
or U13811 (N_13811,N_13532,N_13644);
nand U13812 (N_13812,N_13646,N_13696);
nor U13813 (N_13813,N_13522,N_13658);
nor U13814 (N_13814,N_13662,N_13521);
and U13815 (N_13815,N_13721,N_13596);
nand U13816 (N_13816,N_13670,N_13525);
nand U13817 (N_13817,N_13509,N_13556);
xor U13818 (N_13818,N_13748,N_13631);
and U13819 (N_13819,N_13704,N_13742);
or U13820 (N_13820,N_13507,N_13648);
and U13821 (N_13821,N_13685,N_13597);
or U13822 (N_13822,N_13724,N_13583);
nor U13823 (N_13823,N_13723,N_13698);
and U13824 (N_13824,N_13737,N_13689);
nand U13825 (N_13825,N_13544,N_13735);
nor U13826 (N_13826,N_13581,N_13512);
and U13827 (N_13827,N_13653,N_13555);
or U13828 (N_13828,N_13728,N_13712);
xnor U13829 (N_13829,N_13641,N_13618);
or U13830 (N_13830,N_13738,N_13549);
nor U13831 (N_13831,N_13731,N_13739);
or U13832 (N_13832,N_13515,N_13501);
and U13833 (N_13833,N_13686,N_13705);
or U13834 (N_13834,N_13533,N_13683);
or U13835 (N_13835,N_13591,N_13607);
and U13836 (N_13836,N_13666,N_13682);
or U13837 (N_13837,N_13647,N_13695);
or U13838 (N_13838,N_13729,N_13595);
nor U13839 (N_13839,N_13626,N_13565);
or U13840 (N_13840,N_13575,N_13569);
and U13841 (N_13841,N_13587,N_13594);
nand U13842 (N_13842,N_13598,N_13675);
nand U13843 (N_13843,N_13708,N_13672);
and U13844 (N_13844,N_13659,N_13688);
and U13845 (N_13845,N_13718,N_13633);
nand U13846 (N_13846,N_13543,N_13536);
xor U13847 (N_13847,N_13546,N_13673);
nand U13848 (N_13848,N_13665,N_13518);
or U13849 (N_13849,N_13627,N_13579);
nor U13850 (N_13850,N_13628,N_13570);
and U13851 (N_13851,N_13505,N_13585);
and U13852 (N_13852,N_13511,N_13667);
and U13853 (N_13853,N_13623,N_13694);
and U13854 (N_13854,N_13693,N_13678);
nand U13855 (N_13855,N_13578,N_13584);
nor U13856 (N_13856,N_13734,N_13520);
nor U13857 (N_13857,N_13679,N_13508);
or U13858 (N_13858,N_13684,N_13707);
and U13859 (N_13859,N_13615,N_13642);
or U13860 (N_13860,N_13566,N_13560);
and U13861 (N_13861,N_13510,N_13624);
and U13862 (N_13862,N_13548,N_13690);
or U13863 (N_13863,N_13552,N_13542);
nand U13864 (N_13864,N_13612,N_13622);
and U13865 (N_13865,N_13513,N_13519);
nand U13866 (N_13866,N_13747,N_13740);
or U13867 (N_13867,N_13600,N_13691);
nor U13868 (N_13868,N_13580,N_13567);
nand U13869 (N_13869,N_13663,N_13586);
and U13870 (N_13870,N_13650,N_13592);
or U13871 (N_13871,N_13620,N_13697);
nand U13872 (N_13872,N_13601,N_13541);
and U13873 (N_13873,N_13619,N_13699);
xor U13874 (N_13874,N_13613,N_13538);
or U13875 (N_13875,N_13626,N_13687);
and U13876 (N_13876,N_13576,N_13710);
and U13877 (N_13877,N_13712,N_13708);
nor U13878 (N_13878,N_13632,N_13666);
or U13879 (N_13879,N_13513,N_13683);
and U13880 (N_13880,N_13626,N_13707);
nor U13881 (N_13881,N_13521,N_13612);
or U13882 (N_13882,N_13530,N_13579);
nor U13883 (N_13883,N_13576,N_13572);
nor U13884 (N_13884,N_13741,N_13676);
nor U13885 (N_13885,N_13542,N_13712);
nor U13886 (N_13886,N_13580,N_13680);
nor U13887 (N_13887,N_13588,N_13532);
nand U13888 (N_13888,N_13594,N_13624);
or U13889 (N_13889,N_13603,N_13616);
or U13890 (N_13890,N_13514,N_13716);
nand U13891 (N_13891,N_13518,N_13558);
xnor U13892 (N_13892,N_13631,N_13517);
nand U13893 (N_13893,N_13594,N_13504);
and U13894 (N_13894,N_13669,N_13683);
and U13895 (N_13895,N_13646,N_13531);
or U13896 (N_13896,N_13652,N_13738);
nor U13897 (N_13897,N_13512,N_13566);
or U13898 (N_13898,N_13708,N_13533);
nor U13899 (N_13899,N_13542,N_13555);
nand U13900 (N_13900,N_13635,N_13583);
and U13901 (N_13901,N_13694,N_13655);
and U13902 (N_13902,N_13722,N_13637);
or U13903 (N_13903,N_13627,N_13547);
nor U13904 (N_13904,N_13658,N_13662);
and U13905 (N_13905,N_13594,N_13540);
or U13906 (N_13906,N_13618,N_13546);
or U13907 (N_13907,N_13533,N_13572);
nand U13908 (N_13908,N_13605,N_13734);
and U13909 (N_13909,N_13636,N_13736);
nand U13910 (N_13910,N_13568,N_13689);
nor U13911 (N_13911,N_13714,N_13566);
and U13912 (N_13912,N_13554,N_13607);
nor U13913 (N_13913,N_13633,N_13594);
or U13914 (N_13914,N_13594,N_13640);
and U13915 (N_13915,N_13648,N_13577);
or U13916 (N_13916,N_13714,N_13610);
nand U13917 (N_13917,N_13716,N_13567);
xor U13918 (N_13918,N_13561,N_13698);
and U13919 (N_13919,N_13690,N_13508);
nand U13920 (N_13920,N_13686,N_13536);
and U13921 (N_13921,N_13620,N_13635);
nand U13922 (N_13922,N_13576,N_13684);
and U13923 (N_13923,N_13745,N_13650);
and U13924 (N_13924,N_13596,N_13623);
xnor U13925 (N_13925,N_13689,N_13671);
or U13926 (N_13926,N_13689,N_13629);
or U13927 (N_13927,N_13625,N_13502);
or U13928 (N_13928,N_13588,N_13635);
nor U13929 (N_13929,N_13667,N_13709);
nor U13930 (N_13930,N_13683,N_13510);
nor U13931 (N_13931,N_13731,N_13512);
or U13932 (N_13932,N_13666,N_13670);
nor U13933 (N_13933,N_13533,N_13613);
nor U13934 (N_13934,N_13670,N_13703);
or U13935 (N_13935,N_13540,N_13598);
or U13936 (N_13936,N_13589,N_13708);
or U13937 (N_13937,N_13653,N_13725);
and U13938 (N_13938,N_13683,N_13719);
nor U13939 (N_13939,N_13567,N_13708);
and U13940 (N_13940,N_13632,N_13653);
nor U13941 (N_13941,N_13604,N_13586);
nand U13942 (N_13942,N_13689,N_13682);
nor U13943 (N_13943,N_13585,N_13547);
and U13944 (N_13944,N_13583,N_13596);
and U13945 (N_13945,N_13600,N_13743);
or U13946 (N_13946,N_13710,N_13663);
and U13947 (N_13947,N_13640,N_13624);
or U13948 (N_13948,N_13742,N_13514);
nor U13949 (N_13949,N_13655,N_13565);
nand U13950 (N_13950,N_13518,N_13590);
or U13951 (N_13951,N_13698,N_13677);
or U13952 (N_13952,N_13696,N_13687);
nand U13953 (N_13953,N_13654,N_13534);
xor U13954 (N_13954,N_13653,N_13633);
and U13955 (N_13955,N_13548,N_13536);
nand U13956 (N_13956,N_13719,N_13665);
or U13957 (N_13957,N_13563,N_13539);
nor U13958 (N_13958,N_13676,N_13719);
or U13959 (N_13959,N_13654,N_13625);
or U13960 (N_13960,N_13586,N_13565);
and U13961 (N_13961,N_13631,N_13553);
nand U13962 (N_13962,N_13591,N_13577);
or U13963 (N_13963,N_13682,N_13704);
and U13964 (N_13964,N_13665,N_13534);
nand U13965 (N_13965,N_13728,N_13691);
or U13966 (N_13966,N_13652,N_13598);
nor U13967 (N_13967,N_13654,N_13744);
and U13968 (N_13968,N_13595,N_13670);
or U13969 (N_13969,N_13530,N_13554);
and U13970 (N_13970,N_13536,N_13505);
or U13971 (N_13971,N_13643,N_13584);
xnor U13972 (N_13972,N_13574,N_13586);
and U13973 (N_13973,N_13672,N_13717);
xor U13974 (N_13974,N_13651,N_13543);
and U13975 (N_13975,N_13698,N_13706);
or U13976 (N_13976,N_13712,N_13506);
and U13977 (N_13977,N_13505,N_13684);
nor U13978 (N_13978,N_13689,N_13742);
nand U13979 (N_13979,N_13729,N_13724);
nor U13980 (N_13980,N_13624,N_13595);
or U13981 (N_13981,N_13601,N_13622);
and U13982 (N_13982,N_13629,N_13697);
and U13983 (N_13983,N_13534,N_13712);
nor U13984 (N_13984,N_13719,N_13550);
nor U13985 (N_13985,N_13640,N_13535);
xor U13986 (N_13986,N_13584,N_13503);
or U13987 (N_13987,N_13646,N_13612);
or U13988 (N_13988,N_13596,N_13579);
and U13989 (N_13989,N_13630,N_13623);
and U13990 (N_13990,N_13592,N_13560);
nand U13991 (N_13991,N_13614,N_13591);
nor U13992 (N_13992,N_13691,N_13684);
and U13993 (N_13993,N_13584,N_13690);
nor U13994 (N_13994,N_13622,N_13663);
nand U13995 (N_13995,N_13648,N_13690);
or U13996 (N_13996,N_13725,N_13746);
nor U13997 (N_13997,N_13550,N_13653);
and U13998 (N_13998,N_13539,N_13680);
nor U13999 (N_13999,N_13598,N_13746);
nor U14000 (N_14000,N_13917,N_13777);
and U14001 (N_14001,N_13822,N_13954);
or U14002 (N_14002,N_13758,N_13888);
and U14003 (N_14003,N_13850,N_13967);
xor U14004 (N_14004,N_13936,N_13997);
and U14005 (N_14005,N_13854,N_13893);
nand U14006 (N_14006,N_13763,N_13750);
nor U14007 (N_14007,N_13820,N_13921);
or U14008 (N_14008,N_13867,N_13819);
and U14009 (N_14009,N_13938,N_13885);
nor U14010 (N_14010,N_13895,N_13995);
nor U14011 (N_14011,N_13754,N_13845);
nor U14012 (N_14012,N_13944,N_13767);
nand U14013 (N_14013,N_13875,N_13914);
nor U14014 (N_14014,N_13870,N_13816);
nor U14015 (N_14015,N_13828,N_13860);
or U14016 (N_14016,N_13836,N_13975);
and U14017 (N_14017,N_13915,N_13918);
or U14018 (N_14018,N_13968,N_13868);
nand U14019 (N_14019,N_13825,N_13775);
and U14020 (N_14020,N_13843,N_13942);
nor U14021 (N_14021,N_13841,N_13873);
and U14022 (N_14022,N_13953,N_13956);
or U14023 (N_14023,N_13978,N_13891);
nand U14024 (N_14024,N_13827,N_13826);
or U14025 (N_14025,N_13952,N_13751);
nand U14026 (N_14026,N_13814,N_13821);
or U14027 (N_14027,N_13989,N_13964);
and U14028 (N_14028,N_13797,N_13785);
and U14029 (N_14029,N_13990,N_13906);
nand U14030 (N_14030,N_13815,N_13838);
nor U14031 (N_14031,N_13974,N_13972);
nand U14032 (N_14032,N_13920,N_13892);
nand U14033 (N_14033,N_13999,N_13880);
nor U14034 (N_14034,N_13852,N_13963);
nand U14035 (N_14035,N_13966,N_13903);
xnor U14036 (N_14036,N_13858,N_13837);
nand U14037 (N_14037,N_13948,N_13804);
nand U14038 (N_14038,N_13946,N_13987);
nand U14039 (N_14039,N_13890,N_13960);
nand U14040 (N_14040,N_13807,N_13800);
nor U14041 (N_14041,N_13761,N_13796);
and U14042 (N_14042,N_13752,N_13872);
or U14043 (N_14043,N_13950,N_13992);
nand U14044 (N_14044,N_13774,N_13764);
or U14045 (N_14045,N_13897,N_13865);
nor U14046 (N_14046,N_13790,N_13896);
nor U14047 (N_14047,N_13901,N_13848);
and U14048 (N_14048,N_13983,N_13871);
and U14049 (N_14049,N_13969,N_13817);
or U14050 (N_14050,N_13940,N_13928);
nor U14051 (N_14051,N_13760,N_13788);
and U14052 (N_14052,N_13961,N_13991);
or U14053 (N_14053,N_13929,N_13937);
and U14054 (N_14054,N_13886,N_13834);
xnor U14055 (N_14055,N_13894,N_13830);
nor U14056 (N_14056,N_13916,N_13923);
nand U14057 (N_14057,N_13794,N_13881);
or U14058 (N_14058,N_13857,N_13793);
or U14059 (N_14059,N_13861,N_13769);
nand U14060 (N_14060,N_13933,N_13932);
or U14061 (N_14061,N_13980,N_13776);
or U14062 (N_14062,N_13832,N_13811);
and U14063 (N_14063,N_13787,N_13986);
or U14064 (N_14064,N_13943,N_13922);
xor U14065 (N_14065,N_13981,N_13869);
or U14066 (N_14066,N_13802,N_13905);
nand U14067 (N_14067,N_13846,N_13898);
nand U14068 (N_14068,N_13965,N_13770);
and U14069 (N_14069,N_13782,N_13951);
nor U14070 (N_14070,N_13862,N_13911);
or U14071 (N_14071,N_13959,N_13889);
nor U14072 (N_14072,N_13855,N_13919);
and U14073 (N_14073,N_13924,N_13884);
and U14074 (N_14074,N_13808,N_13945);
or U14075 (N_14075,N_13973,N_13840);
nor U14076 (N_14076,N_13877,N_13783);
or U14077 (N_14077,N_13810,N_13979);
and U14078 (N_14078,N_13912,N_13909);
or U14079 (N_14079,N_13801,N_13910);
nor U14080 (N_14080,N_13795,N_13806);
nor U14081 (N_14081,N_13900,N_13988);
xnor U14082 (N_14082,N_13759,N_13756);
xnor U14083 (N_14083,N_13994,N_13931);
nand U14084 (N_14084,N_13798,N_13913);
and U14085 (N_14085,N_13935,N_13957);
and U14086 (N_14086,N_13934,N_13899);
nor U14087 (N_14087,N_13939,N_13851);
xnor U14088 (N_14088,N_13823,N_13907);
nor U14089 (N_14089,N_13949,N_13925);
nor U14090 (N_14090,N_13813,N_13998);
or U14091 (N_14091,N_13818,N_13766);
and U14092 (N_14092,N_13778,N_13874);
nand U14093 (N_14093,N_13926,N_13864);
or U14094 (N_14094,N_13853,N_13955);
nor U14095 (N_14095,N_13962,N_13835);
or U14096 (N_14096,N_13958,N_13996);
and U14097 (N_14097,N_13984,N_13771);
or U14098 (N_14098,N_13876,N_13930);
or U14099 (N_14099,N_13773,N_13781);
nor U14100 (N_14100,N_13970,N_13849);
and U14101 (N_14101,N_13866,N_13847);
nand U14102 (N_14102,N_13863,N_13762);
xnor U14103 (N_14103,N_13844,N_13784);
nand U14104 (N_14104,N_13799,N_13971);
nor U14105 (N_14105,N_13789,N_13809);
or U14106 (N_14106,N_13902,N_13755);
and U14107 (N_14107,N_13882,N_13879);
nor U14108 (N_14108,N_13887,N_13883);
nand U14109 (N_14109,N_13856,N_13985);
nand U14110 (N_14110,N_13839,N_13792);
and U14111 (N_14111,N_13904,N_13982);
nor U14112 (N_14112,N_13993,N_13908);
and U14113 (N_14113,N_13927,N_13947);
xor U14114 (N_14114,N_13791,N_13786);
nor U14115 (N_14115,N_13803,N_13878);
and U14116 (N_14116,N_13768,N_13977);
or U14117 (N_14117,N_13765,N_13829);
or U14118 (N_14118,N_13753,N_13757);
and U14119 (N_14119,N_13772,N_13941);
nand U14120 (N_14120,N_13824,N_13859);
nand U14121 (N_14121,N_13780,N_13833);
nand U14122 (N_14122,N_13779,N_13812);
and U14123 (N_14123,N_13842,N_13805);
nor U14124 (N_14124,N_13976,N_13831);
or U14125 (N_14125,N_13935,N_13867);
and U14126 (N_14126,N_13781,N_13868);
nor U14127 (N_14127,N_13823,N_13837);
or U14128 (N_14128,N_13810,N_13858);
nand U14129 (N_14129,N_13750,N_13946);
or U14130 (N_14130,N_13782,N_13967);
or U14131 (N_14131,N_13970,N_13824);
and U14132 (N_14132,N_13987,N_13911);
nor U14133 (N_14133,N_13779,N_13772);
nand U14134 (N_14134,N_13966,N_13764);
and U14135 (N_14135,N_13797,N_13766);
nand U14136 (N_14136,N_13793,N_13862);
or U14137 (N_14137,N_13765,N_13773);
nor U14138 (N_14138,N_13863,N_13797);
or U14139 (N_14139,N_13770,N_13827);
or U14140 (N_14140,N_13815,N_13846);
or U14141 (N_14141,N_13901,N_13906);
or U14142 (N_14142,N_13844,N_13972);
xnor U14143 (N_14143,N_13755,N_13938);
or U14144 (N_14144,N_13768,N_13846);
and U14145 (N_14145,N_13965,N_13862);
nor U14146 (N_14146,N_13950,N_13771);
nand U14147 (N_14147,N_13766,N_13847);
nor U14148 (N_14148,N_13798,N_13901);
and U14149 (N_14149,N_13769,N_13913);
nor U14150 (N_14150,N_13835,N_13905);
and U14151 (N_14151,N_13760,N_13857);
nor U14152 (N_14152,N_13751,N_13985);
nand U14153 (N_14153,N_13984,N_13825);
or U14154 (N_14154,N_13951,N_13777);
nor U14155 (N_14155,N_13913,N_13891);
nor U14156 (N_14156,N_13992,N_13816);
or U14157 (N_14157,N_13789,N_13942);
or U14158 (N_14158,N_13808,N_13868);
or U14159 (N_14159,N_13974,N_13932);
nor U14160 (N_14160,N_13953,N_13812);
nand U14161 (N_14161,N_13812,N_13776);
xnor U14162 (N_14162,N_13827,N_13858);
nor U14163 (N_14163,N_13949,N_13940);
nand U14164 (N_14164,N_13963,N_13802);
or U14165 (N_14165,N_13903,N_13885);
or U14166 (N_14166,N_13880,N_13922);
nor U14167 (N_14167,N_13941,N_13971);
or U14168 (N_14168,N_13791,N_13977);
or U14169 (N_14169,N_13836,N_13944);
and U14170 (N_14170,N_13785,N_13802);
nor U14171 (N_14171,N_13755,N_13990);
and U14172 (N_14172,N_13938,N_13774);
xnor U14173 (N_14173,N_13923,N_13857);
nand U14174 (N_14174,N_13859,N_13801);
nand U14175 (N_14175,N_13914,N_13765);
and U14176 (N_14176,N_13978,N_13848);
nand U14177 (N_14177,N_13814,N_13773);
and U14178 (N_14178,N_13846,N_13991);
xor U14179 (N_14179,N_13878,N_13754);
nand U14180 (N_14180,N_13964,N_13951);
or U14181 (N_14181,N_13999,N_13922);
and U14182 (N_14182,N_13998,N_13960);
or U14183 (N_14183,N_13762,N_13963);
and U14184 (N_14184,N_13892,N_13982);
or U14185 (N_14185,N_13913,N_13772);
nor U14186 (N_14186,N_13987,N_13898);
nand U14187 (N_14187,N_13929,N_13774);
or U14188 (N_14188,N_13835,N_13792);
nor U14189 (N_14189,N_13881,N_13889);
nand U14190 (N_14190,N_13804,N_13868);
nor U14191 (N_14191,N_13754,N_13902);
or U14192 (N_14192,N_13968,N_13953);
or U14193 (N_14193,N_13793,N_13785);
nand U14194 (N_14194,N_13943,N_13751);
nor U14195 (N_14195,N_13767,N_13904);
and U14196 (N_14196,N_13911,N_13804);
or U14197 (N_14197,N_13998,N_13797);
or U14198 (N_14198,N_13876,N_13827);
nand U14199 (N_14199,N_13797,N_13853);
or U14200 (N_14200,N_13767,N_13858);
nand U14201 (N_14201,N_13756,N_13864);
nor U14202 (N_14202,N_13885,N_13825);
and U14203 (N_14203,N_13820,N_13755);
nor U14204 (N_14204,N_13828,N_13908);
xnor U14205 (N_14205,N_13959,N_13928);
nor U14206 (N_14206,N_13797,N_13955);
or U14207 (N_14207,N_13999,N_13868);
nor U14208 (N_14208,N_13812,N_13859);
or U14209 (N_14209,N_13944,N_13911);
nand U14210 (N_14210,N_13883,N_13866);
nor U14211 (N_14211,N_13875,N_13769);
and U14212 (N_14212,N_13960,N_13775);
or U14213 (N_14213,N_13846,N_13781);
nor U14214 (N_14214,N_13834,N_13775);
nand U14215 (N_14215,N_13978,N_13821);
and U14216 (N_14216,N_13893,N_13975);
nor U14217 (N_14217,N_13871,N_13872);
nor U14218 (N_14218,N_13909,N_13811);
and U14219 (N_14219,N_13866,N_13823);
or U14220 (N_14220,N_13904,N_13863);
or U14221 (N_14221,N_13973,N_13804);
nor U14222 (N_14222,N_13779,N_13791);
nor U14223 (N_14223,N_13790,N_13761);
and U14224 (N_14224,N_13887,N_13893);
or U14225 (N_14225,N_13906,N_13843);
nand U14226 (N_14226,N_13963,N_13844);
nor U14227 (N_14227,N_13992,N_13789);
and U14228 (N_14228,N_13800,N_13802);
nand U14229 (N_14229,N_13892,N_13843);
or U14230 (N_14230,N_13984,N_13871);
nor U14231 (N_14231,N_13799,N_13926);
nand U14232 (N_14232,N_13931,N_13841);
and U14233 (N_14233,N_13966,N_13997);
nor U14234 (N_14234,N_13832,N_13975);
nand U14235 (N_14235,N_13871,N_13752);
nand U14236 (N_14236,N_13955,N_13772);
and U14237 (N_14237,N_13793,N_13861);
xor U14238 (N_14238,N_13870,N_13756);
and U14239 (N_14239,N_13804,N_13817);
and U14240 (N_14240,N_13910,N_13762);
nand U14241 (N_14241,N_13786,N_13953);
nor U14242 (N_14242,N_13855,N_13788);
and U14243 (N_14243,N_13793,N_13753);
or U14244 (N_14244,N_13750,N_13904);
nor U14245 (N_14245,N_13772,N_13964);
nor U14246 (N_14246,N_13752,N_13933);
and U14247 (N_14247,N_13958,N_13913);
nand U14248 (N_14248,N_13812,N_13901);
nor U14249 (N_14249,N_13909,N_13843);
nor U14250 (N_14250,N_14053,N_14039);
nand U14251 (N_14251,N_14111,N_14170);
and U14252 (N_14252,N_14086,N_14114);
and U14253 (N_14253,N_14018,N_14027);
nand U14254 (N_14254,N_14178,N_14164);
nor U14255 (N_14255,N_14222,N_14213);
nor U14256 (N_14256,N_14110,N_14137);
or U14257 (N_14257,N_14005,N_14192);
xnor U14258 (N_14258,N_14097,N_14067);
and U14259 (N_14259,N_14071,N_14081);
or U14260 (N_14260,N_14020,N_14132);
nand U14261 (N_14261,N_14009,N_14203);
or U14262 (N_14262,N_14182,N_14117);
and U14263 (N_14263,N_14101,N_14022);
and U14264 (N_14264,N_14172,N_14059);
nand U14265 (N_14265,N_14198,N_14136);
and U14266 (N_14266,N_14236,N_14103);
nand U14267 (N_14267,N_14180,N_14011);
nand U14268 (N_14268,N_14133,N_14085);
or U14269 (N_14269,N_14123,N_14229);
or U14270 (N_14270,N_14091,N_14174);
or U14271 (N_14271,N_14211,N_14084);
and U14272 (N_14272,N_14181,N_14036);
and U14273 (N_14273,N_14074,N_14173);
xnor U14274 (N_14274,N_14115,N_14076);
and U14275 (N_14275,N_14077,N_14225);
nor U14276 (N_14276,N_14066,N_14208);
and U14277 (N_14277,N_14026,N_14243);
nor U14278 (N_14278,N_14245,N_14126);
nor U14279 (N_14279,N_14148,N_14043);
or U14280 (N_14280,N_14073,N_14233);
and U14281 (N_14281,N_14215,N_14099);
nor U14282 (N_14282,N_14100,N_14000);
nor U14283 (N_14283,N_14217,N_14207);
nor U14284 (N_14284,N_14201,N_14113);
and U14285 (N_14285,N_14187,N_14144);
and U14286 (N_14286,N_14184,N_14221);
nor U14287 (N_14287,N_14200,N_14216);
nor U14288 (N_14288,N_14134,N_14002);
or U14289 (N_14289,N_14210,N_14008);
or U14290 (N_14290,N_14063,N_14118);
and U14291 (N_14291,N_14241,N_14034);
and U14292 (N_14292,N_14130,N_14062);
xnor U14293 (N_14293,N_14042,N_14121);
nor U14294 (N_14294,N_14021,N_14102);
or U14295 (N_14295,N_14038,N_14035);
or U14296 (N_14296,N_14165,N_14249);
xor U14297 (N_14297,N_14028,N_14185);
and U14298 (N_14298,N_14141,N_14197);
nor U14299 (N_14299,N_14094,N_14196);
nand U14300 (N_14300,N_14017,N_14127);
or U14301 (N_14301,N_14212,N_14010);
or U14302 (N_14302,N_14228,N_14030);
nand U14303 (N_14303,N_14058,N_14041);
or U14304 (N_14304,N_14205,N_14235);
nand U14305 (N_14305,N_14007,N_14112);
nor U14306 (N_14306,N_14057,N_14119);
nand U14307 (N_14307,N_14078,N_14013);
nand U14308 (N_14308,N_14014,N_14093);
or U14309 (N_14309,N_14204,N_14029);
and U14310 (N_14310,N_14140,N_14128);
and U14311 (N_14311,N_14155,N_14048);
nor U14312 (N_14312,N_14049,N_14089);
and U14313 (N_14313,N_14044,N_14191);
nand U14314 (N_14314,N_14023,N_14056);
nand U14315 (N_14315,N_14226,N_14142);
nor U14316 (N_14316,N_14147,N_14032);
nand U14317 (N_14317,N_14146,N_14242);
nand U14318 (N_14318,N_14202,N_14001);
xnor U14319 (N_14319,N_14124,N_14068);
or U14320 (N_14320,N_14194,N_14116);
nor U14321 (N_14321,N_14156,N_14159);
and U14322 (N_14322,N_14167,N_14158);
nor U14323 (N_14323,N_14166,N_14016);
or U14324 (N_14324,N_14168,N_14154);
or U14325 (N_14325,N_14150,N_14177);
and U14326 (N_14326,N_14087,N_14193);
nand U14327 (N_14327,N_14082,N_14092);
nor U14328 (N_14328,N_14145,N_14107);
nor U14329 (N_14329,N_14033,N_14223);
nor U14330 (N_14330,N_14179,N_14139);
and U14331 (N_14331,N_14143,N_14224);
or U14332 (N_14332,N_14248,N_14230);
xnor U14333 (N_14333,N_14183,N_14120);
nand U14334 (N_14334,N_14061,N_14232);
nand U14335 (N_14335,N_14149,N_14247);
nand U14336 (N_14336,N_14135,N_14214);
nand U14337 (N_14337,N_14206,N_14045);
and U14338 (N_14338,N_14238,N_14153);
or U14339 (N_14339,N_14195,N_14070);
and U14340 (N_14340,N_14209,N_14095);
nor U14341 (N_14341,N_14060,N_14088);
and U14342 (N_14342,N_14160,N_14096);
or U14343 (N_14343,N_14175,N_14219);
nor U14344 (N_14344,N_14171,N_14227);
or U14345 (N_14345,N_14131,N_14054);
or U14346 (N_14346,N_14104,N_14239);
nand U14347 (N_14347,N_14106,N_14244);
nor U14348 (N_14348,N_14246,N_14024);
nor U14349 (N_14349,N_14090,N_14015);
nand U14350 (N_14350,N_14186,N_14072);
and U14351 (N_14351,N_14162,N_14050);
and U14352 (N_14352,N_14125,N_14188);
nor U14353 (N_14353,N_14012,N_14138);
nand U14354 (N_14354,N_14055,N_14031);
and U14355 (N_14355,N_14004,N_14163);
and U14356 (N_14356,N_14109,N_14152);
or U14357 (N_14357,N_14069,N_14079);
nor U14358 (N_14358,N_14105,N_14046);
nor U14359 (N_14359,N_14047,N_14199);
and U14360 (N_14360,N_14108,N_14129);
nand U14361 (N_14361,N_14151,N_14003);
and U14362 (N_14362,N_14122,N_14240);
or U14363 (N_14363,N_14065,N_14189);
or U14364 (N_14364,N_14220,N_14218);
nand U14365 (N_14365,N_14176,N_14075);
nor U14366 (N_14366,N_14019,N_14064);
nor U14367 (N_14367,N_14006,N_14098);
nor U14368 (N_14368,N_14157,N_14040);
and U14369 (N_14369,N_14161,N_14025);
or U14370 (N_14370,N_14237,N_14234);
and U14371 (N_14371,N_14190,N_14169);
and U14372 (N_14372,N_14080,N_14231);
nor U14373 (N_14373,N_14052,N_14037);
and U14374 (N_14374,N_14051,N_14083);
nand U14375 (N_14375,N_14055,N_14151);
and U14376 (N_14376,N_14080,N_14033);
or U14377 (N_14377,N_14100,N_14162);
nand U14378 (N_14378,N_14029,N_14087);
or U14379 (N_14379,N_14145,N_14181);
or U14380 (N_14380,N_14239,N_14081);
nor U14381 (N_14381,N_14144,N_14005);
nand U14382 (N_14382,N_14144,N_14031);
nand U14383 (N_14383,N_14158,N_14144);
nor U14384 (N_14384,N_14020,N_14110);
nor U14385 (N_14385,N_14247,N_14181);
nand U14386 (N_14386,N_14003,N_14127);
and U14387 (N_14387,N_14154,N_14190);
and U14388 (N_14388,N_14128,N_14221);
nor U14389 (N_14389,N_14027,N_14088);
and U14390 (N_14390,N_14018,N_14099);
or U14391 (N_14391,N_14134,N_14238);
and U14392 (N_14392,N_14108,N_14128);
xor U14393 (N_14393,N_14189,N_14101);
and U14394 (N_14394,N_14129,N_14097);
and U14395 (N_14395,N_14138,N_14222);
nor U14396 (N_14396,N_14050,N_14074);
xor U14397 (N_14397,N_14027,N_14195);
nand U14398 (N_14398,N_14127,N_14125);
nand U14399 (N_14399,N_14175,N_14161);
or U14400 (N_14400,N_14183,N_14105);
nand U14401 (N_14401,N_14176,N_14092);
and U14402 (N_14402,N_14111,N_14105);
or U14403 (N_14403,N_14100,N_14070);
and U14404 (N_14404,N_14246,N_14228);
nand U14405 (N_14405,N_14141,N_14177);
or U14406 (N_14406,N_14056,N_14100);
nand U14407 (N_14407,N_14159,N_14174);
nand U14408 (N_14408,N_14189,N_14248);
or U14409 (N_14409,N_14117,N_14225);
and U14410 (N_14410,N_14047,N_14192);
nor U14411 (N_14411,N_14049,N_14249);
and U14412 (N_14412,N_14017,N_14152);
nor U14413 (N_14413,N_14004,N_14043);
or U14414 (N_14414,N_14188,N_14052);
or U14415 (N_14415,N_14075,N_14057);
and U14416 (N_14416,N_14213,N_14011);
or U14417 (N_14417,N_14219,N_14115);
or U14418 (N_14418,N_14219,N_14097);
or U14419 (N_14419,N_14125,N_14197);
and U14420 (N_14420,N_14153,N_14185);
or U14421 (N_14421,N_14082,N_14157);
or U14422 (N_14422,N_14128,N_14182);
or U14423 (N_14423,N_14021,N_14222);
nand U14424 (N_14424,N_14089,N_14164);
nand U14425 (N_14425,N_14072,N_14226);
nand U14426 (N_14426,N_14188,N_14197);
and U14427 (N_14427,N_14242,N_14154);
nor U14428 (N_14428,N_14122,N_14100);
xor U14429 (N_14429,N_14167,N_14021);
nor U14430 (N_14430,N_14132,N_14094);
nor U14431 (N_14431,N_14077,N_14128);
or U14432 (N_14432,N_14107,N_14150);
xor U14433 (N_14433,N_14028,N_14205);
nand U14434 (N_14434,N_14053,N_14187);
nor U14435 (N_14435,N_14178,N_14005);
or U14436 (N_14436,N_14062,N_14091);
nand U14437 (N_14437,N_14037,N_14148);
or U14438 (N_14438,N_14215,N_14228);
nor U14439 (N_14439,N_14045,N_14220);
xor U14440 (N_14440,N_14074,N_14051);
or U14441 (N_14441,N_14200,N_14169);
or U14442 (N_14442,N_14242,N_14241);
nor U14443 (N_14443,N_14012,N_14110);
nor U14444 (N_14444,N_14132,N_14008);
or U14445 (N_14445,N_14097,N_14234);
nor U14446 (N_14446,N_14112,N_14143);
or U14447 (N_14447,N_14200,N_14125);
or U14448 (N_14448,N_14191,N_14064);
nand U14449 (N_14449,N_14217,N_14057);
or U14450 (N_14450,N_14044,N_14108);
or U14451 (N_14451,N_14094,N_14224);
and U14452 (N_14452,N_14198,N_14243);
nor U14453 (N_14453,N_14168,N_14075);
nand U14454 (N_14454,N_14169,N_14100);
and U14455 (N_14455,N_14099,N_14220);
and U14456 (N_14456,N_14138,N_14017);
nor U14457 (N_14457,N_14233,N_14039);
nand U14458 (N_14458,N_14171,N_14153);
nor U14459 (N_14459,N_14094,N_14103);
nand U14460 (N_14460,N_14223,N_14050);
nor U14461 (N_14461,N_14056,N_14155);
or U14462 (N_14462,N_14149,N_14243);
and U14463 (N_14463,N_14207,N_14066);
or U14464 (N_14464,N_14101,N_14066);
nor U14465 (N_14465,N_14204,N_14201);
xor U14466 (N_14466,N_14147,N_14201);
nor U14467 (N_14467,N_14200,N_14001);
nor U14468 (N_14468,N_14133,N_14009);
and U14469 (N_14469,N_14236,N_14084);
and U14470 (N_14470,N_14175,N_14146);
nor U14471 (N_14471,N_14209,N_14217);
or U14472 (N_14472,N_14207,N_14046);
or U14473 (N_14473,N_14101,N_14132);
and U14474 (N_14474,N_14211,N_14242);
and U14475 (N_14475,N_14212,N_14143);
and U14476 (N_14476,N_14176,N_14029);
or U14477 (N_14477,N_14086,N_14072);
nand U14478 (N_14478,N_14053,N_14116);
and U14479 (N_14479,N_14142,N_14114);
nor U14480 (N_14480,N_14123,N_14062);
nor U14481 (N_14481,N_14086,N_14183);
or U14482 (N_14482,N_14211,N_14171);
and U14483 (N_14483,N_14077,N_14181);
and U14484 (N_14484,N_14137,N_14134);
nor U14485 (N_14485,N_14055,N_14024);
or U14486 (N_14486,N_14020,N_14007);
or U14487 (N_14487,N_14049,N_14202);
or U14488 (N_14488,N_14170,N_14155);
or U14489 (N_14489,N_14138,N_14229);
and U14490 (N_14490,N_14209,N_14072);
nor U14491 (N_14491,N_14071,N_14096);
nand U14492 (N_14492,N_14105,N_14159);
and U14493 (N_14493,N_14059,N_14129);
or U14494 (N_14494,N_14165,N_14123);
and U14495 (N_14495,N_14028,N_14114);
nand U14496 (N_14496,N_14214,N_14075);
nor U14497 (N_14497,N_14056,N_14181);
or U14498 (N_14498,N_14070,N_14165);
nor U14499 (N_14499,N_14153,N_14239);
or U14500 (N_14500,N_14336,N_14459);
nor U14501 (N_14501,N_14439,N_14297);
and U14502 (N_14502,N_14364,N_14251);
xnor U14503 (N_14503,N_14470,N_14465);
or U14504 (N_14504,N_14306,N_14444);
or U14505 (N_14505,N_14423,N_14256);
and U14506 (N_14506,N_14476,N_14345);
nand U14507 (N_14507,N_14485,N_14283);
nor U14508 (N_14508,N_14281,N_14483);
and U14509 (N_14509,N_14471,N_14494);
nand U14510 (N_14510,N_14310,N_14273);
nor U14511 (N_14511,N_14408,N_14428);
and U14512 (N_14512,N_14398,N_14264);
and U14513 (N_14513,N_14395,N_14429);
nor U14514 (N_14514,N_14302,N_14496);
or U14515 (N_14515,N_14269,N_14323);
nand U14516 (N_14516,N_14315,N_14427);
or U14517 (N_14517,N_14299,N_14413);
and U14518 (N_14518,N_14348,N_14295);
or U14519 (N_14519,N_14335,N_14451);
nand U14520 (N_14520,N_14446,N_14414);
nor U14521 (N_14521,N_14378,N_14409);
and U14522 (N_14522,N_14389,N_14447);
nand U14523 (N_14523,N_14321,N_14394);
or U14524 (N_14524,N_14291,N_14479);
nand U14525 (N_14525,N_14290,N_14346);
nand U14526 (N_14526,N_14337,N_14260);
nand U14527 (N_14527,N_14438,N_14420);
nand U14528 (N_14528,N_14328,N_14426);
nand U14529 (N_14529,N_14294,N_14493);
and U14530 (N_14530,N_14331,N_14387);
or U14531 (N_14531,N_14388,N_14376);
or U14532 (N_14532,N_14275,N_14435);
or U14533 (N_14533,N_14473,N_14432);
and U14534 (N_14534,N_14357,N_14262);
nor U14535 (N_14535,N_14437,N_14367);
or U14536 (N_14536,N_14274,N_14421);
and U14537 (N_14537,N_14332,N_14416);
or U14538 (N_14538,N_14280,N_14448);
nor U14539 (N_14539,N_14440,N_14296);
and U14540 (N_14540,N_14324,N_14466);
or U14541 (N_14541,N_14415,N_14482);
nor U14542 (N_14542,N_14286,N_14338);
or U14543 (N_14543,N_14284,N_14434);
or U14544 (N_14544,N_14361,N_14392);
and U14545 (N_14545,N_14405,N_14450);
and U14546 (N_14546,N_14375,N_14452);
nor U14547 (N_14547,N_14425,N_14343);
and U14548 (N_14548,N_14311,N_14277);
nand U14549 (N_14549,N_14354,N_14467);
nand U14550 (N_14550,N_14288,N_14441);
and U14551 (N_14551,N_14443,N_14353);
nor U14552 (N_14552,N_14430,N_14462);
nand U14553 (N_14553,N_14268,N_14265);
and U14554 (N_14554,N_14350,N_14454);
or U14555 (N_14555,N_14363,N_14362);
or U14556 (N_14556,N_14333,N_14270);
nor U14557 (N_14557,N_14317,N_14271);
or U14558 (N_14558,N_14498,N_14418);
nor U14559 (N_14559,N_14330,N_14318);
or U14560 (N_14560,N_14347,N_14307);
nor U14561 (N_14561,N_14381,N_14356);
nand U14562 (N_14562,N_14329,N_14272);
and U14563 (N_14563,N_14486,N_14340);
xor U14564 (N_14564,N_14368,N_14313);
or U14565 (N_14565,N_14478,N_14391);
nand U14566 (N_14566,N_14492,N_14480);
and U14567 (N_14567,N_14301,N_14488);
or U14568 (N_14568,N_14379,N_14461);
and U14569 (N_14569,N_14431,N_14453);
and U14570 (N_14570,N_14266,N_14285);
nand U14571 (N_14571,N_14474,N_14316);
nand U14572 (N_14572,N_14487,N_14386);
or U14573 (N_14573,N_14358,N_14255);
nand U14574 (N_14574,N_14499,N_14349);
nand U14575 (N_14575,N_14404,N_14322);
or U14576 (N_14576,N_14497,N_14419);
or U14577 (N_14577,N_14351,N_14254);
nand U14578 (N_14578,N_14460,N_14355);
and U14579 (N_14579,N_14339,N_14372);
and U14580 (N_14580,N_14411,N_14393);
nand U14581 (N_14581,N_14373,N_14402);
nand U14582 (N_14582,N_14359,N_14469);
and U14583 (N_14583,N_14257,N_14449);
or U14584 (N_14584,N_14481,N_14377);
nor U14585 (N_14585,N_14309,N_14366);
nand U14586 (N_14586,N_14397,N_14489);
nor U14587 (N_14587,N_14384,N_14458);
and U14588 (N_14588,N_14406,N_14282);
or U14589 (N_14589,N_14495,N_14300);
nor U14590 (N_14590,N_14319,N_14289);
and U14591 (N_14591,N_14491,N_14303);
and U14592 (N_14592,N_14436,N_14400);
nor U14593 (N_14593,N_14325,N_14334);
nand U14594 (N_14594,N_14385,N_14445);
nand U14595 (N_14595,N_14417,N_14250);
nand U14596 (N_14596,N_14369,N_14371);
and U14597 (N_14597,N_14396,N_14308);
and U14598 (N_14598,N_14433,N_14292);
nor U14599 (N_14599,N_14344,N_14442);
nor U14600 (N_14600,N_14463,N_14424);
and U14601 (N_14601,N_14305,N_14468);
nand U14602 (N_14602,N_14365,N_14326);
and U14603 (N_14603,N_14457,N_14276);
and U14604 (N_14604,N_14383,N_14312);
or U14605 (N_14605,N_14382,N_14380);
and U14606 (N_14606,N_14252,N_14267);
nor U14607 (N_14607,N_14253,N_14374);
or U14608 (N_14608,N_14293,N_14490);
nor U14609 (N_14609,N_14279,N_14263);
xnor U14610 (N_14610,N_14352,N_14314);
or U14611 (N_14611,N_14261,N_14403);
and U14612 (N_14612,N_14399,N_14304);
or U14613 (N_14613,N_14320,N_14259);
and U14614 (N_14614,N_14370,N_14410);
and U14615 (N_14615,N_14456,N_14278);
and U14616 (N_14616,N_14401,N_14475);
nand U14617 (N_14617,N_14477,N_14422);
and U14618 (N_14618,N_14341,N_14484);
nand U14619 (N_14619,N_14407,N_14455);
and U14620 (N_14620,N_14464,N_14287);
nand U14621 (N_14621,N_14412,N_14390);
or U14622 (N_14622,N_14258,N_14327);
and U14623 (N_14623,N_14360,N_14298);
nor U14624 (N_14624,N_14342,N_14472);
and U14625 (N_14625,N_14404,N_14295);
nand U14626 (N_14626,N_14431,N_14467);
and U14627 (N_14627,N_14349,N_14351);
nand U14628 (N_14628,N_14349,N_14379);
or U14629 (N_14629,N_14251,N_14489);
and U14630 (N_14630,N_14447,N_14264);
nor U14631 (N_14631,N_14282,N_14338);
nand U14632 (N_14632,N_14361,N_14445);
nand U14633 (N_14633,N_14280,N_14463);
or U14634 (N_14634,N_14478,N_14374);
or U14635 (N_14635,N_14265,N_14319);
nand U14636 (N_14636,N_14291,N_14302);
or U14637 (N_14637,N_14327,N_14437);
or U14638 (N_14638,N_14354,N_14380);
or U14639 (N_14639,N_14400,N_14480);
nand U14640 (N_14640,N_14358,N_14263);
nor U14641 (N_14641,N_14337,N_14355);
or U14642 (N_14642,N_14350,N_14494);
nand U14643 (N_14643,N_14364,N_14386);
nor U14644 (N_14644,N_14314,N_14315);
nor U14645 (N_14645,N_14460,N_14320);
nand U14646 (N_14646,N_14367,N_14381);
nand U14647 (N_14647,N_14487,N_14437);
nor U14648 (N_14648,N_14316,N_14285);
and U14649 (N_14649,N_14321,N_14276);
nor U14650 (N_14650,N_14331,N_14272);
and U14651 (N_14651,N_14333,N_14338);
xnor U14652 (N_14652,N_14371,N_14342);
nand U14653 (N_14653,N_14323,N_14432);
and U14654 (N_14654,N_14343,N_14485);
nor U14655 (N_14655,N_14325,N_14285);
nor U14656 (N_14656,N_14447,N_14420);
nor U14657 (N_14657,N_14320,N_14444);
or U14658 (N_14658,N_14456,N_14369);
or U14659 (N_14659,N_14385,N_14319);
or U14660 (N_14660,N_14354,N_14370);
and U14661 (N_14661,N_14265,N_14424);
nor U14662 (N_14662,N_14446,N_14496);
and U14663 (N_14663,N_14251,N_14318);
nand U14664 (N_14664,N_14446,N_14396);
and U14665 (N_14665,N_14342,N_14376);
nand U14666 (N_14666,N_14480,N_14311);
and U14667 (N_14667,N_14285,N_14263);
or U14668 (N_14668,N_14289,N_14315);
and U14669 (N_14669,N_14272,N_14356);
and U14670 (N_14670,N_14302,N_14441);
nor U14671 (N_14671,N_14415,N_14259);
nor U14672 (N_14672,N_14435,N_14361);
nor U14673 (N_14673,N_14468,N_14382);
nor U14674 (N_14674,N_14411,N_14463);
nor U14675 (N_14675,N_14485,N_14450);
xnor U14676 (N_14676,N_14318,N_14470);
nor U14677 (N_14677,N_14468,N_14442);
or U14678 (N_14678,N_14385,N_14473);
nand U14679 (N_14679,N_14345,N_14442);
xnor U14680 (N_14680,N_14453,N_14496);
nand U14681 (N_14681,N_14418,N_14270);
or U14682 (N_14682,N_14384,N_14388);
and U14683 (N_14683,N_14417,N_14251);
or U14684 (N_14684,N_14311,N_14359);
nand U14685 (N_14685,N_14458,N_14322);
and U14686 (N_14686,N_14435,N_14401);
nor U14687 (N_14687,N_14383,N_14471);
nand U14688 (N_14688,N_14277,N_14463);
nand U14689 (N_14689,N_14320,N_14407);
xnor U14690 (N_14690,N_14348,N_14274);
nor U14691 (N_14691,N_14451,N_14259);
nor U14692 (N_14692,N_14254,N_14326);
and U14693 (N_14693,N_14434,N_14322);
or U14694 (N_14694,N_14362,N_14454);
nand U14695 (N_14695,N_14499,N_14397);
and U14696 (N_14696,N_14327,N_14412);
nand U14697 (N_14697,N_14274,N_14261);
nand U14698 (N_14698,N_14413,N_14385);
nand U14699 (N_14699,N_14450,N_14463);
nand U14700 (N_14700,N_14335,N_14343);
and U14701 (N_14701,N_14386,N_14351);
or U14702 (N_14702,N_14414,N_14251);
nor U14703 (N_14703,N_14356,N_14476);
and U14704 (N_14704,N_14438,N_14308);
or U14705 (N_14705,N_14255,N_14485);
nor U14706 (N_14706,N_14272,N_14391);
and U14707 (N_14707,N_14377,N_14437);
and U14708 (N_14708,N_14273,N_14370);
and U14709 (N_14709,N_14272,N_14477);
nor U14710 (N_14710,N_14250,N_14307);
nor U14711 (N_14711,N_14483,N_14318);
nand U14712 (N_14712,N_14454,N_14399);
nand U14713 (N_14713,N_14354,N_14495);
nand U14714 (N_14714,N_14369,N_14298);
and U14715 (N_14715,N_14349,N_14257);
and U14716 (N_14716,N_14330,N_14342);
xnor U14717 (N_14717,N_14435,N_14329);
nand U14718 (N_14718,N_14301,N_14303);
nand U14719 (N_14719,N_14250,N_14274);
and U14720 (N_14720,N_14346,N_14278);
and U14721 (N_14721,N_14378,N_14361);
nand U14722 (N_14722,N_14366,N_14295);
and U14723 (N_14723,N_14371,N_14490);
nand U14724 (N_14724,N_14439,N_14448);
nor U14725 (N_14725,N_14415,N_14420);
or U14726 (N_14726,N_14419,N_14286);
or U14727 (N_14727,N_14254,N_14327);
nor U14728 (N_14728,N_14286,N_14370);
or U14729 (N_14729,N_14423,N_14253);
or U14730 (N_14730,N_14407,N_14377);
or U14731 (N_14731,N_14464,N_14467);
or U14732 (N_14732,N_14349,N_14252);
and U14733 (N_14733,N_14488,N_14420);
xnor U14734 (N_14734,N_14481,N_14435);
nand U14735 (N_14735,N_14349,N_14465);
and U14736 (N_14736,N_14486,N_14354);
xor U14737 (N_14737,N_14342,N_14265);
or U14738 (N_14738,N_14318,N_14407);
nand U14739 (N_14739,N_14253,N_14415);
or U14740 (N_14740,N_14388,N_14344);
nor U14741 (N_14741,N_14490,N_14253);
or U14742 (N_14742,N_14440,N_14377);
and U14743 (N_14743,N_14296,N_14340);
xnor U14744 (N_14744,N_14426,N_14384);
or U14745 (N_14745,N_14481,N_14439);
or U14746 (N_14746,N_14483,N_14468);
nor U14747 (N_14747,N_14307,N_14297);
or U14748 (N_14748,N_14462,N_14299);
nor U14749 (N_14749,N_14435,N_14414);
nor U14750 (N_14750,N_14734,N_14671);
and U14751 (N_14751,N_14526,N_14708);
and U14752 (N_14752,N_14500,N_14563);
nand U14753 (N_14753,N_14518,N_14697);
nand U14754 (N_14754,N_14561,N_14644);
nor U14755 (N_14755,N_14608,N_14684);
or U14756 (N_14756,N_14728,N_14506);
xor U14757 (N_14757,N_14604,N_14724);
nor U14758 (N_14758,N_14742,N_14638);
nand U14759 (N_14759,N_14596,N_14619);
nor U14760 (N_14760,N_14560,N_14590);
and U14761 (N_14761,N_14562,N_14670);
nor U14762 (N_14762,N_14584,N_14542);
nor U14763 (N_14763,N_14587,N_14629);
or U14764 (N_14764,N_14693,N_14568);
xnor U14765 (N_14765,N_14632,N_14667);
xor U14766 (N_14766,N_14717,N_14741);
nand U14767 (N_14767,N_14598,N_14557);
and U14768 (N_14768,N_14586,N_14656);
xnor U14769 (N_14769,N_14660,N_14532);
nor U14770 (N_14770,N_14744,N_14599);
or U14771 (N_14771,N_14624,N_14680);
nor U14772 (N_14772,N_14544,N_14726);
nor U14773 (N_14773,N_14652,N_14605);
or U14774 (N_14774,N_14621,N_14623);
nand U14775 (N_14775,N_14564,N_14633);
xor U14776 (N_14776,N_14558,N_14649);
and U14777 (N_14777,N_14601,N_14729);
nand U14778 (N_14778,N_14669,N_14740);
nand U14779 (N_14779,N_14748,N_14688);
and U14780 (N_14780,N_14749,N_14646);
nand U14781 (N_14781,N_14522,N_14574);
and U14782 (N_14782,N_14559,N_14578);
nor U14783 (N_14783,N_14692,N_14501);
and U14784 (N_14784,N_14714,N_14556);
nand U14785 (N_14785,N_14746,N_14735);
and U14786 (N_14786,N_14650,N_14612);
nand U14787 (N_14787,N_14687,N_14583);
nand U14788 (N_14788,N_14585,N_14682);
and U14789 (N_14789,N_14627,N_14747);
and U14790 (N_14790,N_14706,N_14527);
nand U14791 (N_14791,N_14739,N_14538);
nand U14792 (N_14792,N_14659,N_14529);
nor U14793 (N_14793,N_14620,N_14700);
and U14794 (N_14794,N_14647,N_14720);
nor U14795 (N_14795,N_14551,N_14615);
xor U14796 (N_14796,N_14645,N_14676);
nand U14797 (N_14797,N_14613,N_14512);
or U14798 (N_14798,N_14639,N_14503);
and U14799 (N_14799,N_14625,N_14514);
nand U14800 (N_14800,N_14548,N_14600);
nor U14801 (N_14801,N_14655,N_14549);
or U14802 (N_14802,N_14709,N_14721);
or U14803 (N_14803,N_14504,N_14642);
nor U14804 (N_14804,N_14530,N_14733);
and U14805 (N_14805,N_14634,N_14705);
or U14806 (N_14806,N_14525,N_14715);
nor U14807 (N_14807,N_14694,N_14609);
nand U14808 (N_14808,N_14580,N_14658);
nand U14809 (N_14809,N_14537,N_14555);
nor U14810 (N_14810,N_14702,N_14622);
nor U14811 (N_14811,N_14505,N_14543);
or U14812 (N_14812,N_14677,N_14571);
and U14813 (N_14813,N_14573,N_14631);
nand U14814 (N_14814,N_14743,N_14554);
or U14815 (N_14815,N_14626,N_14699);
nor U14816 (N_14816,N_14704,N_14679);
or U14817 (N_14817,N_14616,N_14651);
and U14818 (N_14818,N_14535,N_14657);
or U14819 (N_14819,N_14592,N_14534);
or U14820 (N_14820,N_14614,N_14618);
or U14821 (N_14821,N_14691,N_14567);
and U14822 (N_14822,N_14701,N_14540);
and U14823 (N_14823,N_14575,N_14536);
nor U14824 (N_14824,N_14695,N_14738);
and U14825 (N_14825,N_14606,N_14509);
or U14826 (N_14826,N_14519,N_14730);
xor U14827 (N_14827,N_14594,N_14665);
and U14828 (N_14828,N_14610,N_14516);
nand U14829 (N_14829,N_14666,N_14593);
nand U14830 (N_14830,N_14648,N_14528);
or U14831 (N_14831,N_14675,N_14722);
and U14832 (N_14832,N_14588,N_14510);
or U14833 (N_14833,N_14703,N_14672);
xnor U14834 (N_14834,N_14524,N_14508);
and U14835 (N_14835,N_14547,N_14541);
nand U14836 (N_14836,N_14602,N_14582);
and U14837 (N_14837,N_14546,N_14686);
or U14838 (N_14838,N_14552,N_14520);
or U14839 (N_14839,N_14569,N_14607);
and U14840 (N_14840,N_14727,N_14674);
nor U14841 (N_14841,N_14502,N_14523);
or U14842 (N_14842,N_14635,N_14511);
nor U14843 (N_14843,N_14630,N_14597);
or U14844 (N_14844,N_14572,N_14566);
and U14845 (N_14845,N_14617,N_14673);
and U14846 (N_14846,N_14689,N_14661);
nor U14847 (N_14847,N_14531,N_14641);
nor U14848 (N_14848,N_14515,N_14736);
nand U14849 (N_14849,N_14513,N_14517);
nand U14850 (N_14850,N_14685,N_14698);
and U14851 (N_14851,N_14579,N_14710);
nand U14852 (N_14852,N_14595,N_14707);
and U14853 (N_14853,N_14718,N_14550);
and U14854 (N_14854,N_14696,N_14637);
nor U14855 (N_14855,N_14732,N_14663);
or U14856 (N_14856,N_14681,N_14712);
or U14857 (N_14857,N_14719,N_14636);
nand U14858 (N_14858,N_14654,N_14521);
nand U14859 (N_14859,N_14589,N_14662);
and U14860 (N_14860,N_14723,N_14737);
nor U14861 (N_14861,N_14711,N_14581);
or U14862 (N_14862,N_14678,N_14664);
nor U14863 (N_14863,N_14628,N_14731);
xor U14864 (N_14864,N_14591,N_14713);
nand U14865 (N_14865,N_14716,N_14545);
nor U14866 (N_14866,N_14668,N_14745);
and U14867 (N_14867,N_14576,N_14725);
nand U14868 (N_14868,N_14507,N_14643);
nor U14869 (N_14869,N_14653,N_14611);
or U14870 (N_14870,N_14553,N_14640);
and U14871 (N_14871,N_14565,N_14603);
and U14872 (N_14872,N_14533,N_14539);
nand U14873 (N_14873,N_14690,N_14683);
nor U14874 (N_14874,N_14570,N_14577);
or U14875 (N_14875,N_14505,N_14669);
nand U14876 (N_14876,N_14727,N_14581);
nor U14877 (N_14877,N_14544,N_14566);
nand U14878 (N_14878,N_14625,N_14748);
nand U14879 (N_14879,N_14719,N_14608);
and U14880 (N_14880,N_14592,N_14721);
and U14881 (N_14881,N_14523,N_14730);
nand U14882 (N_14882,N_14527,N_14646);
or U14883 (N_14883,N_14679,N_14692);
and U14884 (N_14884,N_14555,N_14642);
xor U14885 (N_14885,N_14690,N_14720);
and U14886 (N_14886,N_14636,N_14599);
or U14887 (N_14887,N_14544,N_14616);
and U14888 (N_14888,N_14739,N_14608);
nor U14889 (N_14889,N_14503,N_14647);
nand U14890 (N_14890,N_14616,N_14541);
or U14891 (N_14891,N_14667,N_14634);
nor U14892 (N_14892,N_14743,N_14541);
nor U14893 (N_14893,N_14555,N_14690);
or U14894 (N_14894,N_14604,N_14688);
and U14895 (N_14895,N_14635,N_14537);
nand U14896 (N_14896,N_14546,N_14617);
or U14897 (N_14897,N_14656,N_14507);
or U14898 (N_14898,N_14542,N_14587);
or U14899 (N_14899,N_14594,N_14708);
nand U14900 (N_14900,N_14712,N_14614);
nor U14901 (N_14901,N_14630,N_14556);
or U14902 (N_14902,N_14675,N_14648);
nor U14903 (N_14903,N_14654,N_14630);
nor U14904 (N_14904,N_14723,N_14720);
nand U14905 (N_14905,N_14563,N_14725);
and U14906 (N_14906,N_14694,N_14698);
nor U14907 (N_14907,N_14746,N_14748);
and U14908 (N_14908,N_14630,N_14650);
xnor U14909 (N_14909,N_14508,N_14519);
nor U14910 (N_14910,N_14635,N_14744);
or U14911 (N_14911,N_14640,N_14548);
nor U14912 (N_14912,N_14549,N_14544);
and U14913 (N_14913,N_14735,N_14700);
and U14914 (N_14914,N_14515,N_14665);
and U14915 (N_14915,N_14543,N_14552);
nor U14916 (N_14916,N_14626,N_14511);
nor U14917 (N_14917,N_14595,N_14747);
nand U14918 (N_14918,N_14703,N_14534);
or U14919 (N_14919,N_14625,N_14691);
and U14920 (N_14920,N_14712,N_14528);
or U14921 (N_14921,N_14654,N_14556);
or U14922 (N_14922,N_14602,N_14559);
nand U14923 (N_14923,N_14500,N_14583);
nor U14924 (N_14924,N_14541,N_14511);
nor U14925 (N_14925,N_14607,N_14585);
nor U14926 (N_14926,N_14661,N_14729);
nand U14927 (N_14927,N_14569,N_14662);
and U14928 (N_14928,N_14662,N_14538);
and U14929 (N_14929,N_14607,N_14581);
nand U14930 (N_14930,N_14682,N_14600);
or U14931 (N_14931,N_14545,N_14602);
nor U14932 (N_14932,N_14554,N_14535);
and U14933 (N_14933,N_14564,N_14603);
and U14934 (N_14934,N_14566,N_14665);
or U14935 (N_14935,N_14737,N_14680);
and U14936 (N_14936,N_14581,N_14694);
or U14937 (N_14937,N_14677,N_14537);
or U14938 (N_14938,N_14637,N_14518);
nor U14939 (N_14939,N_14694,N_14590);
and U14940 (N_14940,N_14651,N_14593);
nor U14941 (N_14941,N_14741,N_14577);
nand U14942 (N_14942,N_14560,N_14665);
or U14943 (N_14943,N_14589,N_14570);
nand U14944 (N_14944,N_14733,N_14636);
nand U14945 (N_14945,N_14722,N_14669);
and U14946 (N_14946,N_14652,N_14739);
or U14947 (N_14947,N_14566,N_14575);
and U14948 (N_14948,N_14585,N_14653);
or U14949 (N_14949,N_14661,N_14731);
nand U14950 (N_14950,N_14617,N_14694);
and U14951 (N_14951,N_14551,N_14715);
or U14952 (N_14952,N_14560,N_14742);
or U14953 (N_14953,N_14605,N_14673);
and U14954 (N_14954,N_14539,N_14670);
nor U14955 (N_14955,N_14514,N_14695);
xnor U14956 (N_14956,N_14682,N_14582);
and U14957 (N_14957,N_14702,N_14685);
nor U14958 (N_14958,N_14513,N_14597);
or U14959 (N_14959,N_14523,N_14608);
or U14960 (N_14960,N_14564,N_14674);
nand U14961 (N_14961,N_14569,N_14691);
or U14962 (N_14962,N_14646,N_14739);
nor U14963 (N_14963,N_14503,N_14582);
or U14964 (N_14964,N_14542,N_14632);
and U14965 (N_14965,N_14566,N_14730);
or U14966 (N_14966,N_14542,N_14596);
or U14967 (N_14967,N_14718,N_14667);
nor U14968 (N_14968,N_14672,N_14567);
nand U14969 (N_14969,N_14637,N_14529);
nand U14970 (N_14970,N_14554,N_14660);
nor U14971 (N_14971,N_14733,N_14702);
and U14972 (N_14972,N_14728,N_14714);
nor U14973 (N_14973,N_14649,N_14714);
or U14974 (N_14974,N_14583,N_14746);
nor U14975 (N_14975,N_14741,N_14638);
and U14976 (N_14976,N_14643,N_14502);
nor U14977 (N_14977,N_14661,N_14559);
nand U14978 (N_14978,N_14522,N_14616);
nor U14979 (N_14979,N_14727,N_14537);
xor U14980 (N_14980,N_14551,N_14691);
or U14981 (N_14981,N_14590,N_14504);
and U14982 (N_14982,N_14615,N_14605);
or U14983 (N_14983,N_14584,N_14711);
nor U14984 (N_14984,N_14634,N_14513);
nand U14985 (N_14985,N_14588,N_14595);
nand U14986 (N_14986,N_14608,N_14678);
or U14987 (N_14987,N_14655,N_14560);
nor U14988 (N_14988,N_14533,N_14623);
or U14989 (N_14989,N_14697,N_14654);
or U14990 (N_14990,N_14712,N_14566);
or U14991 (N_14991,N_14614,N_14518);
or U14992 (N_14992,N_14549,N_14573);
and U14993 (N_14993,N_14673,N_14545);
or U14994 (N_14994,N_14741,N_14526);
and U14995 (N_14995,N_14674,N_14570);
nand U14996 (N_14996,N_14576,N_14583);
nor U14997 (N_14997,N_14590,N_14627);
and U14998 (N_14998,N_14670,N_14512);
nor U14999 (N_14999,N_14670,N_14558);
nand UO_0 (O_0,N_14833,N_14992);
nand UO_1 (O_1,N_14932,N_14779);
nand UO_2 (O_2,N_14822,N_14775);
nor UO_3 (O_3,N_14978,N_14818);
nor UO_4 (O_4,N_14791,N_14814);
and UO_5 (O_5,N_14759,N_14908);
nand UO_6 (O_6,N_14883,N_14807);
nor UO_7 (O_7,N_14935,N_14837);
and UO_8 (O_8,N_14898,N_14783);
and UO_9 (O_9,N_14856,N_14888);
or UO_10 (O_10,N_14868,N_14772);
or UO_11 (O_11,N_14823,N_14918);
or UO_12 (O_12,N_14790,N_14816);
or UO_13 (O_13,N_14892,N_14850);
nor UO_14 (O_14,N_14847,N_14957);
and UO_15 (O_15,N_14991,N_14758);
and UO_16 (O_16,N_14786,N_14889);
nand UO_17 (O_17,N_14828,N_14789);
xnor UO_18 (O_18,N_14801,N_14994);
and UO_19 (O_19,N_14795,N_14980);
or UO_20 (O_20,N_14834,N_14809);
nor UO_21 (O_21,N_14871,N_14975);
and UO_22 (O_22,N_14984,N_14947);
nand UO_23 (O_23,N_14766,N_14841);
nor UO_24 (O_24,N_14948,N_14949);
nand UO_25 (O_25,N_14753,N_14771);
nand UO_26 (O_26,N_14869,N_14925);
xnor UO_27 (O_27,N_14934,N_14757);
nand UO_28 (O_28,N_14910,N_14928);
or UO_29 (O_29,N_14907,N_14803);
or UO_30 (O_30,N_14880,N_14817);
xnor UO_31 (O_31,N_14887,N_14879);
and UO_32 (O_32,N_14829,N_14776);
xor UO_33 (O_33,N_14787,N_14838);
and UO_34 (O_34,N_14813,N_14895);
nor UO_35 (O_35,N_14805,N_14845);
or UO_36 (O_36,N_14930,N_14924);
and UO_37 (O_37,N_14941,N_14913);
nand UO_38 (O_38,N_14794,N_14964);
and UO_39 (O_39,N_14950,N_14893);
nor UO_40 (O_40,N_14974,N_14884);
and UO_41 (O_41,N_14863,N_14959);
nor UO_42 (O_42,N_14826,N_14970);
nor UO_43 (O_43,N_14840,N_14951);
and UO_44 (O_44,N_14848,N_14998);
nand UO_45 (O_45,N_14926,N_14755);
nor UO_46 (O_46,N_14800,N_14990);
nand UO_47 (O_47,N_14812,N_14846);
or UO_48 (O_48,N_14859,N_14979);
and UO_49 (O_49,N_14903,N_14937);
and UO_50 (O_50,N_14989,N_14915);
or UO_51 (O_51,N_14919,N_14986);
or UO_52 (O_52,N_14923,N_14890);
nor UO_53 (O_53,N_14760,N_14894);
nand UO_54 (O_54,N_14774,N_14799);
xor UO_55 (O_55,N_14967,N_14770);
nor UO_56 (O_56,N_14917,N_14969);
and UO_57 (O_57,N_14927,N_14851);
nor UO_58 (O_58,N_14897,N_14977);
or UO_59 (O_59,N_14988,N_14874);
or UO_60 (O_60,N_14839,N_14798);
nand UO_61 (O_61,N_14756,N_14855);
nor UO_62 (O_62,N_14982,N_14768);
nor UO_63 (O_63,N_14909,N_14778);
and UO_64 (O_64,N_14983,N_14796);
nor UO_65 (O_65,N_14832,N_14797);
nor UO_66 (O_66,N_14875,N_14881);
nor UO_67 (O_67,N_14912,N_14905);
xor UO_68 (O_68,N_14804,N_14751);
or UO_69 (O_69,N_14882,N_14831);
xor UO_70 (O_70,N_14938,N_14965);
nor UO_71 (O_71,N_14858,N_14953);
nor UO_72 (O_72,N_14830,N_14784);
and UO_73 (O_73,N_14782,N_14933);
nand UO_74 (O_74,N_14860,N_14844);
or UO_75 (O_75,N_14997,N_14878);
or UO_76 (O_76,N_14849,N_14958);
and UO_77 (O_77,N_14940,N_14802);
or UO_78 (O_78,N_14781,N_14946);
nor UO_79 (O_79,N_14857,N_14763);
nor UO_80 (O_80,N_14921,N_14955);
and UO_81 (O_81,N_14891,N_14825);
or UO_82 (O_82,N_14854,N_14793);
nand UO_83 (O_83,N_14780,N_14864);
nand UO_84 (O_84,N_14999,N_14899);
or UO_85 (O_85,N_14827,N_14931);
nand UO_86 (O_86,N_14963,N_14916);
and UO_87 (O_87,N_14769,N_14767);
nor UO_88 (O_88,N_14993,N_14996);
xor UO_89 (O_89,N_14981,N_14808);
nor UO_90 (O_90,N_14810,N_14985);
and UO_91 (O_91,N_14815,N_14976);
and UO_92 (O_92,N_14853,N_14942);
nor UO_93 (O_93,N_14852,N_14902);
nand UO_94 (O_94,N_14872,N_14995);
nand UO_95 (O_95,N_14956,N_14762);
xnor UO_96 (O_96,N_14945,N_14962);
or UO_97 (O_97,N_14811,N_14877);
nor UO_98 (O_98,N_14911,N_14939);
and UO_99 (O_99,N_14904,N_14922);
or UO_100 (O_100,N_14842,N_14765);
and UO_101 (O_101,N_14806,N_14824);
or UO_102 (O_102,N_14867,N_14886);
nand UO_103 (O_103,N_14987,N_14764);
nor UO_104 (O_104,N_14966,N_14792);
and UO_105 (O_105,N_14865,N_14752);
or UO_106 (O_106,N_14972,N_14896);
or UO_107 (O_107,N_14885,N_14866);
nand UO_108 (O_108,N_14873,N_14968);
and UO_109 (O_109,N_14876,N_14773);
or UO_110 (O_110,N_14901,N_14971);
or UO_111 (O_111,N_14761,N_14943);
nand UO_112 (O_112,N_14936,N_14920);
nor UO_113 (O_113,N_14861,N_14750);
nor UO_114 (O_114,N_14836,N_14835);
or UO_115 (O_115,N_14821,N_14944);
nor UO_116 (O_116,N_14914,N_14960);
or UO_117 (O_117,N_14862,N_14929);
nand UO_118 (O_118,N_14785,N_14973);
or UO_119 (O_119,N_14961,N_14906);
nor UO_120 (O_120,N_14820,N_14952);
nand UO_121 (O_121,N_14954,N_14788);
and UO_122 (O_122,N_14843,N_14777);
or UO_123 (O_123,N_14819,N_14754);
and UO_124 (O_124,N_14900,N_14870);
or UO_125 (O_125,N_14903,N_14897);
nor UO_126 (O_126,N_14846,N_14766);
nor UO_127 (O_127,N_14927,N_14880);
nor UO_128 (O_128,N_14824,N_14771);
or UO_129 (O_129,N_14984,N_14750);
or UO_130 (O_130,N_14788,N_14762);
nor UO_131 (O_131,N_14986,N_14929);
and UO_132 (O_132,N_14769,N_14908);
or UO_133 (O_133,N_14787,N_14764);
nand UO_134 (O_134,N_14835,N_14843);
and UO_135 (O_135,N_14893,N_14835);
nor UO_136 (O_136,N_14978,N_14855);
nand UO_137 (O_137,N_14971,N_14864);
nor UO_138 (O_138,N_14972,N_14763);
and UO_139 (O_139,N_14829,N_14831);
or UO_140 (O_140,N_14794,N_14995);
nand UO_141 (O_141,N_14815,N_14963);
or UO_142 (O_142,N_14893,N_14825);
and UO_143 (O_143,N_14804,N_14988);
nor UO_144 (O_144,N_14951,N_14822);
or UO_145 (O_145,N_14880,N_14900);
nor UO_146 (O_146,N_14880,N_14954);
and UO_147 (O_147,N_14855,N_14794);
nand UO_148 (O_148,N_14971,N_14834);
nand UO_149 (O_149,N_14792,N_14917);
and UO_150 (O_150,N_14906,N_14992);
or UO_151 (O_151,N_14833,N_14751);
and UO_152 (O_152,N_14786,N_14982);
and UO_153 (O_153,N_14998,N_14949);
or UO_154 (O_154,N_14856,N_14759);
nand UO_155 (O_155,N_14953,N_14827);
and UO_156 (O_156,N_14864,N_14954);
xor UO_157 (O_157,N_14953,N_14955);
nor UO_158 (O_158,N_14944,N_14800);
nor UO_159 (O_159,N_14860,N_14957);
or UO_160 (O_160,N_14878,N_14819);
or UO_161 (O_161,N_14850,N_14960);
and UO_162 (O_162,N_14967,N_14949);
nor UO_163 (O_163,N_14796,N_14814);
nor UO_164 (O_164,N_14985,N_14852);
or UO_165 (O_165,N_14792,N_14892);
nor UO_166 (O_166,N_14777,N_14944);
or UO_167 (O_167,N_14838,N_14960);
nor UO_168 (O_168,N_14993,N_14846);
or UO_169 (O_169,N_14815,N_14839);
and UO_170 (O_170,N_14871,N_14948);
and UO_171 (O_171,N_14867,N_14823);
nand UO_172 (O_172,N_14853,N_14751);
and UO_173 (O_173,N_14925,N_14899);
and UO_174 (O_174,N_14912,N_14870);
nand UO_175 (O_175,N_14756,N_14842);
and UO_176 (O_176,N_14935,N_14905);
nand UO_177 (O_177,N_14936,N_14903);
nor UO_178 (O_178,N_14890,N_14848);
nand UO_179 (O_179,N_14813,N_14757);
and UO_180 (O_180,N_14772,N_14754);
xor UO_181 (O_181,N_14771,N_14879);
nor UO_182 (O_182,N_14866,N_14948);
nor UO_183 (O_183,N_14816,N_14821);
or UO_184 (O_184,N_14834,N_14827);
nor UO_185 (O_185,N_14948,N_14755);
or UO_186 (O_186,N_14782,N_14924);
nor UO_187 (O_187,N_14787,N_14836);
and UO_188 (O_188,N_14956,N_14981);
and UO_189 (O_189,N_14922,N_14933);
and UO_190 (O_190,N_14966,N_14952);
nand UO_191 (O_191,N_14994,N_14776);
nand UO_192 (O_192,N_14792,N_14772);
and UO_193 (O_193,N_14807,N_14837);
nor UO_194 (O_194,N_14844,N_14864);
and UO_195 (O_195,N_14957,N_14820);
nor UO_196 (O_196,N_14832,N_14835);
nand UO_197 (O_197,N_14866,N_14925);
and UO_198 (O_198,N_14787,N_14950);
and UO_199 (O_199,N_14851,N_14946);
or UO_200 (O_200,N_14818,N_14813);
and UO_201 (O_201,N_14949,N_14847);
nand UO_202 (O_202,N_14755,N_14847);
and UO_203 (O_203,N_14996,N_14961);
and UO_204 (O_204,N_14999,N_14958);
and UO_205 (O_205,N_14946,N_14827);
or UO_206 (O_206,N_14844,N_14812);
nand UO_207 (O_207,N_14974,N_14808);
nor UO_208 (O_208,N_14812,N_14854);
nor UO_209 (O_209,N_14853,N_14851);
or UO_210 (O_210,N_14796,N_14956);
and UO_211 (O_211,N_14825,N_14931);
nor UO_212 (O_212,N_14956,N_14991);
and UO_213 (O_213,N_14842,N_14931);
and UO_214 (O_214,N_14963,N_14932);
and UO_215 (O_215,N_14976,N_14858);
nor UO_216 (O_216,N_14876,N_14850);
or UO_217 (O_217,N_14871,N_14992);
and UO_218 (O_218,N_14867,N_14759);
nand UO_219 (O_219,N_14858,N_14997);
nand UO_220 (O_220,N_14985,N_14812);
xor UO_221 (O_221,N_14938,N_14970);
or UO_222 (O_222,N_14769,N_14993);
or UO_223 (O_223,N_14962,N_14840);
or UO_224 (O_224,N_14914,N_14966);
nor UO_225 (O_225,N_14762,N_14780);
or UO_226 (O_226,N_14883,N_14803);
nor UO_227 (O_227,N_14944,N_14988);
nand UO_228 (O_228,N_14894,N_14925);
and UO_229 (O_229,N_14825,N_14913);
and UO_230 (O_230,N_14925,N_14753);
or UO_231 (O_231,N_14959,N_14987);
nor UO_232 (O_232,N_14820,N_14939);
nand UO_233 (O_233,N_14956,N_14939);
xnor UO_234 (O_234,N_14789,N_14970);
or UO_235 (O_235,N_14845,N_14853);
or UO_236 (O_236,N_14871,N_14807);
and UO_237 (O_237,N_14974,N_14940);
nand UO_238 (O_238,N_14992,N_14774);
or UO_239 (O_239,N_14993,N_14887);
nor UO_240 (O_240,N_14887,N_14964);
nor UO_241 (O_241,N_14882,N_14950);
nand UO_242 (O_242,N_14963,N_14957);
nor UO_243 (O_243,N_14917,N_14933);
or UO_244 (O_244,N_14750,N_14858);
or UO_245 (O_245,N_14906,N_14935);
or UO_246 (O_246,N_14806,N_14847);
nor UO_247 (O_247,N_14977,N_14984);
nand UO_248 (O_248,N_14928,N_14803);
and UO_249 (O_249,N_14828,N_14928);
nand UO_250 (O_250,N_14753,N_14848);
nor UO_251 (O_251,N_14891,N_14773);
or UO_252 (O_252,N_14992,N_14937);
nor UO_253 (O_253,N_14922,N_14808);
nor UO_254 (O_254,N_14880,N_14803);
and UO_255 (O_255,N_14754,N_14937);
nand UO_256 (O_256,N_14942,N_14817);
nor UO_257 (O_257,N_14958,N_14910);
nor UO_258 (O_258,N_14919,N_14763);
and UO_259 (O_259,N_14903,N_14967);
and UO_260 (O_260,N_14960,N_14851);
nor UO_261 (O_261,N_14893,N_14760);
or UO_262 (O_262,N_14996,N_14767);
nand UO_263 (O_263,N_14844,N_14794);
nor UO_264 (O_264,N_14968,N_14825);
nor UO_265 (O_265,N_14847,N_14807);
or UO_266 (O_266,N_14993,N_14915);
and UO_267 (O_267,N_14870,N_14839);
nand UO_268 (O_268,N_14760,N_14904);
or UO_269 (O_269,N_14774,N_14932);
nor UO_270 (O_270,N_14996,N_14926);
and UO_271 (O_271,N_14763,N_14809);
nor UO_272 (O_272,N_14897,N_14924);
nand UO_273 (O_273,N_14817,N_14990);
nand UO_274 (O_274,N_14873,N_14887);
nor UO_275 (O_275,N_14788,N_14945);
nand UO_276 (O_276,N_14816,N_14964);
and UO_277 (O_277,N_14766,N_14774);
nand UO_278 (O_278,N_14891,N_14923);
nor UO_279 (O_279,N_14792,N_14884);
nor UO_280 (O_280,N_14902,N_14829);
nor UO_281 (O_281,N_14989,N_14953);
and UO_282 (O_282,N_14866,N_14804);
and UO_283 (O_283,N_14883,N_14754);
nand UO_284 (O_284,N_14972,N_14975);
nor UO_285 (O_285,N_14799,N_14893);
and UO_286 (O_286,N_14928,N_14765);
and UO_287 (O_287,N_14853,N_14912);
nand UO_288 (O_288,N_14879,N_14975);
nand UO_289 (O_289,N_14964,N_14780);
nor UO_290 (O_290,N_14767,N_14793);
and UO_291 (O_291,N_14850,N_14824);
nor UO_292 (O_292,N_14838,N_14922);
and UO_293 (O_293,N_14855,N_14903);
or UO_294 (O_294,N_14870,N_14961);
nor UO_295 (O_295,N_14805,N_14781);
nand UO_296 (O_296,N_14799,N_14787);
nand UO_297 (O_297,N_14946,N_14910);
or UO_298 (O_298,N_14751,N_14876);
nor UO_299 (O_299,N_14815,N_14933);
nor UO_300 (O_300,N_14780,N_14859);
or UO_301 (O_301,N_14944,N_14897);
and UO_302 (O_302,N_14788,N_14867);
nand UO_303 (O_303,N_14930,N_14872);
nor UO_304 (O_304,N_14869,N_14913);
nand UO_305 (O_305,N_14895,N_14927);
nor UO_306 (O_306,N_14803,N_14821);
nor UO_307 (O_307,N_14877,N_14787);
or UO_308 (O_308,N_14846,N_14982);
nor UO_309 (O_309,N_14780,N_14961);
and UO_310 (O_310,N_14757,N_14872);
xnor UO_311 (O_311,N_14876,N_14862);
or UO_312 (O_312,N_14799,N_14818);
or UO_313 (O_313,N_14836,N_14935);
and UO_314 (O_314,N_14926,N_14903);
or UO_315 (O_315,N_14927,N_14873);
nor UO_316 (O_316,N_14922,N_14947);
and UO_317 (O_317,N_14927,N_14818);
nor UO_318 (O_318,N_14965,N_14913);
and UO_319 (O_319,N_14781,N_14758);
or UO_320 (O_320,N_14827,N_14904);
or UO_321 (O_321,N_14942,N_14949);
nor UO_322 (O_322,N_14958,N_14898);
and UO_323 (O_323,N_14843,N_14897);
or UO_324 (O_324,N_14801,N_14883);
nand UO_325 (O_325,N_14960,N_14936);
nand UO_326 (O_326,N_14761,N_14797);
nand UO_327 (O_327,N_14752,N_14970);
or UO_328 (O_328,N_14971,N_14982);
xnor UO_329 (O_329,N_14805,N_14875);
nand UO_330 (O_330,N_14787,N_14922);
nor UO_331 (O_331,N_14985,N_14944);
nor UO_332 (O_332,N_14781,N_14912);
nand UO_333 (O_333,N_14757,N_14863);
and UO_334 (O_334,N_14907,N_14793);
nand UO_335 (O_335,N_14781,N_14925);
nand UO_336 (O_336,N_14801,N_14858);
and UO_337 (O_337,N_14977,N_14969);
and UO_338 (O_338,N_14892,N_14912);
or UO_339 (O_339,N_14987,N_14765);
nand UO_340 (O_340,N_14896,N_14978);
nand UO_341 (O_341,N_14757,N_14969);
nand UO_342 (O_342,N_14878,N_14817);
nand UO_343 (O_343,N_14950,N_14785);
nand UO_344 (O_344,N_14882,N_14761);
nand UO_345 (O_345,N_14900,N_14871);
nand UO_346 (O_346,N_14816,N_14928);
nand UO_347 (O_347,N_14914,N_14781);
and UO_348 (O_348,N_14886,N_14970);
or UO_349 (O_349,N_14801,N_14972);
nor UO_350 (O_350,N_14756,N_14908);
nand UO_351 (O_351,N_14911,N_14802);
or UO_352 (O_352,N_14895,N_14751);
and UO_353 (O_353,N_14854,N_14786);
xnor UO_354 (O_354,N_14854,N_14794);
nand UO_355 (O_355,N_14758,N_14895);
and UO_356 (O_356,N_14863,N_14880);
nor UO_357 (O_357,N_14996,N_14974);
and UO_358 (O_358,N_14821,N_14938);
nor UO_359 (O_359,N_14845,N_14771);
or UO_360 (O_360,N_14848,N_14846);
and UO_361 (O_361,N_14777,N_14937);
or UO_362 (O_362,N_14969,N_14781);
nor UO_363 (O_363,N_14898,N_14875);
nor UO_364 (O_364,N_14756,N_14971);
or UO_365 (O_365,N_14852,N_14901);
and UO_366 (O_366,N_14755,N_14994);
nor UO_367 (O_367,N_14953,N_14811);
nor UO_368 (O_368,N_14891,N_14851);
nor UO_369 (O_369,N_14968,N_14979);
nand UO_370 (O_370,N_14891,N_14879);
xor UO_371 (O_371,N_14782,N_14953);
xnor UO_372 (O_372,N_14907,N_14797);
and UO_373 (O_373,N_14850,N_14831);
nor UO_374 (O_374,N_14753,N_14755);
or UO_375 (O_375,N_14958,N_14924);
nor UO_376 (O_376,N_14781,N_14842);
nor UO_377 (O_377,N_14885,N_14998);
and UO_378 (O_378,N_14817,N_14835);
and UO_379 (O_379,N_14793,N_14756);
or UO_380 (O_380,N_14990,N_14985);
nor UO_381 (O_381,N_14856,N_14838);
or UO_382 (O_382,N_14750,N_14950);
or UO_383 (O_383,N_14867,N_14766);
nand UO_384 (O_384,N_14863,N_14905);
nand UO_385 (O_385,N_14925,N_14791);
and UO_386 (O_386,N_14835,N_14756);
nand UO_387 (O_387,N_14834,N_14842);
nand UO_388 (O_388,N_14757,N_14902);
nor UO_389 (O_389,N_14975,N_14865);
xnor UO_390 (O_390,N_14830,N_14839);
xor UO_391 (O_391,N_14977,N_14998);
or UO_392 (O_392,N_14787,N_14923);
nand UO_393 (O_393,N_14972,N_14750);
nand UO_394 (O_394,N_14793,N_14957);
and UO_395 (O_395,N_14882,N_14864);
nor UO_396 (O_396,N_14847,N_14771);
nand UO_397 (O_397,N_14771,N_14866);
or UO_398 (O_398,N_14783,N_14854);
and UO_399 (O_399,N_14991,N_14782);
or UO_400 (O_400,N_14980,N_14774);
nand UO_401 (O_401,N_14935,N_14826);
and UO_402 (O_402,N_14997,N_14891);
nor UO_403 (O_403,N_14963,N_14765);
nand UO_404 (O_404,N_14894,N_14885);
nand UO_405 (O_405,N_14833,N_14820);
nor UO_406 (O_406,N_14978,N_14790);
or UO_407 (O_407,N_14997,N_14841);
nor UO_408 (O_408,N_14782,N_14766);
and UO_409 (O_409,N_14980,N_14886);
nand UO_410 (O_410,N_14981,N_14941);
nand UO_411 (O_411,N_14886,N_14947);
nand UO_412 (O_412,N_14939,N_14800);
or UO_413 (O_413,N_14867,N_14780);
or UO_414 (O_414,N_14751,N_14808);
nor UO_415 (O_415,N_14837,N_14842);
nand UO_416 (O_416,N_14964,N_14754);
nor UO_417 (O_417,N_14845,N_14980);
nand UO_418 (O_418,N_14882,N_14796);
nand UO_419 (O_419,N_14963,N_14991);
or UO_420 (O_420,N_14878,N_14833);
or UO_421 (O_421,N_14901,N_14799);
or UO_422 (O_422,N_14911,N_14952);
nor UO_423 (O_423,N_14934,N_14964);
nor UO_424 (O_424,N_14813,N_14833);
nor UO_425 (O_425,N_14862,N_14908);
or UO_426 (O_426,N_14994,N_14880);
nor UO_427 (O_427,N_14995,N_14856);
or UO_428 (O_428,N_14995,N_14775);
nor UO_429 (O_429,N_14844,N_14865);
and UO_430 (O_430,N_14886,N_14819);
nor UO_431 (O_431,N_14804,N_14815);
and UO_432 (O_432,N_14998,N_14854);
and UO_433 (O_433,N_14846,N_14819);
and UO_434 (O_434,N_14794,N_14982);
and UO_435 (O_435,N_14983,N_14816);
nor UO_436 (O_436,N_14891,N_14850);
and UO_437 (O_437,N_14842,N_14987);
nand UO_438 (O_438,N_14913,N_14873);
nor UO_439 (O_439,N_14926,N_14797);
nor UO_440 (O_440,N_14864,N_14876);
nor UO_441 (O_441,N_14791,N_14890);
nand UO_442 (O_442,N_14971,N_14886);
nor UO_443 (O_443,N_14803,N_14834);
nor UO_444 (O_444,N_14799,N_14878);
or UO_445 (O_445,N_14828,N_14872);
nor UO_446 (O_446,N_14854,N_14763);
nor UO_447 (O_447,N_14792,N_14863);
nor UO_448 (O_448,N_14880,N_14794);
nor UO_449 (O_449,N_14765,N_14767);
or UO_450 (O_450,N_14915,N_14983);
and UO_451 (O_451,N_14783,N_14979);
or UO_452 (O_452,N_14923,N_14804);
and UO_453 (O_453,N_14899,N_14885);
or UO_454 (O_454,N_14982,N_14926);
nor UO_455 (O_455,N_14764,N_14847);
or UO_456 (O_456,N_14896,N_14994);
or UO_457 (O_457,N_14839,N_14818);
and UO_458 (O_458,N_14920,N_14774);
and UO_459 (O_459,N_14889,N_14840);
and UO_460 (O_460,N_14911,N_14975);
and UO_461 (O_461,N_14855,N_14974);
or UO_462 (O_462,N_14901,N_14882);
and UO_463 (O_463,N_14758,N_14948);
nor UO_464 (O_464,N_14866,N_14862);
nor UO_465 (O_465,N_14970,N_14950);
and UO_466 (O_466,N_14840,N_14996);
and UO_467 (O_467,N_14944,N_14942);
nand UO_468 (O_468,N_14890,N_14862);
or UO_469 (O_469,N_14990,N_14834);
or UO_470 (O_470,N_14862,N_14863);
and UO_471 (O_471,N_14880,N_14858);
and UO_472 (O_472,N_14926,N_14833);
and UO_473 (O_473,N_14903,N_14992);
nor UO_474 (O_474,N_14803,N_14978);
nand UO_475 (O_475,N_14788,N_14787);
nand UO_476 (O_476,N_14781,N_14798);
or UO_477 (O_477,N_14965,N_14910);
nor UO_478 (O_478,N_14875,N_14938);
and UO_479 (O_479,N_14948,N_14849);
nor UO_480 (O_480,N_14891,N_14810);
or UO_481 (O_481,N_14919,N_14825);
and UO_482 (O_482,N_14891,N_14847);
nor UO_483 (O_483,N_14943,N_14963);
or UO_484 (O_484,N_14900,N_14917);
or UO_485 (O_485,N_14968,N_14871);
nand UO_486 (O_486,N_14817,N_14944);
nor UO_487 (O_487,N_14797,N_14884);
and UO_488 (O_488,N_14811,N_14758);
and UO_489 (O_489,N_14769,N_14913);
and UO_490 (O_490,N_14966,N_14892);
or UO_491 (O_491,N_14830,N_14938);
or UO_492 (O_492,N_14868,N_14975);
or UO_493 (O_493,N_14805,N_14918);
or UO_494 (O_494,N_14792,N_14988);
nor UO_495 (O_495,N_14982,N_14812);
or UO_496 (O_496,N_14884,N_14782);
nand UO_497 (O_497,N_14995,N_14958);
or UO_498 (O_498,N_14986,N_14821);
or UO_499 (O_499,N_14855,N_14952);
or UO_500 (O_500,N_14812,N_14769);
or UO_501 (O_501,N_14860,N_14907);
nor UO_502 (O_502,N_14804,N_14856);
nor UO_503 (O_503,N_14977,N_14854);
nor UO_504 (O_504,N_14887,N_14903);
nor UO_505 (O_505,N_14758,N_14846);
nand UO_506 (O_506,N_14750,N_14988);
or UO_507 (O_507,N_14804,N_14753);
nor UO_508 (O_508,N_14842,N_14943);
nand UO_509 (O_509,N_14793,N_14875);
or UO_510 (O_510,N_14803,N_14762);
nor UO_511 (O_511,N_14867,N_14909);
and UO_512 (O_512,N_14841,N_14968);
nand UO_513 (O_513,N_14960,N_14926);
or UO_514 (O_514,N_14813,N_14875);
nor UO_515 (O_515,N_14849,N_14919);
nand UO_516 (O_516,N_14787,N_14837);
and UO_517 (O_517,N_14934,N_14931);
and UO_518 (O_518,N_14837,N_14978);
and UO_519 (O_519,N_14767,N_14772);
nor UO_520 (O_520,N_14878,N_14894);
nor UO_521 (O_521,N_14941,N_14862);
and UO_522 (O_522,N_14763,N_14979);
xnor UO_523 (O_523,N_14981,N_14974);
nor UO_524 (O_524,N_14750,N_14884);
and UO_525 (O_525,N_14756,N_14786);
and UO_526 (O_526,N_14989,N_14812);
or UO_527 (O_527,N_14786,N_14774);
or UO_528 (O_528,N_14824,N_14924);
nor UO_529 (O_529,N_14885,N_14974);
or UO_530 (O_530,N_14997,N_14835);
nand UO_531 (O_531,N_14945,N_14769);
nor UO_532 (O_532,N_14929,N_14821);
or UO_533 (O_533,N_14931,N_14998);
and UO_534 (O_534,N_14863,N_14878);
nor UO_535 (O_535,N_14814,N_14790);
or UO_536 (O_536,N_14909,N_14891);
nor UO_537 (O_537,N_14985,N_14800);
or UO_538 (O_538,N_14983,N_14921);
or UO_539 (O_539,N_14988,N_14998);
nand UO_540 (O_540,N_14815,N_14835);
or UO_541 (O_541,N_14811,N_14837);
xor UO_542 (O_542,N_14793,N_14963);
or UO_543 (O_543,N_14915,N_14848);
nor UO_544 (O_544,N_14846,N_14820);
nor UO_545 (O_545,N_14950,N_14887);
or UO_546 (O_546,N_14909,N_14954);
nor UO_547 (O_547,N_14770,N_14962);
or UO_548 (O_548,N_14875,N_14965);
and UO_549 (O_549,N_14963,N_14872);
nand UO_550 (O_550,N_14965,N_14884);
nor UO_551 (O_551,N_14884,N_14843);
nor UO_552 (O_552,N_14894,N_14889);
nand UO_553 (O_553,N_14806,N_14957);
and UO_554 (O_554,N_14785,N_14764);
and UO_555 (O_555,N_14854,N_14878);
nor UO_556 (O_556,N_14818,N_14982);
or UO_557 (O_557,N_14797,N_14854);
and UO_558 (O_558,N_14860,N_14762);
or UO_559 (O_559,N_14924,N_14816);
or UO_560 (O_560,N_14902,N_14842);
nand UO_561 (O_561,N_14927,N_14876);
nor UO_562 (O_562,N_14796,N_14947);
and UO_563 (O_563,N_14784,N_14787);
nor UO_564 (O_564,N_14901,N_14847);
nor UO_565 (O_565,N_14822,N_14886);
nor UO_566 (O_566,N_14917,N_14953);
xnor UO_567 (O_567,N_14863,N_14773);
nor UO_568 (O_568,N_14752,N_14912);
nor UO_569 (O_569,N_14785,N_14928);
or UO_570 (O_570,N_14803,N_14763);
or UO_571 (O_571,N_14793,N_14900);
or UO_572 (O_572,N_14853,N_14971);
nand UO_573 (O_573,N_14786,N_14870);
nand UO_574 (O_574,N_14793,N_14753);
nor UO_575 (O_575,N_14869,N_14864);
and UO_576 (O_576,N_14961,N_14840);
xnor UO_577 (O_577,N_14911,N_14843);
nand UO_578 (O_578,N_14916,N_14818);
nand UO_579 (O_579,N_14755,N_14776);
or UO_580 (O_580,N_14903,N_14800);
nor UO_581 (O_581,N_14948,N_14976);
nor UO_582 (O_582,N_14971,N_14989);
or UO_583 (O_583,N_14800,N_14816);
nor UO_584 (O_584,N_14862,N_14966);
and UO_585 (O_585,N_14968,N_14959);
or UO_586 (O_586,N_14932,N_14902);
nor UO_587 (O_587,N_14785,N_14822);
nand UO_588 (O_588,N_14812,N_14906);
nand UO_589 (O_589,N_14906,N_14969);
nand UO_590 (O_590,N_14820,N_14861);
nor UO_591 (O_591,N_14817,N_14823);
and UO_592 (O_592,N_14900,N_14892);
and UO_593 (O_593,N_14762,N_14869);
or UO_594 (O_594,N_14986,N_14914);
nand UO_595 (O_595,N_14858,N_14787);
nand UO_596 (O_596,N_14756,N_14824);
or UO_597 (O_597,N_14904,N_14999);
nor UO_598 (O_598,N_14771,N_14763);
or UO_599 (O_599,N_14755,N_14900);
and UO_600 (O_600,N_14802,N_14818);
nor UO_601 (O_601,N_14910,N_14757);
or UO_602 (O_602,N_14930,N_14888);
nor UO_603 (O_603,N_14873,N_14782);
and UO_604 (O_604,N_14772,N_14877);
nor UO_605 (O_605,N_14805,N_14942);
or UO_606 (O_606,N_14780,N_14857);
nand UO_607 (O_607,N_14867,N_14932);
or UO_608 (O_608,N_14797,N_14887);
nor UO_609 (O_609,N_14823,N_14932);
and UO_610 (O_610,N_14955,N_14810);
and UO_611 (O_611,N_14897,N_14793);
and UO_612 (O_612,N_14936,N_14916);
and UO_613 (O_613,N_14803,N_14991);
and UO_614 (O_614,N_14931,N_14772);
nand UO_615 (O_615,N_14912,N_14774);
xor UO_616 (O_616,N_14769,N_14915);
nor UO_617 (O_617,N_14805,N_14752);
nor UO_618 (O_618,N_14892,N_14819);
or UO_619 (O_619,N_14824,N_14983);
nand UO_620 (O_620,N_14910,N_14954);
xnor UO_621 (O_621,N_14986,N_14993);
nand UO_622 (O_622,N_14999,N_14858);
nor UO_623 (O_623,N_14772,N_14838);
or UO_624 (O_624,N_14875,N_14949);
nand UO_625 (O_625,N_14953,N_14915);
or UO_626 (O_626,N_14909,N_14822);
and UO_627 (O_627,N_14769,N_14855);
nand UO_628 (O_628,N_14998,N_14843);
and UO_629 (O_629,N_14867,N_14910);
nand UO_630 (O_630,N_14913,N_14964);
nand UO_631 (O_631,N_14777,N_14958);
or UO_632 (O_632,N_14869,N_14779);
or UO_633 (O_633,N_14984,N_14926);
or UO_634 (O_634,N_14975,N_14957);
and UO_635 (O_635,N_14789,N_14975);
nand UO_636 (O_636,N_14996,N_14867);
and UO_637 (O_637,N_14808,N_14893);
and UO_638 (O_638,N_14752,N_14896);
nand UO_639 (O_639,N_14999,N_14829);
nand UO_640 (O_640,N_14758,N_14995);
xnor UO_641 (O_641,N_14994,N_14917);
nand UO_642 (O_642,N_14882,N_14887);
nor UO_643 (O_643,N_14840,N_14796);
and UO_644 (O_644,N_14874,N_14818);
or UO_645 (O_645,N_14796,N_14888);
or UO_646 (O_646,N_14913,N_14797);
and UO_647 (O_647,N_14754,N_14918);
nor UO_648 (O_648,N_14904,N_14774);
and UO_649 (O_649,N_14950,N_14978);
and UO_650 (O_650,N_14759,N_14824);
or UO_651 (O_651,N_14863,N_14758);
or UO_652 (O_652,N_14976,N_14898);
nor UO_653 (O_653,N_14814,N_14997);
or UO_654 (O_654,N_14864,N_14938);
and UO_655 (O_655,N_14947,N_14908);
or UO_656 (O_656,N_14961,N_14831);
nor UO_657 (O_657,N_14962,N_14810);
and UO_658 (O_658,N_14859,N_14990);
nand UO_659 (O_659,N_14772,N_14827);
nor UO_660 (O_660,N_14940,N_14928);
nand UO_661 (O_661,N_14880,N_14778);
or UO_662 (O_662,N_14846,N_14965);
xnor UO_663 (O_663,N_14953,N_14835);
or UO_664 (O_664,N_14805,N_14887);
nand UO_665 (O_665,N_14879,N_14816);
nor UO_666 (O_666,N_14983,N_14756);
nand UO_667 (O_667,N_14998,N_14984);
nand UO_668 (O_668,N_14936,N_14918);
and UO_669 (O_669,N_14967,N_14918);
nand UO_670 (O_670,N_14956,N_14880);
or UO_671 (O_671,N_14796,N_14987);
nor UO_672 (O_672,N_14761,N_14796);
and UO_673 (O_673,N_14829,N_14886);
and UO_674 (O_674,N_14817,N_14955);
nor UO_675 (O_675,N_14986,N_14830);
nand UO_676 (O_676,N_14901,N_14798);
nand UO_677 (O_677,N_14995,N_14792);
nor UO_678 (O_678,N_14946,N_14971);
nand UO_679 (O_679,N_14869,N_14803);
or UO_680 (O_680,N_14782,N_14998);
and UO_681 (O_681,N_14793,N_14818);
nor UO_682 (O_682,N_14822,N_14755);
nor UO_683 (O_683,N_14984,N_14851);
and UO_684 (O_684,N_14809,N_14980);
or UO_685 (O_685,N_14994,N_14846);
or UO_686 (O_686,N_14790,N_14886);
nor UO_687 (O_687,N_14869,N_14847);
xor UO_688 (O_688,N_14755,N_14999);
nor UO_689 (O_689,N_14864,N_14931);
nand UO_690 (O_690,N_14870,N_14824);
nand UO_691 (O_691,N_14943,N_14815);
and UO_692 (O_692,N_14834,N_14787);
or UO_693 (O_693,N_14901,N_14930);
and UO_694 (O_694,N_14843,N_14771);
or UO_695 (O_695,N_14846,N_14946);
xnor UO_696 (O_696,N_14971,N_14947);
or UO_697 (O_697,N_14966,N_14866);
nand UO_698 (O_698,N_14817,N_14951);
or UO_699 (O_699,N_14919,N_14920);
and UO_700 (O_700,N_14927,N_14804);
and UO_701 (O_701,N_14931,N_14858);
nor UO_702 (O_702,N_14995,N_14816);
or UO_703 (O_703,N_14972,N_14946);
nand UO_704 (O_704,N_14963,N_14988);
nor UO_705 (O_705,N_14933,N_14948);
nand UO_706 (O_706,N_14906,N_14960);
xnor UO_707 (O_707,N_14975,N_14942);
nand UO_708 (O_708,N_14774,N_14943);
or UO_709 (O_709,N_14989,N_14926);
nor UO_710 (O_710,N_14890,N_14756);
nand UO_711 (O_711,N_14982,N_14996);
nor UO_712 (O_712,N_14948,N_14970);
and UO_713 (O_713,N_14818,N_14771);
and UO_714 (O_714,N_14894,N_14970);
or UO_715 (O_715,N_14990,N_14991);
nand UO_716 (O_716,N_14844,N_14787);
or UO_717 (O_717,N_14887,N_14849);
and UO_718 (O_718,N_14899,N_14779);
nor UO_719 (O_719,N_14863,N_14829);
nand UO_720 (O_720,N_14901,N_14859);
and UO_721 (O_721,N_14908,N_14834);
and UO_722 (O_722,N_14902,N_14878);
or UO_723 (O_723,N_14946,N_14816);
xnor UO_724 (O_724,N_14987,N_14794);
or UO_725 (O_725,N_14958,N_14830);
and UO_726 (O_726,N_14856,N_14863);
xor UO_727 (O_727,N_14781,N_14935);
or UO_728 (O_728,N_14777,N_14923);
nor UO_729 (O_729,N_14826,N_14943);
nand UO_730 (O_730,N_14773,N_14813);
nor UO_731 (O_731,N_14853,N_14842);
or UO_732 (O_732,N_14833,N_14900);
and UO_733 (O_733,N_14941,N_14924);
or UO_734 (O_734,N_14956,N_14816);
and UO_735 (O_735,N_14906,N_14802);
or UO_736 (O_736,N_14981,N_14782);
and UO_737 (O_737,N_14848,N_14767);
and UO_738 (O_738,N_14786,N_14824);
and UO_739 (O_739,N_14859,N_14793);
and UO_740 (O_740,N_14804,N_14857);
or UO_741 (O_741,N_14944,N_14900);
and UO_742 (O_742,N_14903,N_14822);
and UO_743 (O_743,N_14755,N_14961);
nor UO_744 (O_744,N_14965,N_14818);
or UO_745 (O_745,N_14943,N_14972);
nor UO_746 (O_746,N_14936,N_14823);
nand UO_747 (O_747,N_14932,N_14832);
or UO_748 (O_748,N_14880,N_14922);
and UO_749 (O_749,N_14981,N_14896);
nand UO_750 (O_750,N_14755,N_14922);
or UO_751 (O_751,N_14999,N_14992);
or UO_752 (O_752,N_14849,N_14884);
or UO_753 (O_753,N_14935,N_14782);
and UO_754 (O_754,N_14948,N_14848);
and UO_755 (O_755,N_14927,N_14944);
nand UO_756 (O_756,N_14866,N_14897);
or UO_757 (O_757,N_14995,N_14825);
nor UO_758 (O_758,N_14782,N_14774);
or UO_759 (O_759,N_14893,N_14774);
nor UO_760 (O_760,N_14915,N_14998);
nor UO_761 (O_761,N_14751,N_14776);
nor UO_762 (O_762,N_14889,N_14773);
nor UO_763 (O_763,N_14984,N_14937);
nand UO_764 (O_764,N_14961,N_14967);
and UO_765 (O_765,N_14919,N_14832);
nor UO_766 (O_766,N_14822,N_14882);
nand UO_767 (O_767,N_14970,N_14766);
nand UO_768 (O_768,N_14883,N_14788);
and UO_769 (O_769,N_14824,N_14993);
or UO_770 (O_770,N_14800,N_14963);
and UO_771 (O_771,N_14826,N_14905);
nor UO_772 (O_772,N_14833,N_14770);
nand UO_773 (O_773,N_14767,N_14979);
nand UO_774 (O_774,N_14786,N_14991);
and UO_775 (O_775,N_14916,N_14803);
or UO_776 (O_776,N_14884,N_14833);
nand UO_777 (O_777,N_14797,N_14990);
nand UO_778 (O_778,N_14875,N_14916);
and UO_779 (O_779,N_14808,N_14886);
or UO_780 (O_780,N_14952,N_14909);
and UO_781 (O_781,N_14930,N_14866);
nor UO_782 (O_782,N_14809,N_14765);
and UO_783 (O_783,N_14879,N_14800);
and UO_784 (O_784,N_14887,N_14753);
and UO_785 (O_785,N_14905,N_14920);
or UO_786 (O_786,N_14768,N_14894);
nand UO_787 (O_787,N_14814,N_14865);
nor UO_788 (O_788,N_14912,N_14893);
nor UO_789 (O_789,N_14882,N_14934);
nand UO_790 (O_790,N_14776,N_14880);
nor UO_791 (O_791,N_14792,N_14826);
nand UO_792 (O_792,N_14761,N_14856);
and UO_793 (O_793,N_14854,N_14919);
nor UO_794 (O_794,N_14751,N_14809);
nor UO_795 (O_795,N_14967,N_14758);
nor UO_796 (O_796,N_14775,N_14917);
and UO_797 (O_797,N_14948,N_14932);
and UO_798 (O_798,N_14899,N_14855);
and UO_799 (O_799,N_14917,N_14811);
or UO_800 (O_800,N_14751,N_14995);
and UO_801 (O_801,N_14767,N_14898);
nor UO_802 (O_802,N_14767,N_14977);
nand UO_803 (O_803,N_14892,N_14929);
or UO_804 (O_804,N_14987,N_14761);
or UO_805 (O_805,N_14968,N_14885);
nand UO_806 (O_806,N_14762,N_14988);
nor UO_807 (O_807,N_14994,N_14784);
or UO_808 (O_808,N_14802,N_14786);
nor UO_809 (O_809,N_14982,N_14828);
nor UO_810 (O_810,N_14917,N_14833);
nand UO_811 (O_811,N_14769,N_14805);
xnor UO_812 (O_812,N_14763,N_14950);
nor UO_813 (O_813,N_14871,N_14837);
or UO_814 (O_814,N_14852,N_14750);
or UO_815 (O_815,N_14791,N_14855);
or UO_816 (O_816,N_14990,N_14804);
and UO_817 (O_817,N_14778,N_14987);
nand UO_818 (O_818,N_14966,N_14884);
nand UO_819 (O_819,N_14973,N_14919);
or UO_820 (O_820,N_14935,N_14878);
or UO_821 (O_821,N_14793,N_14878);
xnor UO_822 (O_822,N_14886,N_14998);
nand UO_823 (O_823,N_14879,N_14984);
or UO_824 (O_824,N_14893,N_14769);
or UO_825 (O_825,N_14958,N_14785);
and UO_826 (O_826,N_14907,N_14818);
or UO_827 (O_827,N_14881,N_14886);
and UO_828 (O_828,N_14850,N_14921);
nor UO_829 (O_829,N_14928,N_14880);
nor UO_830 (O_830,N_14750,N_14848);
and UO_831 (O_831,N_14876,N_14886);
or UO_832 (O_832,N_14841,N_14955);
nand UO_833 (O_833,N_14999,N_14929);
and UO_834 (O_834,N_14993,N_14779);
nor UO_835 (O_835,N_14755,N_14750);
nand UO_836 (O_836,N_14897,N_14882);
nor UO_837 (O_837,N_14789,N_14952);
nand UO_838 (O_838,N_14784,N_14826);
nand UO_839 (O_839,N_14965,N_14761);
nor UO_840 (O_840,N_14967,N_14801);
and UO_841 (O_841,N_14949,N_14755);
and UO_842 (O_842,N_14758,N_14834);
nor UO_843 (O_843,N_14977,N_14924);
nand UO_844 (O_844,N_14920,N_14824);
nand UO_845 (O_845,N_14991,N_14806);
and UO_846 (O_846,N_14843,N_14971);
or UO_847 (O_847,N_14969,N_14818);
and UO_848 (O_848,N_14943,N_14786);
or UO_849 (O_849,N_14755,N_14898);
nor UO_850 (O_850,N_14893,N_14846);
nand UO_851 (O_851,N_14807,N_14800);
and UO_852 (O_852,N_14926,N_14949);
or UO_853 (O_853,N_14795,N_14988);
nand UO_854 (O_854,N_14764,N_14851);
nand UO_855 (O_855,N_14899,N_14764);
nand UO_856 (O_856,N_14785,N_14767);
nor UO_857 (O_857,N_14980,N_14847);
nand UO_858 (O_858,N_14899,N_14871);
or UO_859 (O_859,N_14798,N_14865);
or UO_860 (O_860,N_14761,N_14959);
nand UO_861 (O_861,N_14865,N_14801);
or UO_862 (O_862,N_14940,N_14882);
and UO_863 (O_863,N_14987,N_14926);
or UO_864 (O_864,N_14765,N_14913);
or UO_865 (O_865,N_14837,N_14851);
xnor UO_866 (O_866,N_14777,N_14856);
nand UO_867 (O_867,N_14918,N_14765);
or UO_868 (O_868,N_14951,N_14786);
and UO_869 (O_869,N_14769,N_14845);
and UO_870 (O_870,N_14799,N_14883);
and UO_871 (O_871,N_14924,N_14763);
nor UO_872 (O_872,N_14904,N_14910);
xor UO_873 (O_873,N_14884,N_14830);
nor UO_874 (O_874,N_14989,N_14776);
and UO_875 (O_875,N_14899,N_14753);
or UO_876 (O_876,N_14961,N_14890);
and UO_877 (O_877,N_14991,N_14762);
nor UO_878 (O_878,N_14766,N_14944);
nand UO_879 (O_879,N_14803,N_14983);
nor UO_880 (O_880,N_14892,N_14860);
and UO_881 (O_881,N_14944,N_14775);
and UO_882 (O_882,N_14956,N_14932);
and UO_883 (O_883,N_14892,N_14771);
and UO_884 (O_884,N_14814,N_14869);
nor UO_885 (O_885,N_14869,N_14910);
nor UO_886 (O_886,N_14993,N_14853);
or UO_887 (O_887,N_14788,N_14975);
nand UO_888 (O_888,N_14770,N_14925);
and UO_889 (O_889,N_14990,N_14783);
and UO_890 (O_890,N_14786,N_14871);
or UO_891 (O_891,N_14998,N_14906);
nand UO_892 (O_892,N_14836,N_14797);
and UO_893 (O_893,N_14767,N_14956);
or UO_894 (O_894,N_14775,N_14954);
and UO_895 (O_895,N_14776,N_14983);
or UO_896 (O_896,N_14762,N_14902);
nor UO_897 (O_897,N_14873,N_14997);
and UO_898 (O_898,N_14896,N_14977);
nor UO_899 (O_899,N_14770,N_14893);
and UO_900 (O_900,N_14783,N_14758);
and UO_901 (O_901,N_14761,N_14999);
or UO_902 (O_902,N_14957,N_14853);
nor UO_903 (O_903,N_14929,N_14918);
nand UO_904 (O_904,N_14870,N_14909);
or UO_905 (O_905,N_14888,N_14790);
nand UO_906 (O_906,N_14963,N_14915);
nand UO_907 (O_907,N_14786,N_14833);
and UO_908 (O_908,N_14857,N_14936);
nand UO_909 (O_909,N_14852,N_14959);
and UO_910 (O_910,N_14824,N_14944);
and UO_911 (O_911,N_14882,N_14859);
xor UO_912 (O_912,N_14903,N_14990);
nor UO_913 (O_913,N_14787,N_14816);
or UO_914 (O_914,N_14813,N_14776);
or UO_915 (O_915,N_14897,N_14808);
nor UO_916 (O_916,N_14863,N_14873);
or UO_917 (O_917,N_14780,N_14951);
nor UO_918 (O_918,N_14759,N_14938);
nand UO_919 (O_919,N_14878,N_14869);
or UO_920 (O_920,N_14798,N_14766);
and UO_921 (O_921,N_14976,N_14818);
and UO_922 (O_922,N_14940,N_14902);
or UO_923 (O_923,N_14764,N_14936);
nand UO_924 (O_924,N_14848,N_14883);
or UO_925 (O_925,N_14990,N_14790);
or UO_926 (O_926,N_14958,N_14990);
or UO_927 (O_927,N_14922,N_14862);
nor UO_928 (O_928,N_14956,N_14794);
and UO_929 (O_929,N_14891,N_14982);
and UO_930 (O_930,N_14950,N_14794);
nand UO_931 (O_931,N_14875,N_14945);
nor UO_932 (O_932,N_14953,N_14963);
and UO_933 (O_933,N_14986,N_14965);
nor UO_934 (O_934,N_14953,N_14995);
nor UO_935 (O_935,N_14821,N_14836);
and UO_936 (O_936,N_14830,N_14824);
xor UO_937 (O_937,N_14973,N_14856);
and UO_938 (O_938,N_14789,N_14982);
or UO_939 (O_939,N_14841,N_14765);
nand UO_940 (O_940,N_14821,N_14951);
or UO_941 (O_941,N_14840,N_14837);
nand UO_942 (O_942,N_14848,N_14869);
nand UO_943 (O_943,N_14808,N_14752);
and UO_944 (O_944,N_14990,N_14770);
or UO_945 (O_945,N_14879,N_14802);
nor UO_946 (O_946,N_14857,N_14815);
and UO_947 (O_947,N_14929,N_14881);
nor UO_948 (O_948,N_14990,N_14829);
nor UO_949 (O_949,N_14805,N_14858);
or UO_950 (O_950,N_14992,N_14957);
nand UO_951 (O_951,N_14848,N_14865);
and UO_952 (O_952,N_14759,N_14903);
and UO_953 (O_953,N_14754,N_14853);
and UO_954 (O_954,N_14990,N_14762);
or UO_955 (O_955,N_14882,N_14781);
and UO_956 (O_956,N_14843,N_14752);
nor UO_957 (O_957,N_14978,N_14960);
nand UO_958 (O_958,N_14920,N_14979);
or UO_959 (O_959,N_14901,N_14974);
nor UO_960 (O_960,N_14933,N_14754);
and UO_961 (O_961,N_14994,N_14936);
or UO_962 (O_962,N_14906,N_14938);
nor UO_963 (O_963,N_14791,N_14754);
and UO_964 (O_964,N_14787,N_14755);
or UO_965 (O_965,N_14815,N_14903);
and UO_966 (O_966,N_14834,N_14938);
nand UO_967 (O_967,N_14886,N_14934);
nand UO_968 (O_968,N_14857,N_14949);
nor UO_969 (O_969,N_14759,N_14842);
nor UO_970 (O_970,N_14788,N_14960);
and UO_971 (O_971,N_14783,N_14959);
and UO_972 (O_972,N_14780,N_14817);
or UO_973 (O_973,N_14782,N_14982);
and UO_974 (O_974,N_14962,N_14907);
or UO_975 (O_975,N_14950,N_14903);
and UO_976 (O_976,N_14882,N_14929);
nand UO_977 (O_977,N_14943,N_14940);
nor UO_978 (O_978,N_14944,N_14799);
or UO_979 (O_979,N_14770,N_14984);
and UO_980 (O_980,N_14945,N_14980);
and UO_981 (O_981,N_14751,N_14915);
or UO_982 (O_982,N_14813,N_14755);
nor UO_983 (O_983,N_14895,N_14755);
nor UO_984 (O_984,N_14798,N_14866);
nor UO_985 (O_985,N_14868,N_14774);
nand UO_986 (O_986,N_14859,N_14828);
or UO_987 (O_987,N_14804,N_14882);
and UO_988 (O_988,N_14994,N_14794);
and UO_989 (O_989,N_14839,N_14855);
or UO_990 (O_990,N_14985,N_14848);
nor UO_991 (O_991,N_14969,N_14980);
or UO_992 (O_992,N_14897,N_14981);
or UO_993 (O_993,N_14975,N_14935);
nor UO_994 (O_994,N_14796,N_14986);
and UO_995 (O_995,N_14835,N_14831);
nor UO_996 (O_996,N_14879,N_14948);
and UO_997 (O_997,N_14988,N_14869);
nor UO_998 (O_998,N_14767,N_14802);
nand UO_999 (O_999,N_14829,N_14790);
nor UO_1000 (O_1000,N_14915,N_14941);
nor UO_1001 (O_1001,N_14920,N_14960);
nor UO_1002 (O_1002,N_14886,N_14902);
xor UO_1003 (O_1003,N_14901,N_14762);
or UO_1004 (O_1004,N_14766,N_14913);
nand UO_1005 (O_1005,N_14926,N_14890);
and UO_1006 (O_1006,N_14840,N_14907);
nand UO_1007 (O_1007,N_14981,N_14798);
nor UO_1008 (O_1008,N_14750,N_14777);
nor UO_1009 (O_1009,N_14998,N_14835);
nor UO_1010 (O_1010,N_14757,N_14805);
or UO_1011 (O_1011,N_14776,N_14862);
nand UO_1012 (O_1012,N_14772,N_14906);
and UO_1013 (O_1013,N_14797,N_14750);
nor UO_1014 (O_1014,N_14806,N_14969);
nand UO_1015 (O_1015,N_14830,N_14919);
nand UO_1016 (O_1016,N_14774,N_14750);
nand UO_1017 (O_1017,N_14894,N_14947);
nand UO_1018 (O_1018,N_14917,N_14794);
nand UO_1019 (O_1019,N_14906,N_14953);
or UO_1020 (O_1020,N_14823,N_14786);
or UO_1021 (O_1021,N_14769,N_14778);
nand UO_1022 (O_1022,N_14937,N_14869);
and UO_1023 (O_1023,N_14923,N_14803);
and UO_1024 (O_1024,N_14936,N_14933);
xnor UO_1025 (O_1025,N_14834,N_14932);
or UO_1026 (O_1026,N_14892,N_14959);
nand UO_1027 (O_1027,N_14773,N_14989);
nand UO_1028 (O_1028,N_14975,N_14951);
or UO_1029 (O_1029,N_14949,N_14807);
nor UO_1030 (O_1030,N_14895,N_14904);
nand UO_1031 (O_1031,N_14767,N_14828);
nand UO_1032 (O_1032,N_14752,N_14861);
nor UO_1033 (O_1033,N_14937,N_14961);
and UO_1034 (O_1034,N_14956,N_14877);
nor UO_1035 (O_1035,N_14759,N_14766);
and UO_1036 (O_1036,N_14961,N_14803);
nor UO_1037 (O_1037,N_14853,N_14839);
and UO_1038 (O_1038,N_14825,N_14959);
or UO_1039 (O_1039,N_14958,N_14903);
or UO_1040 (O_1040,N_14859,N_14937);
and UO_1041 (O_1041,N_14848,N_14932);
nand UO_1042 (O_1042,N_14767,N_14751);
and UO_1043 (O_1043,N_14783,N_14861);
xnor UO_1044 (O_1044,N_14759,N_14998);
nor UO_1045 (O_1045,N_14841,N_14843);
or UO_1046 (O_1046,N_14761,N_14974);
xnor UO_1047 (O_1047,N_14976,N_14774);
and UO_1048 (O_1048,N_14875,N_14791);
or UO_1049 (O_1049,N_14790,N_14973);
nand UO_1050 (O_1050,N_14781,N_14754);
nand UO_1051 (O_1051,N_14800,N_14926);
or UO_1052 (O_1052,N_14956,N_14894);
or UO_1053 (O_1053,N_14926,N_14840);
nand UO_1054 (O_1054,N_14928,N_14954);
or UO_1055 (O_1055,N_14850,N_14945);
or UO_1056 (O_1056,N_14852,N_14971);
or UO_1057 (O_1057,N_14823,N_14954);
and UO_1058 (O_1058,N_14816,N_14753);
nand UO_1059 (O_1059,N_14965,N_14791);
or UO_1060 (O_1060,N_14770,N_14801);
nand UO_1061 (O_1061,N_14805,N_14754);
nand UO_1062 (O_1062,N_14932,N_14880);
nand UO_1063 (O_1063,N_14776,N_14795);
nor UO_1064 (O_1064,N_14874,N_14807);
and UO_1065 (O_1065,N_14822,N_14752);
nor UO_1066 (O_1066,N_14808,N_14828);
nor UO_1067 (O_1067,N_14889,N_14970);
nor UO_1068 (O_1068,N_14844,N_14901);
nand UO_1069 (O_1069,N_14801,N_14905);
nand UO_1070 (O_1070,N_14881,N_14846);
or UO_1071 (O_1071,N_14975,N_14799);
or UO_1072 (O_1072,N_14903,N_14951);
and UO_1073 (O_1073,N_14800,N_14825);
nor UO_1074 (O_1074,N_14760,N_14978);
nand UO_1075 (O_1075,N_14946,N_14764);
nor UO_1076 (O_1076,N_14878,N_14768);
nor UO_1077 (O_1077,N_14858,N_14932);
nand UO_1078 (O_1078,N_14883,N_14931);
and UO_1079 (O_1079,N_14985,N_14956);
and UO_1080 (O_1080,N_14935,N_14839);
xor UO_1081 (O_1081,N_14838,N_14847);
nor UO_1082 (O_1082,N_14947,N_14801);
or UO_1083 (O_1083,N_14840,N_14922);
or UO_1084 (O_1084,N_14826,N_14886);
nand UO_1085 (O_1085,N_14813,N_14986);
or UO_1086 (O_1086,N_14978,N_14888);
and UO_1087 (O_1087,N_14756,N_14930);
and UO_1088 (O_1088,N_14821,N_14807);
or UO_1089 (O_1089,N_14948,N_14878);
or UO_1090 (O_1090,N_14826,N_14930);
or UO_1091 (O_1091,N_14934,N_14884);
and UO_1092 (O_1092,N_14817,N_14769);
xor UO_1093 (O_1093,N_14798,N_14922);
and UO_1094 (O_1094,N_14751,N_14936);
nor UO_1095 (O_1095,N_14908,N_14877);
nor UO_1096 (O_1096,N_14810,N_14821);
nor UO_1097 (O_1097,N_14866,N_14890);
nor UO_1098 (O_1098,N_14967,N_14890);
or UO_1099 (O_1099,N_14869,N_14943);
nor UO_1100 (O_1100,N_14824,N_14915);
and UO_1101 (O_1101,N_14939,N_14874);
and UO_1102 (O_1102,N_14964,N_14750);
nand UO_1103 (O_1103,N_14962,N_14871);
or UO_1104 (O_1104,N_14756,N_14758);
nor UO_1105 (O_1105,N_14946,N_14877);
nand UO_1106 (O_1106,N_14868,N_14780);
nand UO_1107 (O_1107,N_14830,N_14943);
or UO_1108 (O_1108,N_14769,N_14907);
nor UO_1109 (O_1109,N_14843,N_14949);
or UO_1110 (O_1110,N_14805,N_14802);
nor UO_1111 (O_1111,N_14788,N_14996);
nand UO_1112 (O_1112,N_14925,N_14776);
and UO_1113 (O_1113,N_14783,N_14960);
or UO_1114 (O_1114,N_14969,N_14878);
and UO_1115 (O_1115,N_14773,N_14886);
nor UO_1116 (O_1116,N_14859,N_14878);
or UO_1117 (O_1117,N_14753,N_14789);
and UO_1118 (O_1118,N_14753,N_14860);
nand UO_1119 (O_1119,N_14806,N_14852);
xnor UO_1120 (O_1120,N_14871,N_14921);
nor UO_1121 (O_1121,N_14869,N_14884);
nor UO_1122 (O_1122,N_14977,N_14755);
nand UO_1123 (O_1123,N_14757,N_14876);
nor UO_1124 (O_1124,N_14844,N_14843);
nand UO_1125 (O_1125,N_14779,N_14914);
and UO_1126 (O_1126,N_14940,N_14847);
nand UO_1127 (O_1127,N_14806,N_14921);
and UO_1128 (O_1128,N_14901,N_14813);
or UO_1129 (O_1129,N_14772,N_14926);
and UO_1130 (O_1130,N_14867,N_14758);
nand UO_1131 (O_1131,N_14890,N_14875);
nand UO_1132 (O_1132,N_14789,N_14981);
or UO_1133 (O_1133,N_14766,N_14821);
and UO_1134 (O_1134,N_14960,N_14910);
or UO_1135 (O_1135,N_14898,N_14987);
nor UO_1136 (O_1136,N_14751,N_14954);
nand UO_1137 (O_1137,N_14944,N_14892);
and UO_1138 (O_1138,N_14855,N_14950);
and UO_1139 (O_1139,N_14965,N_14805);
and UO_1140 (O_1140,N_14848,N_14919);
nor UO_1141 (O_1141,N_14919,N_14911);
nor UO_1142 (O_1142,N_14840,N_14763);
and UO_1143 (O_1143,N_14763,N_14940);
or UO_1144 (O_1144,N_14909,N_14965);
nor UO_1145 (O_1145,N_14890,N_14762);
and UO_1146 (O_1146,N_14999,N_14875);
nor UO_1147 (O_1147,N_14808,N_14827);
nor UO_1148 (O_1148,N_14920,N_14997);
nand UO_1149 (O_1149,N_14853,N_14891);
nor UO_1150 (O_1150,N_14808,N_14926);
or UO_1151 (O_1151,N_14998,N_14968);
nor UO_1152 (O_1152,N_14964,N_14942);
nor UO_1153 (O_1153,N_14888,N_14922);
and UO_1154 (O_1154,N_14772,N_14760);
nor UO_1155 (O_1155,N_14893,N_14943);
nor UO_1156 (O_1156,N_14863,N_14840);
or UO_1157 (O_1157,N_14912,N_14876);
and UO_1158 (O_1158,N_14835,N_14853);
and UO_1159 (O_1159,N_14808,N_14946);
or UO_1160 (O_1160,N_14944,N_14960);
and UO_1161 (O_1161,N_14822,N_14846);
nand UO_1162 (O_1162,N_14851,N_14979);
and UO_1163 (O_1163,N_14958,N_14852);
and UO_1164 (O_1164,N_14755,N_14972);
nand UO_1165 (O_1165,N_14911,N_14796);
and UO_1166 (O_1166,N_14891,N_14799);
nand UO_1167 (O_1167,N_14751,N_14887);
and UO_1168 (O_1168,N_14760,N_14980);
or UO_1169 (O_1169,N_14936,N_14863);
or UO_1170 (O_1170,N_14824,N_14827);
nor UO_1171 (O_1171,N_14916,N_14787);
xor UO_1172 (O_1172,N_14860,N_14769);
or UO_1173 (O_1173,N_14807,N_14894);
nand UO_1174 (O_1174,N_14799,N_14976);
or UO_1175 (O_1175,N_14993,N_14984);
nor UO_1176 (O_1176,N_14849,N_14823);
or UO_1177 (O_1177,N_14981,N_14951);
nand UO_1178 (O_1178,N_14764,N_14755);
and UO_1179 (O_1179,N_14931,N_14860);
nor UO_1180 (O_1180,N_14830,N_14978);
nand UO_1181 (O_1181,N_14916,N_14932);
nor UO_1182 (O_1182,N_14942,N_14918);
or UO_1183 (O_1183,N_14850,N_14918);
nor UO_1184 (O_1184,N_14859,N_14969);
nand UO_1185 (O_1185,N_14850,N_14849);
xor UO_1186 (O_1186,N_14781,N_14848);
nand UO_1187 (O_1187,N_14789,N_14930);
nand UO_1188 (O_1188,N_14768,N_14996);
nand UO_1189 (O_1189,N_14855,N_14940);
nand UO_1190 (O_1190,N_14849,N_14914);
or UO_1191 (O_1191,N_14829,N_14922);
or UO_1192 (O_1192,N_14818,N_14909);
nor UO_1193 (O_1193,N_14986,N_14832);
or UO_1194 (O_1194,N_14804,N_14756);
nand UO_1195 (O_1195,N_14988,N_14960);
or UO_1196 (O_1196,N_14846,N_14879);
xor UO_1197 (O_1197,N_14768,N_14958);
and UO_1198 (O_1198,N_14834,N_14863);
nand UO_1199 (O_1199,N_14766,N_14922);
and UO_1200 (O_1200,N_14851,N_14998);
nor UO_1201 (O_1201,N_14861,N_14788);
and UO_1202 (O_1202,N_14858,N_14935);
and UO_1203 (O_1203,N_14895,N_14860);
or UO_1204 (O_1204,N_14986,N_14815);
nor UO_1205 (O_1205,N_14852,N_14980);
or UO_1206 (O_1206,N_14912,N_14968);
nand UO_1207 (O_1207,N_14943,N_14892);
or UO_1208 (O_1208,N_14779,N_14996);
or UO_1209 (O_1209,N_14835,N_14840);
and UO_1210 (O_1210,N_14931,N_14841);
and UO_1211 (O_1211,N_14893,N_14838);
nor UO_1212 (O_1212,N_14830,N_14972);
or UO_1213 (O_1213,N_14817,N_14842);
or UO_1214 (O_1214,N_14898,N_14970);
and UO_1215 (O_1215,N_14894,N_14886);
nor UO_1216 (O_1216,N_14877,N_14981);
or UO_1217 (O_1217,N_14868,N_14797);
nand UO_1218 (O_1218,N_14764,N_14840);
nor UO_1219 (O_1219,N_14818,N_14844);
and UO_1220 (O_1220,N_14809,N_14961);
nand UO_1221 (O_1221,N_14815,N_14843);
and UO_1222 (O_1222,N_14783,N_14894);
and UO_1223 (O_1223,N_14819,N_14992);
and UO_1224 (O_1224,N_14986,N_14861);
or UO_1225 (O_1225,N_14993,N_14917);
nand UO_1226 (O_1226,N_14884,N_14867);
and UO_1227 (O_1227,N_14873,N_14753);
xor UO_1228 (O_1228,N_14986,N_14776);
xor UO_1229 (O_1229,N_14863,N_14964);
and UO_1230 (O_1230,N_14979,N_14821);
nand UO_1231 (O_1231,N_14772,N_14873);
nand UO_1232 (O_1232,N_14880,N_14779);
or UO_1233 (O_1233,N_14880,N_14827);
nor UO_1234 (O_1234,N_14999,N_14913);
xor UO_1235 (O_1235,N_14929,N_14834);
nor UO_1236 (O_1236,N_14924,N_14830);
and UO_1237 (O_1237,N_14864,N_14871);
and UO_1238 (O_1238,N_14798,N_14983);
and UO_1239 (O_1239,N_14918,N_14953);
nand UO_1240 (O_1240,N_14808,N_14995);
and UO_1241 (O_1241,N_14903,N_14963);
nor UO_1242 (O_1242,N_14952,N_14951);
nand UO_1243 (O_1243,N_14833,N_14971);
nor UO_1244 (O_1244,N_14808,N_14853);
nor UO_1245 (O_1245,N_14880,N_14768);
or UO_1246 (O_1246,N_14831,N_14760);
nand UO_1247 (O_1247,N_14848,N_14964);
nand UO_1248 (O_1248,N_14954,N_14971);
nor UO_1249 (O_1249,N_14799,N_14863);
or UO_1250 (O_1250,N_14915,N_14856);
and UO_1251 (O_1251,N_14889,N_14908);
nor UO_1252 (O_1252,N_14789,N_14905);
nand UO_1253 (O_1253,N_14915,N_14862);
and UO_1254 (O_1254,N_14888,N_14783);
and UO_1255 (O_1255,N_14777,N_14858);
nor UO_1256 (O_1256,N_14787,N_14927);
nand UO_1257 (O_1257,N_14965,N_14864);
nor UO_1258 (O_1258,N_14887,N_14861);
nor UO_1259 (O_1259,N_14793,N_14840);
or UO_1260 (O_1260,N_14750,N_14769);
nor UO_1261 (O_1261,N_14871,N_14815);
nand UO_1262 (O_1262,N_14785,N_14825);
nand UO_1263 (O_1263,N_14927,N_14991);
and UO_1264 (O_1264,N_14777,N_14938);
or UO_1265 (O_1265,N_14917,N_14957);
and UO_1266 (O_1266,N_14847,N_14784);
nand UO_1267 (O_1267,N_14936,N_14991);
nor UO_1268 (O_1268,N_14962,N_14861);
nor UO_1269 (O_1269,N_14789,N_14848);
and UO_1270 (O_1270,N_14850,N_14958);
and UO_1271 (O_1271,N_14880,N_14828);
or UO_1272 (O_1272,N_14785,N_14750);
or UO_1273 (O_1273,N_14919,N_14824);
nand UO_1274 (O_1274,N_14886,N_14769);
or UO_1275 (O_1275,N_14885,N_14982);
nand UO_1276 (O_1276,N_14910,N_14962);
nand UO_1277 (O_1277,N_14800,N_14928);
xnor UO_1278 (O_1278,N_14811,N_14925);
nor UO_1279 (O_1279,N_14907,N_14751);
or UO_1280 (O_1280,N_14976,N_14887);
nor UO_1281 (O_1281,N_14796,N_14967);
or UO_1282 (O_1282,N_14914,N_14895);
nor UO_1283 (O_1283,N_14797,N_14975);
nand UO_1284 (O_1284,N_14797,N_14793);
nand UO_1285 (O_1285,N_14788,N_14913);
and UO_1286 (O_1286,N_14938,N_14983);
nand UO_1287 (O_1287,N_14846,N_14964);
nand UO_1288 (O_1288,N_14852,N_14812);
nor UO_1289 (O_1289,N_14812,N_14890);
or UO_1290 (O_1290,N_14810,N_14847);
nor UO_1291 (O_1291,N_14863,N_14810);
nand UO_1292 (O_1292,N_14904,N_14840);
nand UO_1293 (O_1293,N_14829,N_14851);
and UO_1294 (O_1294,N_14981,N_14860);
nand UO_1295 (O_1295,N_14971,N_14800);
and UO_1296 (O_1296,N_14860,N_14757);
and UO_1297 (O_1297,N_14997,N_14854);
and UO_1298 (O_1298,N_14865,N_14875);
nor UO_1299 (O_1299,N_14824,N_14951);
nand UO_1300 (O_1300,N_14823,N_14869);
and UO_1301 (O_1301,N_14868,N_14906);
or UO_1302 (O_1302,N_14838,N_14864);
nor UO_1303 (O_1303,N_14819,N_14875);
or UO_1304 (O_1304,N_14903,N_14891);
nor UO_1305 (O_1305,N_14867,N_14944);
and UO_1306 (O_1306,N_14816,N_14934);
nand UO_1307 (O_1307,N_14943,N_14756);
or UO_1308 (O_1308,N_14761,N_14799);
and UO_1309 (O_1309,N_14840,N_14829);
or UO_1310 (O_1310,N_14919,N_14953);
or UO_1311 (O_1311,N_14826,N_14993);
nor UO_1312 (O_1312,N_14901,N_14834);
nand UO_1313 (O_1313,N_14799,N_14789);
nand UO_1314 (O_1314,N_14813,N_14903);
or UO_1315 (O_1315,N_14809,N_14902);
and UO_1316 (O_1316,N_14794,N_14811);
or UO_1317 (O_1317,N_14906,N_14918);
or UO_1318 (O_1318,N_14928,N_14771);
or UO_1319 (O_1319,N_14848,N_14993);
or UO_1320 (O_1320,N_14901,N_14794);
xnor UO_1321 (O_1321,N_14946,N_14822);
nor UO_1322 (O_1322,N_14880,N_14862);
and UO_1323 (O_1323,N_14980,N_14786);
and UO_1324 (O_1324,N_14783,N_14984);
nand UO_1325 (O_1325,N_14939,N_14925);
nand UO_1326 (O_1326,N_14937,N_14986);
and UO_1327 (O_1327,N_14931,N_14927);
and UO_1328 (O_1328,N_14977,N_14973);
or UO_1329 (O_1329,N_14849,N_14790);
nand UO_1330 (O_1330,N_14945,N_14882);
nor UO_1331 (O_1331,N_14801,N_14885);
or UO_1332 (O_1332,N_14788,N_14866);
nand UO_1333 (O_1333,N_14911,N_14829);
nand UO_1334 (O_1334,N_14921,N_14855);
and UO_1335 (O_1335,N_14868,N_14941);
xnor UO_1336 (O_1336,N_14895,N_14788);
or UO_1337 (O_1337,N_14802,N_14994);
nor UO_1338 (O_1338,N_14947,N_14772);
nand UO_1339 (O_1339,N_14923,N_14981);
nand UO_1340 (O_1340,N_14918,N_14859);
nor UO_1341 (O_1341,N_14880,N_14781);
and UO_1342 (O_1342,N_14753,N_14985);
nor UO_1343 (O_1343,N_14978,N_14878);
or UO_1344 (O_1344,N_14763,N_14853);
and UO_1345 (O_1345,N_14821,N_14997);
or UO_1346 (O_1346,N_14870,N_14761);
and UO_1347 (O_1347,N_14901,N_14919);
and UO_1348 (O_1348,N_14797,N_14891);
or UO_1349 (O_1349,N_14944,N_14813);
nand UO_1350 (O_1350,N_14984,N_14854);
nor UO_1351 (O_1351,N_14786,N_14877);
nor UO_1352 (O_1352,N_14760,N_14765);
and UO_1353 (O_1353,N_14770,N_14861);
nor UO_1354 (O_1354,N_14991,N_14907);
nand UO_1355 (O_1355,N_14821,N_14966);
and UO_1356 (O_1356,N_14952,N_14761);
or UO_1357 (O_1357,N_14808,N_14935);
nor UO_1358 (O_1358,N_14920,N_14783);
nand UO_1359 (O_1359,N_14839,N_14816);
nor UO_1360 (O_1360,N_14924,N_14864);
nor UO_1361 (O_1361,N_14884,N_14871);
or UO_1362 (O_1362,N_14971,N_14908);
xor UO_1363 (O_1363,N_14906,N_14884);
xor UO_1364 (O_1364,N_14803,N_14884);
xnor UO_1365 (O_1365,N_14835,N_14896);
and UO_1366 (O_1366,N_14963,N_14757);
nand UO_1367 (O_1367,N_14767,N_14954);
and UO_1368 (O_1368,N_14777,N_14983);
nand UO_1369 (O_1369,N_14836,N_14946);
nand UO_1370 (O_1370,N_14859,N_14753);
nand UO_1371 (O_1371,N_14766,N_14900);
nor UO_1372 (O_1372,N_14859,N_14809);
nor UO_1373 (O_1373,N_14901,N_14843);
nand UO_1374 (O_1374,N_14838,N_14961);
and UO_1375 (O_1375,N_14790,N_14885);
and UO_1376 (O_1376,N_14830,N_14957);
nand UO_1377 (O_1377,N_14884,N_14890);
nand UO_1378 (O_1378,N_14942,N_14834);
nor UO_1379 (O_1379,N_14750,N_14955);
nor UO_1380 (O_1380,N_14812,N_14903);
nand UO_1381 (O_1381,N_14894,N_14839);
or UO_1382 (O_1382,N_14756,N_14946);
and UO_1383 (O_1383,N_14990,N_14871);
and UO_1384 (O_1384,N_14883,N_14998);
nor UO_1385 (O_1385,N_14913,N_14792);
nand UO_1386 (O_1386,N_14966,N_14907);
and UO_1387 (O_1387,N_14756,N_14945);
nand UO_1388 (O_1388,N_14874,N_14758);
or UO_1389 (O_1389,N_14877,N_14774);
nor UO_1390 (O_1390,N_14808,N_14985);
or UO_1391 (O_1391,N_14897,N_14922);
nand UO_1392 (O_1392,N_14940,N_14824);
or UO_1393 (O_1393,N_14848,N_14884);
and UO_1394 (O_1394,N_14958,N_14833);
nor UO_1395 (O_1395,N_14941,N_14770);
and UO_1396 (O_1396,N_14960,N_14877);
nor UO_1397 (O_1397,N_14935,N_14763);
or UO_1398 (O_1398,N_14765,N_14829);
or UO_1399 (O_1399,N_14894,N_14904);
nor UO_1400 (O_1400,N_14978,N_14811);
nor UO_1401 (O_1401,N_14828,N_14784);
nand UO_1402 (O_1402,N_14986,N_14804);
or UO_1403 (O_1403,N_14845,N_14941);
nand UO_1404 (O_1404,N_14854,N_14925);
or UO_1405 (O_1405,N_14816,N_14883);
xor UO_1406 (O_1406,N_14813,N_14940);
and UO_1407 (O_1407,N_14911,N_14922);
nand UO_1408 (O_1408,N_14771,N_14808);
and UO_1409 (O_1409,N_14909,N_14931);
or UO_1410 (O_1410,N_14750,N_14923);
nand UO_1411 (O_1411,N_14943,N_14938);
nor UO_1412 (O_1412,N_14865,N_14960);
or UO_1413 (O_1413,N_14911,N_14861);
nor UO_1414 (O_1414,N_14943,N_14809);
nor UO_1415 (O_1415,N_14975,N_14984);
nand UO_1416 (O_1416,N_14896,N_14833);
and UO_1417 (O_1417,N_14868,N_14888);
nand UO_1418 (O_1418,N_14965,N_14890);
nand UO_1419 (O_1419,N_14951,N_14916);
nand UO_1420 (O_1420,N_14926,N_14956);
nand UO_1421 (O_1421,N_14887,N_14813);
or UO_1422 (O_1422,N_14765,N_14843);
nor UO_1423 (O_1423,N_14788,N_14905);
and UO_1424 (O_1424,N_14969,N_14925);
nor UO_1425 (O_1425,N_14785,N_14977);
and UO_1426 (O_1426,N_14753,N_14900);
or UO_1427 (O_1427,N_14942,N_14774);
or UO_1428 (O_1428,N_14874,N_14928);
and UO_1429 (O_1429,N_14828,N_14795);
nand UO_1430 (O_1430,N_14936,N_14959);
nand UO_1431 (O_1431,N_14911,N_14758);
nand UO_1432 (O_1432,N_14988,N_14948);
nand UO_1433 (O_1433,N_14762,N_14962);
nor UO_1434 (O_1434,N_14868,N_14782);
xnor UO_1435 (O_1435,N_14865,N_14998);
nand UO_1436 (O_1436,N_14957,N_14914);
and UO_1437 (O_1437,N_14932,N_14897);
nand UO_1438 (O_1438,N_14788,N_14801);
nor UO_1439 (O_1439,N_14773,N_14935);
and UO_1440 (O_1440,N_14890,N_14796);
nand UO_1441 (O_1441,N_14798,N_14769);
xor UO_1442 (O_1442,N_14793,N_14851);
nand UO_1443 (O_1443,N_14961,N_14776);
nor UO_1444 (O_1444,N_14840,N_14979);
or UO_1445 (O_1445,N_14950,N_14994);
nor UO_1446 (O_1446,N_14760,N_14942);
nand UO_1447 (O_1447,N_14843,N_14855);
and UO_1448 (O_1448,N_14773,N_14966);
or UO_1449 (O_1449,N_14853,N_14870);
nand UO_1450 (O_1450,N_14784,N_14917);
or UO_1451 (O_1451,N_14801,N_14822);
nand UO_1452 (O_1452,N_14957,N_14760);
nor UO_1453 (O_1453,N_14909,N_14751);
or UO_1454 (O_1454,N_14759,N_14975);
nand UO_1455 (O_1455,N_14938,N_14808);
and UO_1456 (O_1456,N_14936,N_14819);
nor UO_1457 (O_1457,N_14753,N_14820);
or UO_1458 (O_1458,N_14764,N_14857);
and UO_1459 (O_1459,N_14781,N_14767);
nor UO_1460 (O_1460,N_14905,N_14934);
and UO_1461 (O_1461,N_14964,N_14999);
nor UO_1462 (O_1462,N_14832,N_14890);
or UO_1463 (O_1463,N_14982,N_14896);
nor UO_1464 (O_1464,N_14966,N_14824);
nor UO_1465 (O_1465,N_14789,N_14757);
xor UO_1466 (O_1466,N_14950,N_14930);
xor UO_1467 (O_1467,N_14861,N_14798);
or UO_1468 (O_1468,N_14968,N_14796);
and UO_1469 (O_1469,N_14963,N_14881);
and UO_1470 (O_1470,N_14892,N_14991);
nand UO_1471 (O_1471,N_14871,N_14801);
nor UO_1472 (O_1472,N_14925,N_14812);
nand UO_1473 (O_1473,N_14938,N_14788);
or UO_1474 (O_1474,N_14997,N_14857);
or UO_1475 (O_1475,N_14854,N_14971);
and UO_1476 (O_1476,N_14756,N_14986);
xor UO_1477 (O_1477,N_14909,N_14837);
nand UO_1478 (O_1478,N_14822,N_14839);
nor UO_1479 (O_1479,N_14903,N_14872);
nand UO_1480 (O_1480,N_14863,N_14793);
nor UO_1481 (O_1481,N_14751,N_14888);
and UO_1482 (O_1482,N_14765,N_14844);
nand UO_1483 (O_1483,N_14949,N_14886);
nor UO_1484 (O_1484,N_14893,N_14960);
xnor UO_1485 (O_1485,N_14808,N_14990);
nand UO_1486 (O_1486,N_14784,N_14808);
and UO_1487 (O_1487,N_14802,N_14950);
nor UO_1488 (O_1488,N_14902,N_14816);
nand UO_1489 (O_1489,N_14771,N_14904);
or UO_1490 (O_1490,N_14908,N_14852);
and UO_1491 (O_1491,N_14817,N_14776);
or UO_1492 (O_1492,N_14870,N_14860);
or UO_1493 (O_1493,N_14839,N_14950);
nor UO_1494 (O_1494,N_14874,N_14994);
or UO_1495 (O_1495,N_14884,N_14815);
nand UO_1496 (O_1496,N_14850,N_14919);
nor UO_1497 (O_1497,N_14875,N_14802);
or UO_1498 (O_1498,N_14956,N_14876);
or UO_1499 (O_1499,N_14788,N_14803);
or UO_1500 (O_1500,N_14930,N_14867);
nand UO_1501 (O_1501,N_14970,N_14793);
and UO_1502 (O_1502,N_14965,N_14798);
nand UO_1503 (O_1503,N_14806,N_14871);
nand UO_1504 (O_1504,N_14815,N_14870);
nand UO_1505 (O_1505,N_14909,N_14752);
nor UO_1506 (O_1506,N_14944,N_14818);
nand UO_1507 (O_1507,N_14787,N_14778);
and UO_1508 (O_1508,N_14772,N_14837);
nand UO_1509 (O_1509,N_14889,N_14841);
and UO_1510 (O_1510,N_14906,N_14977);
nand UO_1511 (O_1511,N_14904,N_14821);
nand UO_1512 (O_1512,N_14962,N_14946);
xor UO_1513 (O_1513,N_14846,N_14792);
nor UO_1514 (O_1514,N_14757,N_14978);
nand UO_1515 (O_1515,N_14877,N_14950);
and UO_1516 (O_1516,N_14787,N_14960);
xnor UO_1517 (O_1517,N_14834,N_14814);
nand UO_1518 (O_1518,N_14905,N_14758);
or UO_1519 (O_1519,N_14782,N_14892);
and UO_1520 (O_1520,N_14931,N_14921);
nand UO_1521 (O_1521,N_14861,N_14972);
or UO_1522 (O_1522,N_14987,N_14984);
nand UO_1523 (O_1523,N_14878,N_14980);
nand UO_1524 (O_1524,N_14890,N_14925);
or UO_1525 (O_1525,N_14940,N_14917);
and UO_1526 (O_1526,N_14813,N_14810);
nand UO_1527 (O_1527,N_14959,N_14868);
nand UO_1528 (O_1528,N_14759,N_14774);
and UO_1529 (O_1529,N_14766,N_14894);
nor UO_1530 (O_1530,N_14941,N_14931);
nand UO_1531 (O_1531,N_14927,N_14894);
or UO_1532 (O_1532,N_14885,N_14851);
xor UO_1533 (O_1533,N_14927,N_14945);
and UO_1534 (O_1534,N_14766,N_14959);
or UO_1535 (O_1535,N_14957,N_14889);
or UO_1536 (O_1536,N_14999,N_14796);
nor UO_1537 (O_1537,N_14800,N_14995);
xor UO_1538 (O_1538,N_14933,N_14756);
nand UO_1539 (O_1539,N_14957,N_14882);
and UO_1540 (O_1540,N_14797,N_14940);
and UO_1541 (O_1541,N_14945,N_14942);
nand UO_1542 (O_1542,N_14891,N_14871);
and UO_1543 (O_1543,N_14895,N_14776);
nor UO_1544 (O_1544,N_14938,N_14953);
nor UO_1545 (O_1545,N_14836,N_14816);
nor UO_1546 (O_1546,N_14824,N_14911);
and UO_1547 (O_1547,N_14987,N_14978);
or UO_1548 (O_1548,N_14943,N_14772);
or UO_1549 (O_1549,N_14814,N_14882);
nand UO_1550 (O_1550,N_14780,N_14826);
nor UO_1551 (O_1551,N_14791,N_14996);
and UO_1552 (O_1552,N_14971,N_14838);
nor UO_1553 (O_1553,N_14913,N_14853);
nor UO_1554 (O_1554,N_14931,N_14874);
nand UO_1555 (O_1555,N_14884,N_14911);
nand UO_1556 (O_1556,N_14756,N_14979);
or UO_1557 (O_1557,N_14806,N_14880);
nand UO_1558 (O_1558,N_14982,N_14900);
nor UO_1559 (O_1559,N_14968,N_14813);
xnor UO_1560 (O_1560,N_14910,N_14810);
nand UO_1561 (O_1561,N_14779,N_14861);
nand UO_1562 (O_1562,N_14995,N_14984);
nand UO_1563 (O_1563,N_14953,N_14864);
nor UO_1564 (O_1564,N_14963,N_14969);
or UO_1565 (O_1565,N_14953,N_14802);
nand UO_1566 (O_1566,N_14927,N_14907);
and UO_1567 (O_1567,N_14841,N_14969);
and UO_1568 (O_1568,N_14888,N_14821);
nor UO_1569 (O_1569,N_14939,N_14754);
or UO_1570 (O_1570,N_14827,N_14842);
and UO_1571 (O_1571,N_14906,N_14778);
nor UO_1572 (O_1572,N_14926,N_14878);
or UO_1573 (O_1573,N_14756,N_14844);
and UO_1574 (O_1574,N_14882,N_14983);
and UO_1575 (O_1575,N_14898,N_14810);
and UO_1576 (O_1576,N_14750,N_14835);
and UO_1577 (O_1577,N_14892,N_14993);
and UO_1578 (O_1578,N_14903,N_14841);
and UO_1579 (O_1579,N_14992,N_14792);
nand UO_1580 (O_1580,N_14965,N_14990);
or UO_1581 (O_1581,N_14789,N_14991);
and UO_1582 (O_1582,N_14990,N_14944);
or UO_1583 (O_1583,N_14934,N_14777);
or UO_1584 (O_1584,N_14992,N_14983);
or UO_1585 (O_1585,N_14836,N_14851);
nor UO_1586 (O_1586,N_14880,N_14935);
nor UO_1587 (O_1587,N_14874,N_14904);
and UO_1588 (O_1588,N_14831,N_14985);
and UO_1589 (O_1589,N_14818,N_14946);
nand UO_1590 (O_1590,N_14928,N_14784);
nor UO_1591 (O_1591,N_14825,N_14907);
or UO_1592 (O_1592,N_14984,N_14808);
nor UO_1593 (O_1593,N_14993,N_14796);
and UO_1594 (O_1594,N_14781,N_14896);
xor UO_1595 (O_1595,N_14912,N_14866);
xor UO_1596 (O_1596,N_14926,N_14844);
or UO_1597 (O_1597,N_14840,N_14873);
or UO_1598 (O_1598,N_14985,N_14791);
or UO_1599 (O_1599,N_14791,N_14909);
and UO_1600 (O_1600,N_14882,N_14914);
nand UO_1601 (O_1601,N_14942,N_14888);
and UO_1602 (O_1602,N_14905,N_14804);
and UO_1603 (O_1603,N_14912,N_14969);
and UO_1604 (O_1604,N_14916,N_14931);
nor UO_1605 (O_1605,N_14810,N_14909);
nand UO_1606 (O_1606,N_14762,N_14997);
nand UO_1607 (O_1607,N_14872,N_14804);
xor UO_1608 (O_1608,N_14932,N_14907);
or UO_1609 (O_1609,N_14862,N_14819);
nor UO_1610 (O_1610,N_14948,N_14962);
or UO_1611 (O_1611,N_14919,N_14820);
nand UO_1612 (O_1612,N_14909,N_14803);
or UO_1613 (O_1613,N_14797,N_14831);
and UO_1614 (O_1614,N_14787,N_14774);
xor UO_1615 (O_1615,N_14788,N_14818);
nand UO_1616 (O_1616,N_14870,N_14876);
nor UO_1617 (O_1617,N_14993,N_14903);
and UO_1618 (O_1618,N_14907,N_14981);
nor UO_1619 (O_1619,N_14889,N_14789);
and UO_1620 (O_1620,N_14817,N_14774);
nor UO_1621 (O_1621,N_14764,N_14994);
and UO_1622 (O_1622,N_14883,N_14914);
and UO_1623 (O_1623,N_14996,N_14950);
nor UO_1624 (O_1624,N_14762,N_14895);
nand UO_1625 (O_1625,N_14997,N_14837);
nand UO_1626 (O_1626,N_14752,N_14866);
xnor UO_1627 (O_1627,N_14973,N_14885);
and UO_1628 (O_1628,N_14849,N_14802);
or UO_1629 (O_1629,N_14766,N_14832);
xnor UO_1630 (O_1630,N_14835,N_14933);
nor UO_1631 (O_1631,N_14753,N_14832);
or UO_1632 (O_1632,N_14840,N_14834);
nor UO_1633 (O_1633,N_14889,N_14778);
nand UO_1634 (O_1634,N_14890,N_14784);
and UO_1635 (O_1635,N_14901,N_14783);
nor UO_1636 (O_1636,N_14849,N_14826);
nand UO_1637 (O_1637,N_14916,N_14776);
xnor UO_1638 (O_1638,N_14899,N_14911);
and UO_1639 (O_1639,N_14854,N_14980);
and UO_1640 (O_1640,N_14993,N_14947);
nor UO_1641 (O_1641,N_14862,N_14914);
nand UO_1642 (O_1642,N_14960,N_14894);
or UO_1643 (O_1643,N_14893,N_14986);
nor UO_1644 (O_1644,N_14868,N_14993);
and UO_1645 (O_1645,N_14956,N_14961);
or UO_1646 (O_1646,N_14771,N_14963);
or UO_1647 (O_1647,N_14925,N_14941);
nor UO_1648 (O_1648,N_14874,N_14888);
and UO_1649 (O_1649,N_14850,N_14852);
nor UO_1650 (O_1650,N_14882,N_14819);
or UO_1651 (O_1651,N_14759,N_14974);
or UO_1652 (O_1652,N_14976,N_14846);
xor UO_1653 (O_1653,N_14965,N_14987);
nand UO_1654 (O_1654,N_14808,N_14819);
and UO_1655 (O_1655,N_14763,N_14923);
xnor UO_1656 (O_1656,N_14947,N_14760);
or UO_1657 (O_1657,N_14937,N_14834);
nor UO_1658 (O_1658,N_14991,N_14799);
and UO_1659 (O_1659,N_14866,N_14750);
and UO_1660 (O_1660,N_14995,N_14876);
nor UO_1661 (O_1661,N_14766,N_14925);
xnor UO_1662 (O_1662,N_14753,N_14847);
or UO_1663 (O_1663,N_14941,N_14946);
nand UO_1664 (O_1664,N_14910,N_14832);
or UO_1665 (O_1665,N_14956,N_14882);
nand UO_1666 (O_1666,N_14793,N_14980);
and UO_1667 (O_1667,N_14883,N_14858);
or UO_1668 (O_1668,N_14860,N_14991);
or UO_1669 (O_1669,N_14999,N_14832);
or UO_1670 (O_1670,N_14843,N_14941);
nor UO_1671 (O_1671,N_14756,N_14871);
and UO_1672 (O_1672,N_14931,N_14972);
nor UO_1673 (O_1673,N_14852,N_14853);
nor UO_1674 (O_1674,N_14927,N_14941);
nand UO_1675 (O_1675,N_14895,N_14770);
nor UO_1676 (O_1676,N_14959,N_14828);
nand UO_1677 (O_1677,N_14970,N_14794);
xor UO_1678 (O_1678,N_14931,N_14798);
nand UO_1679 (O_1679,N_14943,N_14958);
nand UO_1680 (O_1680,N_14914,N_14805);
or UO_1681 (O_1681,N_14952,N_14921);
nand UO_1682 (O_1682,N_14964,N_14974);
and UO_1683 (O_1683,N_14806,N_14983);
nand UO_1684 (O_1684,N_14854,N_14765);
nor UO_1685 (O_1685,N_14965,N_14792);
and UO_1686 (O_1686,N_14805,N_14943);
and UO_1687 (O_1687,N_14841,N_14807);
and UO_1688 (O_1688,N_14821,N_14854);
or UO_1689 (O_1689,N_14996,N_14825);
or UO_1690 (O_1690,N_14990,N_14961);
nand UO_1691 (O_1691,N_14950,N_14764);
or UO_1692 (O_1692,N_14867,N_14891);
nor UO_1693 (O_1693,N_14962,N_14797);
or UO_1694 (O_1694,N_14978,N_14798);
nand UO_1695 (O_1695,N_14891,N_14950);
xor UO_1696 (O_1696,N_14992,N_14840);
nor UO_1697 (O_1697,N_14801,N_14785);
nor UO_1698 (O_1698,N_14775,N_14920);
or UO_1699 (O_1699,N_14817,N_14798);
or UO_1700 (O_1700,N_14924,N_14792);
and UO_1701 (O_1701,N_14837,N_14880);
nand UO_1702 (O_1702,N_14966,N_14900);
nand UO_1703 (O_1703,N_14784,N_14882);
or UO_1704 (O_1704,N_14952,N_14993);
or UO_1705 (O_1705,N_14969,N_14898);
nor UO_1706 (O_1706,N_14965,N_14945);
or UO_1707 (O_1707,N_14962,N_14800);
and UO_1708 (O_1708,N_14927,N_14823);
and UO_1709 (O_1709,N_14981,N_14866);
nor UO_1710 (O_1710,N_14787,N_14956);
and UO_1711 (O_1711,N_14789,N_14886);
nand UO_1712 (O_1712,N_14831,N_14758);
and UO_1713 (O_1713,N_14912,N_14768);
nand UO_1714 (O_1714,N_14825,N_14982);
and UO_1715 (O_1715,N_14946,N_14997);
nor UO_1716 (O_1716,N_14953,N_14813);
nand UO_1717 (O_1717,N_14791,N_14772);
nand UO_1718 (O_1718,N_14834,N_14753);
and UO_1719 (O_1719,N_14758,N_14981);
and UO_1720 (O_1720,N_14954,N_14861);
nand UO_1721 (O_1721,N_14812,N_14780);
nand UO_1722 (O_1722,N_14972,N_14803);
and UO_1723 (O_1723,N_14917,N_14766);
or UO_1724 (O_1724,N_14799,N_14936);
nor UO_1725 (O_1725,N_14786,N_14845);
or UO_1726 (O_1726,N_14903,N_14858);
nor UO_1727 (O_1727,N_14936,N_14895);
or UO_1728 (O_1728,N_14997,N_14763);
and UO_1729 (O_1729,N_14972,N_14884);
and UO_1730 (O_1730,N_14896,N_14933);
and UO_1731 (O_1731,N_14983,N_14859);
or UO_1732 (O_1732,N_14808,N_14997);
and UO_1733 (O_1733,N_14933,N_14876);
nand UO_1734 (O_1734,N_14784,N_14801);
nor UO_1735 (O_1735,N_14818,N_14987);
nor UO_1736 (O_1736,N_14804,N_14939);
nor UO_1737 (O_1737,N_14916,N_14948);
nor UO_1738 (O_1738,N_14957,N_14753);
nand UO_1739 (O_1739,N_14965,N_14994);
nor UO_1740 (O_1740,N_14896,N_14783);
or UO_1741 (O_1741,N_14948,N_14931);
nor UO_1742 (O_1742,N_14971,N_14997);
and UO_1743 (O_1743,N_14823,N_14877);
nor UO_1744 (O_1744,N_14813,N_14921);
and UO_1745 (O_1745,N_14898,N_14854);
or UO_1746 (O_1746,N_14999,N_14967);
nand UO_1747 (O_1747,N_14919,N_14861);
or UO_1748 (O_1748,N_14934,N_14954);
and UO_1749 (O_1749,N_14966,N_14947);
or UO_1750 (O_1750,N_14862,N_14778);
nand UO_1751 (O_1751,N_14868,N_14831);
and UO_1752 (O_1752,N_14872,N_14992);
or UO_1753 (O_1753,N_14932,N_14943);
nand UO_1754 (O_1754,N_14852,N_14923);
or UO_1755 (O_1755,N_14797,N_14949);
and UO_1756 (O_1756,N_14996,N_14917);
and UO_1757 (O_1757,N_14764,N_14867);
nand UO_1758 (O_1758,N_14842,N_14980);
and UO_1759 (O_1759,N_14852,N_14802);
nor UO_1760 (O_1760,N_14828,N_14863);
nor UO_1761 (O_1761,N_14774,N_14795);
and UO_1762 (O_1762,N_14957,N_14911);
or UO_1763 (O_1763,N_14830,N_14926);
nor UO_1764 (O_1764,N_14890,N_14979);
nand UO_1765 (O_1765,N_14871,N_14910);
nor UO_1766 (O_1766,N_14864,N_14918);
nand UO_1767 (O_1767,N_14802,N_14785);
nor UO_1768 (O_1768,N_14757,N_14800);
nor UO_1769 (O_1769,N_14995,N_14944);
and UO_1770 (O_1770,N_14913,N_14946);
or UO_1771 (O_1771,N_14894,N_14912);
or UO_1772 (O_1772,N_14758,N_14962);
or UO_1773 (O_1773,N_14826,N_14883);
or UO_1774 (O_1774,N_14916,N_14968);
and UO_1775 (O_1775,N_14948,N_14881);
and UO_1776 (O_1776,N_14871,N_14993);
and UO_1777 (O_1777,N_14969,N_14849);
nor UO_1778 (O_1778,N_14985,N_14779);
or UO_1779 (O_1779,N_14971,N_14986);
nor UO_1780 (O_1780,N_14970,N_14905);
and UO_1781 (O_1781,N_14807,N_14992);
and UO_1782 (O_1782,N_14919,N_14807);
nor UO_1783 (O_1783,N_14968,N_14892);
and UO_1784 (O_1784,N_14944,N_14764);
and UO_1785 (O_1785,N_14767,N_14969);
nor UO_1786 (O_1786,N_14760,N_14956);
or UO_1787 (O_1787,N_14929,N_14832);
and UO_1788 (O_1788,N_14817,N_14811);
or UO_1789 (O_1789,N_14766,N_14927);
xnor UO_1790 (O_1790,N_14775,N_14816);
nor UO_1791 (O_1791,N_14778,N_14920);
nand UO_1792 (O_1792,N_14950,N_14901);
xor UO_1793 (O_1793,N_14932,N_14893);
nand UO_1794 (O_1794,N_14774,N_14969);
or UO_1795 (O_1795,N_14981,N_14756);
nand UO_1796 (O_1796,N_14926,N_14836);
and UO_1797 (O_1797,N_14931,N_14946);
or UO_1798 (O_1798,N_14771,N_14858);
or UO_1799 (O_1799,N_14817,N_14840);
and UO_1800 (O_1800,N_14798,N_14894);
nand UO_1801 (O_1801,N_14965,N_14978);
and UO_1802 (O_1802,N_14979,N_14764);
nand UO_1803 (O_1803,N_14999,N_14972);
nor UO_1804 (O_1804,N_14821,N_14994);
or UO_1805 (O_1805,N_14884,N_14904);
nand UO_1806 (O_1806,N_14765,N_14880);
nand UO_1807 (O_1807,N_14979,N_14858);
nor UO_1808 (O_1808,N_14894,N_14806);
nand UO_1809 (O_1809,N_14926,N_14875);
nand UO_1810 (O_1810,N_14938,N_14785);
nor UO_1811 (O_1811,N_14874,N_14772);
nand UO_1812 (O_1812,N_14760,N_14898);
nor UO_1813 (O_1813,N_14763,N_14981);
or UO_1814 (O_1814,N_14964,N_14916);
or UO_1815 (O_1815,N_14757,N_14918);
and UO_1816 (O_1816,N_14944,N_14875);
and UO_1817 (O_1817,N_14945,N_14813);
nand UO_1818 (O_1818,N_14811,N_14808);
and UO_1819 (O_1819,N_14751,N_14818);
nand UO_1820 (O_1820,N_14899,N_14837);
or UO_1821 (O_1821,N_14777,N_14844);
and UO_1822 (O_1822,N_14998,N_14928);
xor UO_1823 (O_1823,N_14858,N_14764);
nand UO_1824 (O_1824,N_14978,N_14796);
or UO_1825 (O_1825,N_14939,N_14986);
or UO_1826 (O_1826,N_14927,N_14850);
or UO_1827 (O_1827,N_14900,N_14883);
or UO_1828 (O_1828,N_14761,N_14998);
nand UO_1829 (O_1829,N_14783,N_14751);
or UO_1830 (O_1830,N_14751,N_14931);
and UO_1831 (O_1831,N_14821,N_14953);
or UO_1832 (O_1832,N_14850,N_14810);
nor UO_1833 (O_1833,N_14817,N_14964);
or UO_1834 (O_1834,N_14786,N_14858);
nor UO_1835 (O_1835,N_14841,N_14771);
nor UO_1836 (O_1836,N_14846,N_14801);
and UO_1837 (O_1837,N_14803,N_14874);
nand UO_1838 (O_1838,N_14849,N_14933);
or UO_1839 (O_1839,N_14845,N_14754);
and UO_1840 (O_1840,N_14961,N_14841);
xnor UO_1841 (O_1841,N_14937,N_14956);
or UO_1842 (O_1842,N_14943,N_14823);
xnor UO_1843 (O_1843,N_14813,N_14870);
and UO_1844 (O_1844,N_14923,N_14844);
nand UO_1845 (O_1845,N_14784,N_14834);
or UO_1846 (O_1846,N_14955,N_14936);
nor UO_1847 (O_1847,N_14941,N_14788);
nand UO_1848 (O_1848,N_14947,N_14858);
or UO_1849 (O_1849,N_14821,N_14943);
nand UO_1850 (O_1850,N_14772,N_14934);
nand UO_1851 (O_1851,N_14852,N_14987);
nand UO_1852 (O_1852,N_14989,N_14874);
or UO_1853 (O_1853,N_14937,N_14987);
and UO_1854 (O_1854,N_14901,N_14918);
and UO_1855 (O_1855,N_14781,N_14750);
or UO_1856 (O_1856,N_14904,N_14882);
nor UO_1857 (O_1857,N_14992,N_14933);
and UO_1858 (O_1858,N_14788,N_14780);
nand UO_1859 (O_1859,N_14897,N_14988);
or UO_1860 (O_1860,N_14873,N_14870);
nor UO_1861 (O_1861,N_14869,N_14920);
nor UO_1862 (O_1862,N_14945,N_14915);
or UO_1863 (O_1863,N_14857,N_14904);
and UO_1864 (O_1864,N_14863,N_14768);
or UO_1865 (O_1865,N_14910,N_14926);
nor UO_1866 (O_1866,N_14790,N_14823);
nor UO_1867 (O_1867,N_14996,N_14838);
and UO_1868 (O_1868,N_14911,N_14994);
and UO_1869 (O_1869,N_14763,N_14807);
or UO_1870 (O_1870,N_14766,N_14942);
nor UO_1871 (O_1871,N_14910,N_14780);
and UO_1872 (O_1872,N_14863,N_14912);
nand UO_1873 (O_1873,N_14821,N_14964);
nand UO_1874 (O_1874,N_14891,N_14837);
or UO_1875 (O_1875,N_14816,N_14994);
or UO_1876 (O_1876,N_14813,N_14758);
nand UO_1877 (O_1877,N_14837,N_14950);
nor UO_1878 (O_1878,N_14902,N_14993);
xnor UO_1879 (O_1879,N_14802,N_14841);
nor UO_1880 (O_1880,N_14963,N_14770);
and UO_1881 (O_1881,N_14816,N_14763);
or UO_1882 (O_1882,N_14975,N_14848);
nand UO_1883 (O_1883,N_14801,N_14897);
or UO_1884 (O_1884,N_14912,N_14874);
and UO_1885 (O_1885,N_14832,N_14917);
or UO_1886 (O_1886,N_14871,N_14918);
and UO_1887 (O_1887,N_14868,N_14851);
xor UO_1888 (O_1888,N_14972,N_14990);
nand UO_1889 (O_1889,N_14956,N_14820);
nand UO_1890 (O_1890,N_14923,N_14811);
nor UO_1891 (O_1891,N_14907,N_14894);
or UO_1892 (O_1892,N_14899,N_14793);
and UO_1893 (O_1893,N_14801,N_14793);
or UO_1894 (O_1894,N_14867,N_14783);
nand UO_1895 (O_1895,N_14901,N_14849);
nand UO_1896 (O_1896,N_14803,N_14970);
nand UO_1897 (O_1897,N_14784,N_14772);
and UO_1898 (O_1898,N_14923,N_14925);
or UO_1899 (O_1899,N_14787,N_14965);
nand UO_1900 (O_1900,N_14969,N_14860);
or UO_1901 (O_1901,N_14754,N_14807);
nand UO_1902 (O_1902,N_14883,N_14797);
nand UO_1903 (O_1903,N_14845,N_14981);
and UO_1904 (O_1904,N_14998,N_14980);
or UO_1905 (O_1905,N_14891,N_14769);
and UO_1906 (O_1906,N_14836,N_14882);
and UO_1907 (O_1907,N_14946,N_14821);
nand UO_1908 (O_1908,N_14933,N_14966);
or UO_1909 (O_1909,N_14774,N_14929);
nand UO_1910 (O_1910,N_14926,N_14792);
nor UO_1911 (O_1911,N_14959,N_14893);
and UO_1912 (O_1912,N_14837,N_14766);
nor UO_1913 (O_1913,N_14761,N_14992);
and UO_1914 (O_1914,N_14909,N_14785);
nor UO_1915 (O_1915,N_14828,N_14857);
nand UO_1916 (O_1916,N_14925,N_14906);
or UO_1917 (O_1917,N_14804,N_14783);
and UO_1918 (O_1918,N_14907,N_14822);
or UO_1919 (O_1919,N_14887,N_14871);
and UO_1920 (O_1920,N_14974,N_14904);
nand UO_1921 (O_1921,N_14985,N_14813);
nand UO_1922 (O_1922,N_14769,N_14861);
or UO_1923 (O_1923,N_14848,N_14914);
or UO_1924 (O_1924,N_14852,N_14930);
nand UO_1925 (O_1925,N_14871,N_14869);
and UO_1926 (O_1926,N_14900,N_14960);
nor UO_1927 (O_1927,N_14919,N_14783);
nor UO_1928 (O_1928,N_14930,N_14792);
and UO_1929 (O_1929,N_14880,N_14851);
nor UO_1930 (O_1930,N_14866,N_14880);
and UO_1931 (O_1931,N_14767,N_14981);
and UO_1932 (O_1932,N_14935,N_14853);
xor UO_1933 (O_1933,N_14752,N_14915);
and UO_1934 (O_1934,N_14791,N_14846);
and UO_1935 (O_1935,N_14894,N_14819);
nor UO_1936 (O_1936,N_14953,N_14769);
and UO_1937 (O_1937,N_14881,N_14845);
or UO_1938 (O_1938,N_14759,N_14996);
nor UO_1939 (O_1939,N_14835,N_14803);
and UO_1940 (O_1940,N_14803,N_14850);
nand UO_1941 (O_1941,N_14868,N_14820);
nor UO_1942 (O_1942,N_14781,N_14870);
and UO_1943 (O_1943,N_14863,N_14963);
and UO_1944 (O_1944,N_14845,N_14802);
nor UO_1945 (O_1945,N_14924,N_14767);
or UO_1946 (O_1946,N_14825,N_14832);
or UO_1947 (O_1947,N_14907,N_14888);
and UO_1948 (O_1948,N_14977,N_14818);
nand UO_1949 (O_1949,N_14848,N_14836);
and UO_1950 (O_1950,N_14951,N_14879);
nor UO_1951 (O_1951,N_14846,N_14764);
nor UO_1952 (O_1952,N_14841,N_14831);
nor UO_1953 (O_1953,N_14940,N_14852);
nor UO_1954 (O_1954,N_14900,N_14779);
nand UO_1955 (O_1955,N_14791,N_14950);
nand UO_1956 (O_1956,N_14756,N_14771);
or UO_1957 (O_1957,N_14842,N_14814);
nor UO_1958 (O_1958,N_14943,N_14854);
nor UO_1959 (O_1959,N_14913,N_14934);
nand UO_1960 (O_1960,N_14782,N_14966);
nor UO_1961 (O_1961,N_14976,N_14888);
or UO_1962 (O_1962,N_14751,N_14900);
and UO_1963 (O_1963,N_14935,N_14866);
nand UO_1964 (O_1964,N_14933,N_14767);
and UO_1965 (O_1965,N_14962,N_14892);
nor UO_1966 (O_1966,N_14763,N_14776);
nor UO_1967 (O_1967,N_14876,N_14808);
nor UO_1968 (O_1968,N_14801,N_14754);
and UO_1969 (O_1969,N_14818,N_14956);
nor UO_1970 (O_1970,N_14930,N_14856);
or UO_1971 (O_1971,N_14978,N_14899);
and UO_1972 (O_1972,N_14898,N_14769);
nor UO_1973 (O_1973,N_14907,N_14875);
or UO_1974 (O_1974,N_14975,N_14982);
and UO_1975 (O_1975,N_14998,N_14941);
nor UO_1976 (O_1976,N_14871,N_14859);
and UO_1977 (O_1977,N_14793,N_14833);
xor UO_1978 (O_1978,N_14772,N_14970);
and UO_1979 (O_1979,N_14824,N_14780);
or UO_1980 (O_1980,N_14859,N_14823);
and UO_1981 (O_1981,N_14811,N_14780);
or UO_1982 (O_1982,N_14870,N_14916);
or UO_1983 (O_1983,N_14950,N_14824);
nand UO_1984 (O_1984,N_14969,N_14993);
nand UO_1985 (O_1985,N_14833,N_14823);
nor UO_1986 (O_1986,N_14855,N_14824);
nor UO_1987 (O_1987,N_14948,N_14979);
nor UO_1988 (O_1988,N_14980,N_14812);
and UO_1989 (O_1989,N_14995,N_14945);
xor UO_1990 (O_1990,N_14920,N_14841);
or UO_1991 (O_1991,N_14989,N_14758);
nor UO_1992 (O_1992,N_14798,N_14800);
or UO_1993 (O_1993,N_14929,N_14916);
nor UO_1994 (O_1994,N_14814,N_14990);
nor UO_1995 (O_1995,N_14953,N_14812);
nand UO_1996 (O_1996,N_14987,N_14991);
nor UO_1997 (O_1997,N_14905,N_14975);
and UO_1998 (O_1998,N_14849,N_14967);
nand UO_1999 (O_1999,N_14758,N_14845);
endmodule