module basic_1000_10000_1500_10_levels_2xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_483,In_410);
or U1 (N_1,In_575,In_317);
nand U2 (N_2,In_722,In_670);
nand U3 (N_3,In_791,In_466);
nand U4 (N_4,In_35,In_877);
nor U5 (N_5,In_43,In_332);
and U6 (N_6,In_739,In_621);
or U7 (N_7,In_93,In_197);
and U8 (N_8,In_29,In_540);
and U9 (N_9,In_781,In_685);
and U10 (N_10,In_924,In_452);
nor U11 (N_11,In_443,In_57);
nor U12 (N_12,In_464,In_942);
xnor U13 (N_13,In_899,In_480);
nor U14 (N_14,In_773,In_566);
and U15 (N_15,In_103,In_66);
or U16 (N_16,In_819,In_285);
nor U17 (N_17,In_850,In_714);
nand U18 (N_18,In_358,In_174);
nor U19 (N_19,In_952,In_854);
or U20 (N_20,In_698,In_210);
nand U21 (N_21,In_516,In_439);
and U22 (N_22,In_918,In_327);
or U23 (N_23,In_765,In_709);
and U24 (N_24,In_65,In_926);
nor U25 (N_25,In_239,In_852);
nor U26 (N_26,In_553,In_651);
nor U27 (N_27,In_624,In_376);
nor U28 (N_28,In_196,In_118);
nor U29 (N_29,In_761,In_719);
nand U30 (N_30,In_727,In_237);
or U31 (N_31,In_231,In_969);
nor U32 (N_32,In_808,In_705);
nor U33 (N_33,In_862,In_973);
and U34 (N_34,In_726,In_129);
nand U35 (N_35,In_929,In_559);
or U36 (N_36,In_92,In_989);
or U37 (N_37,In_731,In_342);
nor U38 (N_38,In_999,In_419);
nand U39 (N_39,In_244,In_33);
and U40 (N_40,In_113,In_763);
and U41 (N_41,In_785,In_992);
and U42 (N_42,In_655,In_644);
nor U43 (N_43,In_914,In_672);
nor U44 (N_44,In_707,In_178);
nand U45 (N_45,In_526,In_472);
or U46 (N_46,In_179,In_135);
and U47 (N_47,In_76,In_95);
xor U48 (N_48,In_863,In_512);
nor U49 (N_49,In_905,In_499);
and U50 (N_50,In_202,In_673);
xnor U51 (N_51,In_520,In_701);
nand U52 (N_52,In_167,In_356);
and U53 (N_53,In_31,In_414);
xor U54 (N_54,In_552,In_52);
nand U55 (N_55,In_617,In_416);
nor U56 (N_56,In_787,In_832);
nor U57 (N_57,In_334,In_886);
nand U58 (N_58,In_923,In_176);
and U59 (N_59,In_408,In_485);
nor U60 (N_60,In_858,In_501);
nand U61 (N_61,In_505,In_157);
or U62 (N_62,In_15,In_804);
nand U63 (N_63,In_625,In_823);
and U64 (N_64,In_551,In_68);
nor U65 (N_65,In_126,In_421);
nor U66 (N_66,In_311,In_557);
or U67 (N_67,In_451,In_534);
or U68 (N_68,In_8,In_982);
or U69 (N_69,In_919,In_561);
or U70 (N_70,In_404,In_475);
xnor U71 (N_71,In_912,In_943);
and U72 (N_72,In_909,In_184);
nand U73 (N_73,In_836,In_381);
or U74 (N_74,In_164,In_54);
nor U75 (N_75,In_870,In_693);
and U76 (N_76,In_903,In_881);
nor U77 (N_77,In_588,In_90);
nand U78 (N_78,In_322,In_663);
or U79 (N_79,In_712,In_435);
or U80 (N_80,In_73,In_345);
nand U81 (N_81,In_977,In_742);
nor U82 (N_82,In_793,In_240);
or U83 (N_83,In_812,In_704);
nand U84 (N_84,In_266,In_611);
nand U85 (N_85,In_309,In_971);
or U86 (N_86,In_0,In_851);
xnor U87 (N_87,In_411,In_252);
nor U88 (N_88,In_567,In_777);
nor U89 (N_89,In_541,In_107);
nor U90 (N_90,In_831,In_106);
nor U91 (N_91,In_981,In_97);
nor U92 (N_92,In_955,In_128);
and U93 (N_93,In_716,In_199);
and U94 (N_94,In_333,In_98);
nor U95 (N_95,In_945,In_359);
and U96 (N_96,In_58,In_121);
or U97 (N_97,In_876,In_161);
and U98 (N_98,In_491,In_323);
nor U99 (N_99,In_647,In_799);
or U100 (N_100,In_1,In_703);
nor U101 (N_101,In_904,In_610);
or U102 (N_102,In_995,In_980);
nor U103 (N_103,In_151,In_99);
nand U104 (N_104,In_769,In_771);
nand U105 (N_105,In_548,In_104);
or U106 (N_106,In_163,In_294);
or U107 (N_107,In_778,In_286);
and U108 (N_108,In_415,In_717);
nand U109 (N_109,In_222,In_966);
nand U110 (N_110,In_79,In_521);
nand U111 (N_111,In_535,In_3);
or U112 (N_112,In_509,In_738);
nor U113 (N_113,In_585,In_983);
nor U114 (N_114,In_312,In_185);
xor U115 (N_115,In_604,In_127);
nor U116 (N_116,In_361,In_502);
nor U117 (N_117,In_384,In_511);
and U118 (N_118,In_896,In_759);
nand U119 (N_119,In_490,In_20);
nand U120 (N_120,In_331,In_387);
or U121 (N_121,In_389,In_214);
nand U122 (N_122,In_676,In_120);
or U123 (N_123,In_867,In_786);
nor U124 (N_124,In_233,In_28);
nor U125 (N_125,In_613,In_578);
and U126 (N_126,In_513,In_690);
nand U127 (N_127,In_965,In_142);
nor U128 (N_128,In_232,In_123);
nor U129 (N_129,In_438,In_460);
and U130 (N_130,In_463,In_906);
nand U131 (N_131,In_378,In_735);
and U132 (N_132,In_382,In_148);
nor U133 (N_133,In_353,In_348);
or U134 (N_134,In_82,In_399);
nand U135 (N_135,In_730,In_375);
xor U136 (N_136,In_394,In_476);
or U137 (N_137,In_132,In_874);
or U138 (N_138,In_547,In_207);
nand U139 (N_139,In_577,In_56);
or U140 (N_140,In_556,In_951);
nand U141 (N_141,In_679,In_713);
or U142 (N_142,In_170,In_440);
and U143 (N_143,In_927,In_803);
nand U144 (N_144,In_349,In_287);
nor U145 (N_145,In_650,In_189);
nand U146 (N_146,In_397,In_635);
or U147 (N_147,In_290,In_236);
nand U148 (N_148,In_269,In_109);
and U149 (N_149,In_291,In_783);
and U150 (N_150,In_879,In_426);
nor U151 (N_151,In_263,In_453);
xor U152 (N_152,In_70,In_883);
and U153 (N_153,In_94,In_921);
nor U154 (N_154,In_117,In_367);
and U155 (N_155,In_871,In_657);
nor U156 (N_156,In_855,In_221);
or U157 (N_157,In_620,In_193);
and U158 (N_158,In_506,In_50);
and U159 (N_159,In_619,In_841);
nor U160 (N_160,In_493,In_39);
nand U161 (N_161,In_162,In_865);
nor U162 (N_162,In_976,In_171);
nand U163 (N_163,In_319,In_542);
nand U164 (N_164,In_366,In_779);
nor U165 (N_165,In_935,In_797);
or U166 (N_166,In_328,In_733);
nand U167 (N_167,In_915,In_796);
or U168 (N_168,In_868,In_86);
xor U169 (N_169,In_860,In_259);
nor U170 (N_170,In_44,In_743);
and U171 (N_171,In_531,In_201);
and U172 (N_172,In_504,In_271);
and U173 (N_173,In_589,In_36);
and U174 (N_174,In_816,In_26);
or U175 (N_175,In_514,In_861);
nor U176 (N_176,In_10,In_363);
xnor U177 (N_177,In_159,In_139);
or U178 (N_178,In_622,In_338);
and U179 (N_179,In_274,In_975);
nand U180 (N_180,In_265,In_165);
nand U181 (N_181,In_42,In_62);
and U182 (N_182,In_710,In_145);
and U183 (N_183,In_450,In_418);
nand U184 (N_184,In_427,In_393);
nand U185 (N_185,In_790,In_27);
nor U186 (N_186,In_887,In_194);
nor U187 (N_187,In_153,In_489);
nor U188 (N_188,In_864,In_218);
or U189 (N_189,In_643,In_347);
nand U190 (N_190,In_425,In_337);
or U191 (N_191,In_19,In_664);
or U192 (N_192,In_192,In_306);
and U193 (N_193,In_674,In_217);
or U194 (N_194,In_5,In_702);
or U195 (N_195,In_325,In_902);
nand U196 (N_196,In_937,In_661);
nand U197 (N_197,In_750,In_970);
nand U198 (N_198,In_143,In_571);
and U199 (N_199,In_229,In_91);
nor U200 (N_200,In_302,In_696);
or U201 (N_201,In_433,In_293);
or U202 (N_202,In_9,In_351);
and U203 (N_203,In_364,In_754);
nand U204 (N_204,In_96,In_102);
or U205 (N_205,In_253,In_38);
and U206 (N_206,In_947,In_968);
or U207 (N_207,In_209,In_608);
nor U208 (N_208,In_155,In_30);
xor U209 (N_209,In_596,In_396);
and U210 (N_210,In_205,In_242);
or U211 (N_211,In_63,In_821);
and U212 (N_212,In_314,In_597);
or U213 (N_213,In_187,In_431);
or U214 (N_214,In_724,In_67);
or U215 (N_215,In_454,In_447);
nor U216 (N_216,In_402,In_296);
or U217 (N_217,In_634,In_303);
and U218 (N_218,In_517,In_448);
or U219 (N_219,In_130,In_468);
nor U220 (N_220,In_262,In_388);
nand U221 (N_221,In_304,In_49);
and U222 (N_222,In_108,In_14);
nor U223 (N_223,In_340,In_297);
and U224 (N_224,In_115,In_191);
nand U225 (N_225,In_747,In_160);
or U226 (N_226,In_72,In_316);
nand U227 (N_227,In_321,In_758);
and U228 (N_228,In_849,In_522);
and U229 (N_229,In_536,In_254);
nor U230 (N_230,In_795,In_188);
or U231 (N_231,In_668,In_789);
and U232 (N_232,In_152,In_149);
nand U233 (N_233,In_748,In_979);
and U234 (N_234,In_400,In_329);
or U235 (N_235,In_554,In_219);
and U236 (N_236,In_658,In_628);
and U237 (N_237,In_728,In_930);
nand U238 (N_238,In_800,In_500);
xnor U239 (N_239,In_69,In_273);
or U240 (N_240,In_458,In_6);
nor U241 (N_241,In_687,In_767);
or U242 (N_242,In_944,In_241);
nor U243 (N_243,In_295,In_374);
nand U244 (N_244,In_948,In_277);
and U245 (N_245,In_462,In_568);
nand U246 (N_246,In_246,In_788);
nor U247 (N_247,In_250,In_605);
and U248 (N_248,In_495,In_371);
nand U249 (N_249,In_580,In_124);
and U250 (N_250,In_873,In_671);
xor U251 (N_251,In_916,In_830);
xor U252 (N_252,In_428,In_933);
nand U253 (N_253,In_558,In_465);
nand U254 (N_254,In_649,In_17);
nor U255 (N_255,In_344,In_180);
or U256 (N_256,In_318,In_835);
xnor U257 (N_257,In_928,In_570);
xnor U258 (N_258,In_343,In_996);
nor U259 (N_259,In_662,In_890);
or U260 (N_260,In_776,In_715);
nand U261 (N_261,In_372,In_430);
and U262 (N_262,In_562,In_477);
nor U263 (N_263,In_467,In_582);
or U264 (N_264,In_642,In_938);
nand U265 (N_265,In_482,In_801);
nand U266 (N_266,In_114,In_473);
and U267 (N_267,In_195,In_105);
and U268 (N_268,In_544,In_45);
and U269 (N_269,In_292,In_931);
nor U270 (N_270,In_936,In_456);
nand U271 (N_271,In_412,In_324);
nand U272 (N_272,In_227,In_564);
or U273 (N_273,In_498,In_950);
or U274 (N_274,In_607,In_299);
nand U275 (N_275,In_137,In_760);
or U276 (N_276,In_820,In_474);
nand U277 (N_277,In_959,In_249);
nor U278 (N_278,In_882,In_892);
or U279 (N_279,In_827,In_407);
and U280 (N_280,In_639,In_768);
or U281 (N_281,In_510,In_654);
or U282 (N_282,In_432,In_225);
nand U283 (N_283,In_395,In_424);
nand U284 (N_284,In_811,In_998);
nand U285 (N_285,In_563,In_326);
or U286 (N_286,In_87,In_711);
and U287 (N_287,In_12,In_962);
and U288 (N_288,In_618,In_75);
nand U289 (N_289,In_680,In_683);
and U290 (N_290,In_708,In_984);
and U291 (N_291,In_48,In_838);
nor U292 (N_292,In_298,In_720);
nor U293 (N_293,In_626,In_636);
and U294 (N_294,In_543,In_166);
and U295 (N_295,In_383,In_910);
nor U296 (N_296,In_565,In_974);
or U297 (N_297,In_721,In_601);
or U298 (N_298,In_507,In_243);
and U299 (N_299,In_857,In_891);
or U300 (N_300,In_208,In_352);
nand U301 (N_301,In_737,In_700);
and U302 (N_302,In_251,In_261);
or U303 (N_303,In_745,In_818);
nor U304 (N_304,In_486,In_84);
or U305 (N_305,In_18,In_590);
or U306 (N_306,In_181,In_665);
nor U307 (N_307,In_508,In_775);
or U308 (N_308,In_834,In_469);
nor U309 (N_309,In_546,In_689);
and U310 (N_310,In_158,In_678);
nor U311 (N_311,In_774,In_81);
and U312 (N_312,In_436,In_925);
nor U313 (N_313,In_591,In_606);
nand U314 (N_314,In_963,In_23);
nor U315 (N_315,In_560,In_40);
and U316 (N_316,In_341,In_77);
and U317 (N_317,In_784,In_320);
nand U318 (N_318,In_630,In_16);
and U319 (N_319,In_527,In_885);
or U320 (N_320,In_813,In_487);
nor U321 (N_321,In_484,In_756);
and U322 (N_322,In_686,In_446);
or U323 (N_323,In_814,In_136);
nor U324 (N_324,In_330,In_119);
nand U325 (N_325,In_220,In_986);
and U326 (N_326,In_741,In_183);
nand U327 (N_327,In_146,In_616);
nor U328 (N_328,In_275,In_991);
nor U329 (N_329,In_572,In_940);
nand U330 (N_330,In_762,In_972);
nand U331 (N_331,In_200,In_782);
nor U332 (N_332,In_752,In_78);
and U333 (N_333,In_666,In_496);
and U334 (N_334,In_894,In_357);
nor U335 (N_335,In_32,In_772);
nand U336 (N_336,In_22,In_350);
xor U337 (N_337,In_523,In_260);
nand U338 (N_338,In_4,In_279);
nand U339 (N_339,In_525,In_893);
or U340 (N_340,In_853,In_583);
and U341 (N_341,In_900,In_405);
nand U342 (N_342,In_398,In_681);
nand U343 (N_343,In_422,In_211);
and U344 (N_344,In_956,In_539);
nor U345 (N_345,In_631,In_815);
and U346 (N_346,In_7,In_718);
nor U347 (N_347,In_660,In_494);
nor U348 (N_348,In_629,In_386);
nand U349 (N_349,In_602,In_889);
or U350 (N_350,In_528,In_549);
nor U351 (N_351,In_614,In_985);
nand U352 (N_352,In_257,In_60);
or U353 (N_353,In_826,In_839);
and U354 (N_354,In_844,In_593);
and U355 (N_355,In_958,In_335);
and U356 (N_356,In_798,In_845);
and U357 (N_357,In_100,In_574);
or U358 (N_358,In_88,In_988);
or U359 (N_359,In_391,In_751);
nor U360 (N_360,In_216,In_584);
nor U361 (N_361,In_946,In_503);
nor U362 (N_362,In_792,In_122);
nor U363 (N_363,In_833,In_888);
nand U364 (N_364,In_434,In_939);
or U365 (N_365,In_212,In_51);
and U366 (N_366,In_169,In_470);
or U367 (N_367,In_282,In_336);
nor U368 (N_368,In_805,In_2);
nor U369 (N_369,In_133,In_360);
nor U370 (N_370,In_638,In_268);
or U371 (N_371,In_697,In_579);
nor U372 (N_372,In_213,In_21);
or U373 (N_373,In_669,In_71);
or U374 (N_374,In_368,In_652);
and U375 (N_375,In_417,In_729);
and U376 (N_376,In_288,In_744);
and U377 (N_377,In_101,In_215);
nand U378 (N_378,In_645,In_569);
nor U379 (N_379,In_550,In_110);
or U380 (N_380,In_85,In_755);
or U381 (N_381,In_623,In_581);
nor U382 (N_382,In_444,In_455);
nor U383 (N_383,In_147,In_369);
and U384 (N_384,In_390,In_706);
xor U385 (N_385,In_964,In_961);
or U386 (N_386,In_954,In_355);
and U387 (N_387,In_272,In_633);
or U388 (N_388,In_587,In_173);
nor U389 (N_389,In_300,In_770);
xnor U390 (N_390,In_198,In_609);
or U391 (N_391,In_573,In_406);
nor U392 (N_392,In_866,In_445);
and U393 (N_393,In_492,In_449);
nor U394 (N_394,In_824,In_112);
nor U395 (N_395,In_545,In_278);
nor U396 (N_396,In_646,In_289);
or U397 (N_397,In_682,In_156);
or U398 (N_398,In_880,In_640);
or U399 (N_399,In_691,In_807);
nand U400 (N_400,In_822,In_809);
xnor U401 (N_401,In_828,In_190);
nand U402 (N_402,In_154,In_598);
nand U403 (N_403,In_627,In_37);
nor U404 (N_404,In_695,In_204);
nor U405 (N_405,In_226,In_684);
nand U406 (N_406,In_967,In_248);
or U407 (N_407,In_481,In_413);
nor U408 (N_408,In_442,In_41);
nand U409 (N_409,In_732,In_429);
and U410 (N_410,In_595,In_911);
nor U411 (N_411,In_632,In_960);
and U412 (N_412,In_441,In_667);
nand U413 (N_413,In_603,In_125);
nand U414 (N_414,In_224,In_766);
nor U415 (N_415,In_258,In_284);
nor U416 (N_416,In_47,In_978);
nand U417 (N_417,In_884,In_901);
or U418 (N_418,In_538,In_459);
or U419 (N_419,In_941,In_403);
and U420 (N_420,In_53,In_537);
nor U421 (N_421,In_897,In_310);
and U422 (N_422,In_281,In_401);
and U423 (N_423,In_872,In_895);
or U424 (N_424,In_920,In_692);
and U425 (N_425,In_177,In_409);
nor U426 (N_426,In_878,In_725);
nor U427 (N_427,In_847,In_576);
or U428 (N_428,In_599,In_111);
and U429 (N_429,In_354,In_780);
or U430 (N_430,In_307,In_373);
nor U431 (N_431,In_917,In_255);
nor U432 (N_432,In_80,In_806);
nor U433 (N_433,In_256,In_757);
or U434 (N_434,In_234,In_235);
nand U435 (N_435,In_457,In_346);
nand U436 (N_436,In_83,In_471);
nor U437 (N_437,In_533,In_339);
and U438 (N_438,In_829,In_817);
nand U439 (N_439,In_203,In_934);
or U440 (N_440,In_61,In_313);
or U441 (N_441,In_524,In_515);
nor U442 (N_442,In_753,In_437);
and U443 (N_443,In_461,In_846);
nand U444 (N_444,In_140,In_270);
or U445 (N_445,In_25,In_997);
and U446 (N_446,In_842,In_186);
nor U447 (N_447,In_138,In_11);
nand U448 (N_448,In_848,In_423);
nor U449 (N_449,In_478,In_34);
nor U450 (N_450,In_380,In_764);
or U451 (N_451,In_907,In_46);
nor U452 (N_452,In_856,In_932);
nor U453 (N_453,In_24,In_530);
nand U454 (N_454,In_385,In_875);
nor U455 (N_455,In_116,In_74);
and U456 (N_456,In_675,In_908);
and U457 (N_457,In_144,In_228);
and U458 (N_458,In_555,In_301);
nor U459 (N_459,In_168,In_736);
nor U460 (N_460,In_734,In_648);
and U461 (N_461,In_922,In_869);
nor U462 (N_462,In_659,In_594);
or U463 (N_463,In_280,In_370);
and U464 (N_464,In_479,In_637);
or U465 (N_465,In_247,In_55);
and U466 (N_466,In_740,In_794);
or U467 (N_467,In_131,In_843);
nand U468 (N_468,In_586,In_245);
nand U469 (N_469,In_957,In_532);
or U470 (N_470,In_182,In_840);
and U471 (N_471,In_592,In_172);
nor U472 (N_472,In_749,In_723);
or U473 (N_473,In_134,In_994);
and U474 (N_474,In_308,In_315);
or U475 (N_475,In_283,In_699);
nor U476 (N_476,In_267,In_13);
and U477 (N_477,In_825,In_898);
nor U478 (N_478,In_653,In_953);
nand U479 (N_479,In_238,In_420);
nor U480 (N_480,In_59,In_175);
nand U481 (N_481,In_206,In_488);
or U482 (N_482,In_230,In_615);
and U483 (N_483,In_519,In_392);
nand U484 (N_484,In_677,In_859);
or U485 (N_485,In_612,In_949);
or U486 (N_486,In_802,In_600);
nand U487 (N_487,In_656,In_223);
and U488 (N_488,In_837,In_362);
or U489 (N_489,In_688,In_150);
or U490 (N_490,In_365,In_89);
and U491 (N_491,In_379,In_810);
or U492 (N_492,In_993,In_746);
nand U493 (N_493,In_913,In_529);
and U494 (N_494,In_987,In_641);
xnor U495 (N_495,In_305,In_990);
or U496 (N_496,In_64,In_276);
and U497 (N_497,In_377,In_497);
and U498 (N_498,In_518,In_141);
or U499 (N_499,In_694,In_264);
nor U500 (N_500,In_545,In_99);
and U501 (N_501,In_860,In_50);
nand U502 (N_502,In_21,In_666);
or U503 (N_503,In_415,In_509);
and U504 (N_504,In_367,In_655);
or U505 (N_505,In_312,In_146);
nor U506 (N_506,In_761,In_342);
xor U507 (N_507,In_210,In_609);
or U508 (N_508,In_67,In_945);
and U509 (N_509,In_9,In_122);
nand U510 (N_510,In_844,In_530);
nor U511 (N_511,In_183,In_711);
nand U512 (N_512,In_820,In_193);
nor U513 (N_513,In_994,In_110);
nor U514 (N_514,In_68,In_111);
nand U515 (N_515,In_423,In_416);
nor U516 (N_516,In_907,In_806);
and U517 (N_517,In_141,In_657);
nand U518 (N_518,In_487,In_810);
and U519 (N_519,In_889,In_688);
or U520 (N_520,In_405,In_542);
or U521 (N_521,In_828,In_602);
and U522 (N_522,In_618,In_175);
or U523 (N_523,In_107,In_715);
and U524 (N_524,In_619,In_200);
nand U525 (N_525,In_735,In_655);
nor U526 (N_526,In_942,In_988);
nor U527 (N_527,In_95,In_55);
nor U528 (N_528,In_546,In_782);
nand U529 (N_529,In_838,In_221);
xnor U530 (N_530,In_109,In_564);
or U531 (N_531,In_496,In_315);
or U532 (N_532,In_26,In_86);
nor U533 (N_533,In_448,In_350);
nand U534 (N_534,In_201,In_88);
nor U535 (N_535,In_134,In_537);
and U536 (N_536,In_772,In_118);
or U537 (N_537,In_747,In_955);
or U538 (N_538,In_171,In_375);
xnor U539 (N_539,In_160,In_295);
nor U540 (N_540,In_366,In_360);
and U541 (N_541,In_104,In_495);
nor U542 (N_542,In_510,In_5);
and U543 (N_543,In_25,In_567);
or U544 (N_544,In_535,In_854);
nor U545 (N_545,In_654,In_449);
and U546 (N_546,In_670,In_897);
nand U547 (N_547,In_897,In_110);
nand U548 (N_548,In_508,In_366);
nand U549 (N_549,In_132,In_806);
nor U550 (N_550,In_891,In_917);
and U551 (N_551,In_235,In_818);
or U552 (N_552,In_706,In_468);
nand U553 (N_553,In_130,In_870);
and U554 (N_554,In_461,In_966);
or U555 (N_555,In_414,In_685);
nor U556 (N_556,In_420,In_535);
and U557 (N_557,In_904,In_45);
nor U558 (N_558,In_232,In_550);
or U559 (N_559,In_890,In_190);
and U560 (N_560,In_547,In_942);
nor U561 (N_561,In_998,In_542);
nand U562 (N_562,In_270,In_77);
nor U563 (N_563,In_862,In_889);
or U564 (N_564,In_111,In_967);
and U565 (N_565,In_624,In_403);
or U566 (N_566,In_716,In_102);
nand U567 (N_567,In_254,In_493);
and U568 (N_568,In_372,In_385);
nor U569 (N_569,In_344,In_263);
xor U570 (N_570,In_681,In_483);
nand U571 (N_571,In_773,In_851);
or U572 (N_572,In_511,In_562);
nor U573 (N_573,In_213,In_695);
nand U574 (N_574,In_219,In_703);
nand U575 (N_575,In_864,In_990);
nor U576 (N_576,In_895,In_788);
xnor U577 (N_577,In_637,In_95);
nor U578 (N_578,In_180,In_113);
nor U579 (N_579,In_273,In_821);
nand U580 (N_580,In_55,In_204);
nor U581 (N_581,In_41,In_781);
and U582 (N_582,In_729,In_258);
nor U583 (N_583,In_469,In_288);
xor U584 (N_584,In_683,In_766);
nor U585 (N_585,In_939,In_249);
or U586 (N_586,In_871,In_415);
and U587 (N_587,In_804,In_814);
or U588 (N_588,In_696,In_866);
nand U589 (N_589,In_411,In_688);
and U590 (N_590,In_920,In_203);
or U591 (N_591,In_662,In_823);
and U592 (N_592,In_359,In_416);
or U593 (N_593,In_211,In_312);
xor U594 (N_594,In_105,In_638);
nor U595 (N_595,In_521,In_871);
xor U596 (N_596,In_922,In_321);
or U597 (N_597,In_693,In_215);
nor U598 (N_598,In_330,In_905);
or U599 (N_599,In_947,In_932);
nand U600 (N_600,In_761,In_247);
or U601 (N_601,In_57,In_132);
and U602 (N_602,In_397,In_818);
and U603 (N_603,In_356,In_99);
and U604 (N_604,In_875,In_228);
or U605 (N_605,In_264,In_688);
and U606 (N_606,In_566,In_258);
nand U607 (N_607,In_466,In_456);
and U608 (N_608,In_35,In_933);
nor U609 (N_609,In_443,In_107);
nor U610 (N_610,In_407,In_60);
xnor U611 (N_611,In_586,In_880);
and U612 (N_612,In_222,In_941);
xor U613 (N_613,In_379,In_386);
nand U614 (N_614,In_875,In_709);
or U615 (N_615,In_548,In_773);
nor U616 (N_616,In_383,In_36);
or U617 (N_617,In_579,In_901);
or U618 (N_618,In_727,In_593);
nand U619 (N_619,In_93,In_325);
nand U620 (N_620,In_395,In_368);
nor U621 (N_621,In_448,In_913);
nand U622 (N_622,In_913,In_711);
nor U623 (N_623,In_597,In_140);
nand U624 (N_624,In_449,In_770);
or U625 (N_625,In_93,In_342);
nor U626 (N_626,In_108,In_427);
or U627 (N_627,In_42,In_335);
or U628 (N_628,In_248,In_540);
nand U629 (N_629,In_140,In_29);
nor U630 (N_630,In_41,In_17);
and U631 (N_631,In_67,In_198);
or U632 (N_632,In_652,In_809);
nor U633 (N_633,In_617,In_836);
nand U634 (N_634,In_848,In_296);
nand U635 (N_635,In_183,In_854);
or U636 (N_636,In_310,In_340);
and U637 (N_637,In_727,In_112);
nor U638 (N_638,In_521,In_643);
nand U639 (N_639,In_29,In_450);
and U640 (N_640,In_254,In_260);
nand U641 (N_641,In_629,In_42);
nand U642 (N_642,In_410,In_587);
nand U643 (N_643,In_132,In_982);
or U644 (N_644,In_630,In_933);
nor U645 (N_645,In_641,In_250);
nor U646 (N_646,In_306,In_438);
and U647 (N_647,In_163,In_884);
and U648 (N_648,In_192,In_705);
nand U649 (N_649,In_164,In_432);
nor U650 (N_650,In_316,In_127);
and U651 (N_651,In_953,In_229);
nor U652 (N_652,In_424,In_810);
nor U653 (N_653,In_164,In_564);
nand U654 (N_654,In_357,In_817);
nor U655 (N_655,In_557,In_564);
nand U656 (N_656,In_554,In_431);
nand U657 (N_657,In_615,In_109);
and U658 (N_658,In_352,In_639);
or U659 (N_659,In_728,In_666);
nand U660 (N_660,In_974,In_238);
and U661 (N_661,In_696,In_221);
and U662 (N_662,In_764,In_391);
and U663 (N_663,In_80,In_348);
nand U664 (N_664,In_830,In_586);
and U665 (N_665,In_902,In_335);
nand U666 (N_666,In_461,In_742);
nor U667 (N_667,In_754,In_367);
nor U668 (N_668,In_624,In_785);
or U669 (N_669,In_285,In_317);
or U670 (N_670,In_174,In_415);
or U671 (N_671,In_929,In_475);
and U672 (N_672,In_940,In_173);
nor U673 (N_673,In_644,In_845);
and U674 (N_674,In_432,In_220);
nor U675 (N_675,In_515,In_325);
or U676 (N_676,In_944,In_740);
nor U677 (N_677,In_679,In_589);
nand U678 (N_678,In_579,In_689);
nor U679 (N_679,In_35,In_323);
and U680 (N_680,In_80,In_231);
and U681 (N_681,In_553,In_808);
nand U682 (N_682,In_698,In_793);
and U683 (N_683,In_993,In_714);
and U684 (N_684,In_649,In_561);
nand U685 (N_685,In_490,In_952);
or U686 (N_686,In_225,In_947);
nor U687 (N_687,In_647,In_346);
or U688 (N_688,In_756,In_843);
nor U689 (N_689,In_636,In_63);
or U690 (N_690,In_894,In_724);
and U691 (N_691,In_345,In_592);
nor U692 (N_692,In_233,In_468);
nor U693 (N_693,In_726,In_710);
or U694 (N_694,In_327,In_329);
nand U695 (N_695,In_943,In_48);
and U696 (N_696,In_171,In_350);
xor U697 (N_697,In_751,In_82);
or U698 (N_698,In_343,In_228);
nand U699 (N_699,In_497,In_679);
nand U700 (N_700,In_520,In_900);
or U701 (N_701,In_544,In_495);
or U702 (N_702,In_712,In_729);
or U703 (N_703,In_466,In_666);
nand U704 (N_704,In_649,In_333);
nand U705 (N_705,In_337,In_472);
or U706 (N_706,In_826,In_555);
or U707 (N_707,In_221,In_743);
or U708 (N_708,In_696,In_322);
nand U709 (N_709,In_38,In_161);
nand U710 (N_710,In_349,In_725);
nor U711 (N_711,In_465,In_786);
or U712 (N_712,In_24,In_814);
and U713 (N_713,In_108,In_814);
or U714 (N_714,In_298,In_421);
nor U715 (N_715,In_596,In_857);
xnor U716 (N_716,In_663,In_176);
nor U717 (N_717,In_556,In_625);
nor U718 (N_718,In_500,In_358);
nor U719 (N_719,In_727,In_944);
or U720 (N_720,In_613,In_263);
nor U721 (N_721,In_808,In_143);
or U722 (N_722,In_826,In_135);
nor U723 (N_723,In_211,In_343);
xnor U724 (N_724,In_14,In_11);
and U725 (N_725,In_927,In_125);
xnor U726 (N_726,In_378,In_486);
and U727 (N_727,In_345,In_308);
nand U728 (N_728,In_776,In_838);
nand U729 (N_729,In_228,In_150);
and U730 (N_730,In_554,In_283);
nand U731 (N_731,In_136,In_293);
and U732 (N_732,In_78,In_413);
and U733 (N_733,In_571,In_35);
or U734 (N_734,In_402,In_945);
nor U735 (N_735,In_361,In_495);
nor U736 (N_736,In_748,In_936);
nor U737 (N_737,In_248,In_919);
and U738 (N_738,In_488,In_754);
nand U739 (N_739,In_347,In_814);
and U740 (N_740,In_656,In_854);
nand U741 (N_741,In_425,In_818);
nor U742 (N_742,In_788,In_775);
nand U743 (N_743,In_500,In_245);
nand U744 (N_744,In_209,In_858);
nor U745 (N_745,In_713,In_979);
and U746 (N_746,In_422,In_296);
or U747 (N_747,In_907,In_604);
and U748 (N_748,In_104,In_118);
nand U749 (N_749,In_334,In_960);
nand U750 (N_750,In_63,In_161);
nand U751 (N_751,In_872,In_248);
and U752 (N_752,In_160,In_677);
nor U753 (N_753,In_458,In_201);
nand U754 (N_754,In_555,In_90);
or U755 (N_755,In_587,In_852);
and U756 (N_756,In_566,In_867);
and U757 (N_757,In_378,In_641);
and U758 (N_758,In_213,In_229);
or U759 (N_759,In_417,In_288);
nand U760 (N_760,In_939,In_536);
or U761 (N_761,In_50,In_664);
and U762 (N_762,In_281,In_869);
nand U763 (N_763,In_675,In_47);
or U764 (N_764,In_549,In_24);
or U765 (N_765,In_690,In_911);
or U766 (N_766,In_271,In_846);
and U767 (N_767,In_953,In_54);
nand U768 (N_768,In_23,In_899);
xor U769 (N_769,In_48,In_78);
nor U770 (N_770,In_62,In_401);
nand U771 (N_771,In_472,In_487);
nor U772 (N_772,In_691,In_929);
nand U773 (N_773,In_281,In_297);
nor U774 (N_774,In_960,In_397);
or U775 (N_775,In_727,In_826);
nor U776 (N_776,In_611,In_695);
or U777 (N_777,In_699,In_720);
and U778 (N_778,In_916,In_657);
or U779 (N_779,In_852,In_161);
and U780 (N_780,In_666,In_754);
nand U781 (N_781,In_442,In_173);
xor U782 (N_782,In_915,In_995);
and U783 (N_783,In_598,In_325);
or U784 (N_784,In_1,In_163);
nand U785 (N_785,In_334,In_259);
or U786 (N_786,In_108,In_815);
and U787 (N_787,In_709,In_253);
and U788 (N_788,In_161,In_3);
nor U789 (N_789,In_393,In_859);
nand U790 (N_790,In_50,In_159);
or U791 (N_791,In_290,In_916);
and U792 (N_792,In_891,In_204);
or U793 (N_793,In_856,In_890);
nand U794 (N_794,In_461,In_985);
nand U795 (N_795,In_961,In_975);
or U796 (N_796,In_739,In_784);
and U797 (N_797,In_656,In_792);
and U798 (N_798,In_211,In_872);
nand U799 (N_799,In_182,In_573);
nor U800 (N_800,In_80,In_432);
nand U801 (N_801,In_961,In_275);
and U802 (N_802,In_931,In_281);
or U803 (N_803,In_819,In_755);
and U804 (N_804,In_908,In_218);
nand U805 (N_805,In_516,In_673);
nor U806 (N_806,In_0,In_609);
and U807 (N_807,In_356,In_406);
xnor U808 (N_808,In_766,In_888);
nor U809 (N_809,In_473,In_464);
and U810 (N_810,In_208,In_801);
xor U811 (N_811,In_1,In_342);
nor U812 (N_812,In_555,In_102);
xor U813 (N_813,In_366,In_988);
nor U814 (N_814,In_392,In_855);
or U815 (N_815,In_81,In_168);
and U816 (N_816,In_761,In_34);
nor U817 (N_817,In_250,In_380);
nor U818 (N_818,In_191,In_274);
xnor U819 (N_819,In_210,In_190);
nor U820 (N_820,In_445,In_208);
nand U821 (N_821,In_752,In_459);
and U822 (N_822,In_694,In_665);
nand U823 (N_823,In_596,In_704);
and U824 (N_824,In_232,In_675);
nand U825 (N_825,In_132,In_755);
nand U826 (N_826,In_708,In_785);
nor U827 (N_827,In_500,In_40);
or U828 (N_828,In_749,In_816);
nor U829 (N_829,In_552,In_398);
or U830 (N_830,In_459,In_235);
nor U831 (N_831,In_647,In_123);
nor U832 (N_832,In_402,In_143);
or U833 (N_833,In_763,In_807);
nand U834 (N_834,In_395,In_694);
nor U835 (N_835,In_549,In_343);
or U836 (N_836,In_156,In_547);
or U837 (N_837,In_383,In_982);
nor U838 (N_838,In_821,In_250);
and U839 (N_839,In_354,In_875);
and U840 (N_840,In_546,In_443);
and U841 (N_841,In_768,In_724);
nand U842 (N_842,In_209,In_318);
nand U843 (N_843,In_50,In_147);
and U844 (N_844,In_628,In_676);
nand U845 (N_845,In_267,In_671);
or U846 (N_846,In_729,In_648);
nand U847 (N_847,In_497,In_966);
or U848 (N_848,In_394,In_781);
or U849 (N_849,In_778,In_937);
nor U850 (N_850,In_274,In_979);
nand U851 (N_851,In_26,In_253);
or U852 (N_852,In_973,In_237);
nand U853 (N_853,In_84,In_53);
or U854 (N_854,In_507,In_661);
nand U855 (N_855,In_507,In_948);
and U856 (N_856,In_409,In_297);
nand U857 (N_857,In_238,In_44);
nand U858 (N_858,In_26,In_656);
or U859 (N_859,In_171,In_182);
and U860 (N_860,In_919,In_247);
and U861 (N_861,In_240,In_242);
or U862 (N_862,In_349,In_983);
and U863 (N_863,In_12,In_438);
nor U864 (N_864,In_518,In_416);
nor U865 (N_865,In_531,In_576);
or U866 (N_866,In_386,In_188);
nand U867 (N_867,In_381,In_112);
nand U868 (N_868,In_283,In_64);
nand U869 (N_869,In_189,In_60);
xnor U870 (N_870,In_227,In_826);
nand U871 (N_871,In_130,In_229);
nand U872 (N_872,In_642,In_988);
nand U873 (N_873,In_968,In_267);
nand U874 (N_874,In_639,In_223);
nor U875 (N_875,In_359,In_529);
nand U876 (N_876,In_599,In_840);
or U877 (N_877,In_149,In_839);
nor U878 (N_878,In_233,In_363);
or U879 (N_879,In_390,In_974);
nor U880 (N_880,In_655,In_573);
nand U881 (N_881,In_223,In_502);
nand U882 (N_882,In_991,In_614);
xnor U883 (N_883,In_624,In_484);
nor U884 (N_884,In_657,In_921);
and U885 (N_885,In_524,In_135);
nand U886 (N_886,In_833,In_338);
nor U887 (N_887,In_797,In_695);
nor U888 (N_888,In_972,In_530);
nor U889 (N_889,In_104,In_587);
nor U890 (N_890,In_988,In_676);
nand U891 (N_891,In_696,In_72);
nor U892 (N_892,In_72,In_61);
nor U893 (N_893,In_248,In_857);
or U894 (N_894,In_388,In_140);
nor U895 (N_895,In_520,In_116);
nand U896 (N_896,In_618,In_39);
nor U897 (N_897,In_876,In_606);
or U898 (N_898,In_989,In_324);
and U899 (N_899,In_730,In_528);
nand U900 (N_900,In_192,In_529);
xor U901 (N_901,In_289,In_439);
nand U902 (N_902,In_235,In_150);
and U903 (N_903,In_372,In_327);
or U904 (N_904,In_393,In_661);
nand U905 (N_905,In_512,In_776);
nor U906 (N_906,In_101,In_957);
nor U907 (N_907,In_232,In_700);
or U908 (N_908,In_39,In_661);
or U909 (N_909,In_388,In_316);
and U910 (N_910,In_127,In_792);
nand U911 (N_911,In_642,In_987);
nand U912 (N_912,In_408,In_50);
nor U913 (N_913,In_794,In_487);
nor U914 (N_914,In_305,In_997);
nor U915 (N_915,In_310,In_288);
or U916 (N_916,In_389,In_196);
nand U917 (N_917,In_173,In_641);
nand U918 (N_918,In_587,In_131);
and U919 (N_919,In_842,In_650);
and U920 (N_920,In_305,In_917);
nor U921 (N_921,In_663,In_316);
or U922 (N_922,In_444,In_33);
nand U923 (N_923,In_495,In_565);
nand U924 (N_924,In_55,In_121);
and U925 (N_925,In_108,In_850);
nor U926 (N_926,In_593,In_125);
or U927 (N_927,In_168,In_126);
nand U928 (N_928,In_88,In_112);
nor U929 (N_929,In_780,In_52);
nor U930 (N_930,In_713,In_563);
nor U931 (N_931,In_964,In_785);
nor U932 (N_932,In_263,In_369);
and U933 (N_933,In_840,In_614);
nand U934 (N_934,In_441,In_889);
nor U935 (N_935,In_25,In_163);
nand U936 (N_936,In_128,In_374);
or U937 (N_937,In_640,In_183);
or U938 (N_938,In_171,In_668);
and U939 (N_939,In_514,In_320);
nor U940 (N_940,In_563,In_299);
nor U941 (N_941,In_25,In_821);
nor U942 (N_942,In_129,In_900);
and U943 (N_943,In_822,In_513);
or U944 (N_944,In_423,In_626);
nor U945 (N_945,In_272,In_647);
or U946 (N_946,In_421,In_838);
nand U947 (N_947,In_471,In_12);
nor U948 (N_948,In_328,In_120);
nand U949 (N_949,In_255,In_450);
or U950 (N_950,In_60,In_174);
nor U951 (N_951,In_215,In_14);
nand U952 (N_952,In_724,In_513);
or U953 (N_953,In_887,In_26);
or U954 (N_954,In_384,In_8);
and U955 (N_955,In_554,In_469);
or U956 (N_956,In_633,In_837);
nand U957 (N_957,In_156,In_439);
or U958 (N_958,In_293,In_193);
or U959 (N_959,In_10,In_560);
nor U960 (N_960,In_322,In_563);
and U961 (N_961,In_54,In_118);
or U962 (N_962,In_127,In_256);
xnor U963 (N_963,In_136,In_297);
nand U964 (N_964,In_781,In_799);
nor U965 (N_965,In_184,In_760);
nand U966 (N_966,In_732,In_251);
and U967 (N_967,In_865,In_914);
nand U968 (N_968,In_627,In_315);
nand U969 (N_969,In_184,In_467);
nand U970 (N_970,In_989,In_405);
nand U971 (N_971,In_757,In_660);
or U972 (N_972,In_46,In_809);
nor U973 (N_973,In_274,In_614);
nor U974 (N_974,In_273,In_326);
and U975 (N_975,In_318,In_189);
and U976 (N_976,In_976,In_337);
and U977 (N_977,In_426,In_411);
and U978 (N_978,In_737,In_714);
or U979 (N_979,In_441,In_4);
and U980 (N_980,In_361,In_329);
and U981 (N_981,In_905,In_383);
nand U982 (N_982,In_280,In_156);
nand U983 (N_983,In_634,In_44);
or U984 (N_984,In_249,In_540);
or U985 (N_985,In_354,In_924);
or U986 (N_986,In_193,In_486);
or U987 (N_987,In_635,In_563);
or U988 (N_988,In_863,In_376);
and U989 (N_989,In_934,In_838);
nand U990 (N_990,In_941,In_649);
nor U991 (N_991,In_841,In_609);
nor U992 (N_992,In_187,In_818);
nor U993 (N_993,In_372,In_188);
nand U994 (N_994,In_781,In_49);
nand U995 (N_995,In_753,In_257);
nand U996 (N_996,In_124,In_897);
nand U997 (N_997,In_419,In_943);
or U998 (N_998,In_690,In_435);
nand U999 (N_999,In_658,In_282);
nand U1000 (N_1000,N_192,N_44);
nand U1001 (N_1001,N_349,N_686);
nand U1002 (N_1002,N_858,N_391);
nor U1003 (N_1003,N_143,N_559);
nand U1004 (N_1004,N_567,N_377);
nor U1005 (N_1005,N_325,N_129);
or U1006 (N_1006,N_658,N_132);
and U1007 (N_1007,N_303,N_948);
nor U1008 (N_1008,N_824,N_262);
xor U1009 (N_1009,N_964,N_615);
and U1010 (N_1010,N_447,N_563);
and U1011 (N_1011,N_697,N_694);
and U1012 (N_1012,N_234,N_779);
nor U1013 (N_1013,N_238,N_855);
nor U1014 (N_1014,N_908,N_154);
nand U1015 (N_1015,N_628,N_860);
and U1016 (N_1016,N_937,N_347);
and U1017 (N_1017,N_576,N_570);
nand U1018 (N_1018,N_895,N_804);
nand U1019 (N_1019,N_983,N_420);
nand U1020 (N_1020,N_6,N_604);
and U1021 (N_1021,N_105,N_621);
nor U1022 (N_1022,N_654,N_987);
and U1023 (N_1023,N_373,N_75);
and U1024 (N_1024,N_287,N_513);
and U1025 (N_1025,N_643,N_700);
nor U1026 (N_1026,N_137,N_423);
nand U1027 (N_1027,N_297,N_729);
and U1028 (N_1028,N_20,N_32);
nand U1029 (N_1029,N_501,N_190);
or U1030 (N_1030,N_560,N_655);
nand U1031 (N_1031,N_225,N_722);
or U1032 (N_1032,N_889,N_668);
and U1033 (N_1033,N_726,N_758);
nand U1034 (N_1034,N_87,N_947);
and U1035 (N_1035,N_81,N_69);
or U1036 (N_1036,N_134,N_293);
or U1037 (N_1037,N_631,N_892);
nor U1038 (N_1038,N_395,N_484);
and U1039 (N_1039,N_408,N_728);
nand U1040 (N_1040,N_483,N_845);
or U1041 (N_1041,N_684,N_381);
nor U1042 (N_1042,N_19,N_323);
nand U1043 (N_1043,N_650,N_723);
nand U1044 (N_1044,N_317,N_548);
or U1045 (N_1045,N_685,N_91);
nor U1046 (N_1046,N_847,N_690);
and U1047 (N_1047,N_2,N_691);
nand U1048 (N_1048,N_575,N_837);
or U1049 (N_1049,N_836,N_304);
or U1050 (N_1050,N_56,N_789);
nor U1051 (N_1051,N_394,N_520);
or U1052 (N_1052,N_295,N_857);
nor U1053 (N_1053,N_22,N_361);
or U1054 (N_1054,N_122,N_438);
and U1055 (N_1055,N_308,N_276);
or U1056 (N_1056,N_644,N_663);
and U1057 (N_1057,N_653,N_107);
and U1058 (N_1058,N_339,N_637);
nor U1059 (N_1059,N_128,N_738);
and U1060 (N_1060,N_616,N_121);
nor U1061 (N_1061,N_750,N_707);
nor U1062 (N_1062,N_975,N_526);
nor U1063 (N_1063,N_98,N_550);
nor U1064 (N_1064,N_430,N_24);
xnor U1065 (N_1065,N_573,N_278);
nand U1066 (N_1066,N_819,N_961);
nand U1067 (N_1067,N_929,N_138);
or U1068 (N_1068,N_479,N_353);
nor U1069 (N_1069,N_301,N_827);
nor U1070 (N_1070,N_850,N_392);
and U1071 (N_1071,N_16,N_418);
and U1072 (N_1072,N_578,N_792);
nor U1073 (N_1073,N_133,N_798);
nand U1074 (N_1074,N_508,N_907);
or U1075 (N_1075,N_571,N_195);
and U1076 (N_1076,N_42,N_842);
or U1077 (N_1077,N_759,N_939);
nor U1078 (N_1078,N_329,N_248);
or U1079 (N_1079,N_481,N_568);
and U1080 (N_1080,N_485,N_613);
and U1081 (N_1081,N_246,N_147);
nor U1082 (N_1082,N_358,N_498);
nor U1083 (N_1083,N_510,N_296);
nor U1084 (N_1084,N_523,N_181);
nand U1085 (N_1085,N_218,N_184);
or U1086 (N_1086,N_635,N_396);
nor U1087 (N_1087,N_76,N_936);
xnor U1088 (N_1088,N_564,N_232);
nand U1089 (N_1089,N_117,N_84);
nand U1090 (N_1090,N_865,N_856);
or U1091 (N_1091,N_923,N_74);
nor U1092 (N_1092,N_477,N_187);
nor U1093 (N_1093,N_66,N_351);
and U1094 (N_1094,N_743,N_490);
nand U1095 (N_1095,N_572,N_18);
and U1096 (N_1096,N_906,N_168);
nor U1097 (N_1097,N_191,N_413);
nor U1098 (N_1098,N_846,N_673);
nor U1099 (N_1099,N_404,N_424);
nor U1100 (N_1100,N_415,N_51);
nor U1101 (N_1101,N_566,N_551);
and U1102 (N_1102,N_769,N_712);
xnor U1103 (N_1103,N_155,N_272);
nand U1104 (N_1104,N_884,N_183);
and U1105 (N_1105,N_125,N_815);
nor U1106 (N_1106,N_886,N_590);
and U1107 (N_1107,N_957,N_687);
nand U1108 (N_1108,N_749,N_145);
nor U1109 (N_1109,N_768,N_33);
nor U1110 (N_1110,N_878,N_896);
nor U1111 (N_1111,N_221,N_940);
nand U1112 (N_1112,N_338,N_163);
or U1113 (N_1113,N_113,N_201);
nor U1114 (N_1114,N_370,N_103);
nand U1115 (N_1115,N_453,N_166);
nand U1116 (N_1116,N_503,N_718);
and U1117 (N_1117,N_693,N_933);
or U1118 (N_1118,N_286,N_397);
nand U1119 (N_1119,N_289,N_164);
and U1120 (N_1120,N_368,N_336);
nor U1121 (N_1121,N_342,N_375);
or U1122 (N_1122,N_812,N_390);
xnor U1123 (N_1123,N_814,N_607);
and U1124 (N_1124,N_215,N_671);
nand U1125 (N_1125,N_49,N_417);
or U1126 (N_1126,N_3,N_588);
nand U1127 (N_1127,N_497,N_156);
and U1128 (N_1128,N_974,N_989);
xor U1129 (N_1129,N_0,N_680);
xor U1130 (N_1130,N_844,N_151);
nor U1131 (N_1131,N_206,N_148);
and U1132 (N_1132,N_997,N_640);
nand U1133 (N_1133,N_782,N_705);
nor U1134 (N_1134,N_786,N_67);
or U1135 (N_1135,N_322,N_874);
or U1136 (N_1136,N_612,N_902);
nor U1137 (N_1137,N_597,N_403);
nand U1138 (N_1138,N_161,N_582);
nor U1139 (N_1139,N_364,N_665);
nor U1140 (N_1140,N_826,N_434);
or U1141 (N_1141,N_152,N_231);
or U1142 (N_1142,N_745,N_314);
nand U1143 (N_1143,N_435,N_126);
nor U1144 (N_1144,N_530,N_139);
and U1145 (N_1145,N_808,N_606);
nor U1146 (N_1146,N_801,N_492);
and U1147 (N_1147,N_493,N_244);
and U1148 (N_1148,N_747,N_639);
or U1149 (N_1149,N_710,N_73);
nand U1150 (N_1150,N_407,N_79);
nor U1151 (N_1151,N_48,N_185);
and U1152 (N_1152,N_159,N_527);
or U1153 (N_1153,N_647,N_399);
and U1154 (N_1154,N_656,N_95);
or U1155 (N_1155,N_379,N_883);
nor U1156 (N_1156,N_414,N_901);
and U1157 (N_1157,N_505,N_871);
and U1158 (N_1158,N_952,N_822);
and U1159 (N_1159,N_21,N_380);
or U1160 (N_1160,N_514,N_701);
and U1161 (N_1161,N_809,N_714);
nand U1162 (N_1162,N_800,N_715);
nand U1163 (N_1163,N_834,N_692);
nor U1164 (N_1164,N_97,N_796);
and U1165 (N_1165,N_835,N_868);
and U1166 (N_1166,N_799,N_315);
nor U1167 (N_1167,N_806,N_976);
xor U1168 (N_1168,N_241,N_569);
or U1169 (N_1169,N_545,N_471);
or U1170 (N_1170,N_695,N_609);
and U1171 (N_1171,N_764,N_446);
and U1172 (N_1172,N_869,N_867);
or U1173 (N_1173,N_816,N_533);
or U1174 (N_1174,N_599,N_893);
and U1175 (N_1175,N_367,N_864);
nand U1176 (N_1176,N_35,N_197);
and U1177 (N_1177,N_13,N_45);
and U1178 (N_1178,N_131,N_735);
nor U1179 (N_1179,N_38,N_112);
nand U1180 (N_1180,N_502,N_316);
nand U1181 (N_1181,N_267,N_130);
and U1182 (N_1182,N_925,N_730);
and U1183 (N_1183,N_223,N_667);
nand U1184 (N_1184,N_626,N_919);
nor U1185 (N_1185,N_186,N_270);
nand U1186 (N_1186,N_12,N_558);
or U1187 (N_1187,N_802,N_746);
and U1188 (N_1188,N_877,N_401);
or U1189 (N_1189,N_384,N_124);
nand U1190 (N_1190,N_775,N_553);
and U1191 (N_1191,N_998,N_557);
or U1192 (N_1192,N_666,N_229);
nor U1193 (N_1193,N_954,N_217);
nor U1194 (N_1194,N_70,N_284);
nor U1195 (N_1195,N_465,N_509);
nor U1196 (N_1196,N_160,N_180);
nor U1197 (N_1197,N_172,N_115);
or U1198 (N_1198,N_972,N_648);
nand U1199 (N_1199,N_698,N_529);
and U1200 (N_1200,N_271,N_50);
or U1201 (N_1201,N_788,N_452);
or U1202 (N_1202,N_910,N_535);
and U1203 (N_1203,N_602,N_178);
or U1204 (N_1204,N_849,N_744);
and U1205 (N_1205,N_641,N_818);
xor U1206 (N_1206,N_751,N_670);
nand U1207 (N_1207,N_990,N_382);
and U1208 (N_1208,N_277,N_354);
nand U1209 (N_1209,N_15,N_611);
or U1210 (N_1210,N_903,N_158);
and U1211 (N_1211,N_862,N_623);
nand U1212 (N_1212,N_118,N_887);
nand U1213 (N_1213,N_562,N_475);
nor U1214 (N_1214,N_682,N_92);
and U1215 (N_1215,N_26,N_771);
nor U1216 (N_1216,N_486,N_922);
nor U1217 (N_1217,N_879,N_524);
nor U1218 (N_1218,N_27,N_805);
and U1219 (N_1219,N_935,N_68);
or U1220 (N_1220,N_25,N_332);
or U1221 (N_1221,N_448,N_546);
or U1222 (N_1222,N_696,N_931);
or U1223 (N_1223,N_672,N_760);
nand U1224 (N_1224,N_71,N_94);
xor U1225 (N_1225,N_83,N_460);
nor U1226 (N_1226,N_721,N_978);
or U1227 (N_1227,N_511,N_817);
and U1228 (N_1228,N_247,N_737);
nor U1229 (N_1229,N_268,N_203);
and U1230 (N_1230,N_324,N_425);
nand U1231 (N_1231,N_646,N_515);
or U1232 (N_1232,N_982,N_480);
or U1233 (N_1233,N_212,N_675);
xor U1234 (N_1234,N_104,N_402);
nand U1235 (N_1235,N_708,N_393);
and U1236 (N_1236,N_622,N_872);
or U1237 (N_1237,N_59,N_594);
nor U1238 (N_1238,N_752,N_863);
nand U1239 (N_1239,N_433,N_911);
nand U1240 (N_1240,N_36,N_388);
or U1241 (N_1241,N_372,N_734);
nor U1242 (N_1242,N_210,N_756);
and U1243 (N_1243,N_299,N_713);
and U1244 (N_1244,N_307,N_106);
or U1245 (N_1245,N_891,N_633);
xnor U1246 (N_1246,N_488,N_114);
nand U1247 (N_1247,N_90,N_135);
and U1248 (N_1248,N_699,N_472);
nand U1249 (N_1249,N_755,N_165);
or U1250 (N_1250,N_400,N_432);
nand U1251 (N_1251,N_679,N_440);
nand U1252 (N_1252,N_285,N_333);
or U1253 (N_1253,N_449,N_93);
nand U1254 (N_1254,N_521,N_476);
nand U1255 (N_1255,N_162,N_281);
nor U1256 (N_1256,N_984,N_320);
and U1257 (N_1257,N_598,N_740);
nor U1258 (N_1258,N_263,N_64);
or U1259 (N_1259,N_774,N_848);
nor U1260 (N_1260,N_427,N_732);
nor U1261 (N_1261,N_866,N_385);
nand U1262 (N_1262,N_992,N_220);
nand U1263 (N_1263,N_146,N_346);
and U1264 (N_1264,N_683,N_959);
or U1265 (N_1265,N_43,N_383);
and U1266 (N_1266,N_763,N_651);
nand U1267 (N_1267,N_150,N_830);
and U1268 (N_1268,N_96,N_915);
and U1269 (N_1269,N_345,N_99);
and U1270 (N_1270,N_620,N_116);
nor U1271 (N_1271,N_111,N_23);
or U1272 (N_1272,N_312,N_859);
and U1273 (N_1273,N_674,N_555);
nand U1274 (N_1274,N_260,N_932);
nor U1275 (N_1275,N_885,N_795);
nor U1276 (N_1276,N_525,N_945);
nand U1277 (N_1277,N_494,N_634);
xor U1278 (N_1278,N_11,N_426);
nor U1279 (N_1279,N_214,N_781);
nand U1280 (N_1280,N_854,N_642);
nand U1281 (N_1281,N_870,N_4);
nand U1282 (N_1282,N_953,N_914);
and U1283 (N_1283,N_742,N_532);
nor U1284 (N_1284,N_980,N_706);
or U1285 (N_1285,N_366,N_956);
nand U1286 (N_1286,N_765,N_776);
or U1287 (N_1287,N_709,N_888);
nand U1288 (N_1288,N_662,N_264);
and U1289 (N_1289,N_343,N_140);
nor U1290 (N_1290,N_60,N_52);
and U1291 (N_1291,N_177,N_950);
nor U1292 (N_1292,N_843,N_319);
or U1293 (N_1293,N_409,N_274);
nor U1294 (N_1294,N_337,N_282);
and U1295 (N_1295,N_321,N_627);
and U1296 (N_1296,N_256,N_359);
or U1297 (N_1297,N_554,N_944);
nand U1298 (N_1298,N_72,N_958);
or U1299 (N_1299,N_504,N_739);
and U1300 (N_1300,N_938,N_240);
nor U1301 (N_1301,N_176,N_233);
nor U1302 (N_1302,N_678,N_995);
and U1303 (N_1303,N_283,N_14);
and U1304 (N_1304,N_77,N_927);
and U1305 (N_1305,N_519,N_930);
and U1306 (N_1306,N_335,N_474);
nor U1307 (N_1307,N_577,N_890);
nand U1308 (N_1308,N_136,N_783);
nor U1309 (N_1309,N_470,N_290);
nor U1310 (N_1310,N_873,N_790);
nor U1311 (N_1311,N_688,N_996);
nand U1312 (N_1312,N_820,N_54);
or U1313 (N_1313,N_61,N_926);
or U1314 (N_1314,N_587,N_450);
nand U1315 (N_1315,N_369,N_838);
or U1316 (N_1316,N_119,N_552);
and U1317 (N_1317,N_542,N_258);
nand U1318 (N_1318,N_716,N_199);
or U1319 (N_1319,N_37,N_561);
nand U1320 (N_1320,N_605,N_239);
and U1321 (N_1321,N_142,N_78);
or U1322 (N_1322,N_811,N_211);
and U1323 (N_1323,N_149,N_179);
nor U1324 (N_1324,N_610,N_664);
nor U1325 (N_1325,N_861,N_254);
nand U1326 (N_1326,N_311,N_853);
nor U1327 (N_1327,N_951,N_600);
and U1328 (N_1328,N_540,N_534);
nand U1329 (N_1329,N_968,N_541);
or U1330 (N_1330,N_265,N_832);
nand U1331 (N_1331,N_89,N_757);
and U1332 (N_1332,N_657,N_702);
nand U1333 (N_1333,N_979,N_897);
nor U1334 (N_1334,N_292,N_300);
nor U1335 (N_1335,N_473,N_917);
or U1336 (N_1336,N_288,N_144);
nand U1337 (N_1337,N_778,N_57);
and U1338 (N_1338,N_522,N_1);
xor U1339 (N_1339,N_591,N_157);
nand U1340 (N_1340,N_608,N_330);
nand U1341 (N_1341,N_916,N_468);
or U1342 (N_1342,N_88,N_326);
nand U1343 (N_1343,N_437,N_120);
nand U1344 (N_1344,N_833,N_467);
nand U1345 (N_1345,N_921,N_389);
nand U1346 (N_1346,N_825,N_894);
or U1347 (N_1347,N_243,N_8);
xnor U1348 (N_1348,N_279,N_362);
and U1349 (N_1349,N_603,N_251);
and U1350 (N_1350,N_363,N_762);
nand U1351 (N_1351,N_309,N_823);
and U1352 (N_1352,N_273,N_518);
or U1353 (N_1353,N_660,N_770);
nor U1354 (N_1354,N_882,N_422);
or U1355 (N_1355,N_596,N_766);
nor U1356 (N_1356,N_405,N_153);
and U1357 (N_1357,N_242,N_249);
nand U1358 (N_1358,N_986,N_110);
and U1359 (N_1359,N_618,N_205);
nand U1360 (N_1360,N_506,N_200);
nand U1361 (N_1361,N_767,N_585);
or U1362 (N_1362,N_410,N_720);
and U1363 (N_1363,N_967,N_507);
or U1364 (N_1364,N_202,N_291);
nand U1365 (N_1365,N_579,N_207);
and U1366 (N_1366,N_188,N_661);
and U1367 (N_1367,N_193,N_31);
or U1368 (N_1368,N_840,N_638);
nor U1369 (N_1369,N_985,N_294);
nor U1370 (N_1370,N_965,N_348);
xnor U1371 (N_1371,N_516,N_970);
and U1372 (N_1372,N_574,N_416);
nor U1373 (N_1373,N_17,N_9);
nand U1374 (N_1374,N_780,N_583);
and U1375 (N_1375,N_85,N_334);
nand U1376 (N_1376,N_645,N_428);
nor U1377 (N_1377,N_681,N_466);
nand U1378 (N_1378,N_298,N_841);
nor U1379 (N_1379,N_39,N_275);
nor U1380 (N_1380,N_724,N_973);
or U1381 (N_1381,N_717,N_556);
nor U1382 (N_1382,N_630,N_960);
nor U1383 (N_1383,N_100,N_318);
or U1384 (N_1384,N_436,N_269);
and U1385 (N_1385,N_443,N_528);
and U1386 (N_1386,N_941,N_360);
nor U1387 (N_1387,N_456,N_439);
nor U1388 (N_1388,N_549,N_629);
nand U1389 (N_1389,N_198,N_109);
or U1390 (N_1390,N_669,N_966);
and U1391 (N_1391,N_880,N_753);
or U1392 (N_1392,N_170,N_34);
nor U1393 (N_1393,N_761,N_398);
xnor U1394 (N_1394,N_305,N_876);
nand U1395 (N_1395,N_994,N_371);
nor U1396 (N_1396,N_881,N_459);
or U1397 (N_1397,N_257,N_127);
nor U1398 (N_1398,N_208,N_614);
or U1399 (N_1399,N_544,N_536);
and U1400 (N_1400,N_543,N_727);
nand U1401 (N_1401,N_733,N_387);
nand U1402 (N_1402,N_539,N_235);
and U1403 (N_1403,N_80,N_65);
xnor U1404 (N_1404,N_592,N_141);
xor U1405 (N_1405,N_174,N_928);
or U1406 (N_1406,N_341,N_245);
or U1407 (N_1407,N_386,N_946);
xnor U1408 (N_1408,N_352,N_624);
nor U1409 (N_1409,N_365,N_7);
or U1410 (N_1410,N_357,N_236);
nor U1411 (N_1411,N_828,N_189);
and U1412 (N_1412,N_376,N_169);
nand U1413 (N_1413,N_586,N_632);
nor U1414 (N_1414,N_204,N_489);
and U1415 (N_1415,N_704,N_123);
nor U1416 (N_1416,N_495,N_491);
and U1417 (N_1417,N_302,N_182);
nor U1418 (N_1418,N_306,N_455);
nor U1419 (N_1419,N_10,N_898);
or U1420 (N_1420,N_313,N_942);
nand U1421 (N_1421,N_444,N_565);
nor U1422 (N_1422,N_82,N_617);
and U1423 (N_1423,N_374,N_787);
and U1424 (N_1424,N_216,N_175);
nand U1425 (N_1425,N_580,N_962);
and U1426 (N_1426,N_821,N_625);
nor U1427 (N_1427,N_259,N_463);
or U1428 (N_1428,N_237,N_595);
nor U1429 (N_1429,N_458,N_659);
or U1430 (N_1430,N_676,N_62);
and U1431 (N_1431,N_41,N_266);
nor U1432 (N_1432,N_839,N_711);
nand U1433 (N_1433,N_904,N_601);
nand U1434 (N_1434,N_803,N_46);
or U1435 (N_1435,N_356,N_900);
or U1436 (N_1436,N_652,N_496);
or U1437 (N_1437,N_943,N_981);
or U1438 (N_1438,N_547,N_280);
and U1439 (N_1439,N_253,N_327);
nor U1440 (N_1440,N_852,N_677);
nand U1441 (N_1441,N_171,N_86);
nor U1442 (N_1442,N_794,N_793);
and U1443 (N_1443,N_754,N_807);
nor U1444 (N_1444,N_512,N_28);
or U1445 (N_1445,N_797,N_167);
nor U1446 (N_1446,N_331,N_102);
nor U1447 (N_1447,N_636,N_40);
and U1448 (N_1448,N_411,N_228);
xnor U1449 (N_1449,N_920,N_487);
nand U1450 (N_1450,N_255,N_589);
nor U1451 (N_1451,N_581,N_649);
or U1452 (N_1452,N_194,N_227);
or U1453 (N_1453,N_810,N_785);
and U1454 (N_1454,N_791,N_538);
and U1455 (N_1455,N_913,N_209);
nand U1456 (N_1456,N_991,N_482);
nand U1457 (N_1457,N_350,N_47);
or U1458 (N_1458,N_328,N_53);
nor U1459 (N_1459,N_457,N_988);
or U1460 (N_1460,N_213,N_531);
nand U1461 (N_1461,N_777,N_773);
nand U1462 (N_1462,N_934,N_955);
nand U1463 (N_1463,N_55,N_619);
or U1464 (N_1464,N_784,N_378);
nand U1465 (N_1465,N_689,N_593);
nor U1466 (N_1466,N_478,N_261);
nor U1467 (N_1467,N_5,N_537);
and U1468 (N_1468,N_462,N_340);
nand U1469 (N_1469,N_442,N_58);
nand U1470 (N_1470,N_993,N_431);
nand U1471 (N_1471,N_222,N_899);
and U1472 (N_1472,N_406,N_741);
nor U1473 (N_1473,N_451,N_310);
or U1474 (N_1474,N_108,N_250);
and U1475 (N_1475,N_252,N_905);
and U1476 (N_1476,N_909,N_999);
and U1477 (N_1477,N_963,N_918);
and U1478 (N_1478,N_464,N_412);
nor U1479 (N_1479,N_731,N_829);
nor U1480 (N_1480,N_748,N_971);
nand U1481 (N_1481,N_703,N_736);
and U1482 (N_1482,N_429,N_454);
and U1483 (N_1483,N_469,N_969);
nand U1484 (N_1484,N_173,N_355);
nand U1485 (N_1485,N_912,N_344);
or U1486 (N_1486,N_441,N_230);
nor U1487 (N_1487,N_224,N_461);
nor U1488 (N_1488,N_499,N_419);
and U1489 (N_1489,N_949,N_772);
and U1490 (N_1490,N_813,N_584);
and U1491 (N_1491,N_445,N_63);
or U1492 (N_1492,N_851,N_196);
nand U1493 (N_1493,N_219,N_517);
or U1494 (N_1494,N_30,N_924);
and U1495 (N_1495,N_831,N_875);
nor U1496 (N_1496,N_719,N_977);
nand U1497 (N_1497,N_226,N_29);
or U1498 (N_1498,N_101,N_500);
or U1499 (N_1499,N_421,N_725);
and U1500 (N_1500,N_905,N_873);
or U1501 (N_1501,N_81,N_490);
nand U1502 (N_1502,N_476,N_985);
or U1503 (N_1503,N_90,N_602);
or U1504 (N_1504,N_737,N_836);
or U1505 (N_1505,N_487,N_55);
nand U1506 (N_1506,N_40,N_269);
nor U1507 (N_1507,N_775,N_146);
and U1508 (N_1508,N_465,N_957);
and U1509 (N_1509,N_605,N_14);
and U1510 (N_1510,N_37,N_116);
nor U1511 (N_1511,N_683,N_135);
and U1512 (N_1512,N_102,N_309);
or U1513 (N_1513,N_12,N_911);
or U1514 (N_1514,N_36,N_515);
nor U1515 (N_1515,N_660,N_411);
or U1516 (N_1516,N_327,N_136);
or U1517 (N_1517,N_172,N_933);
nor U1518 (N_1518,N_715,N_355);
nor U1519 (N_1519,N_245,N_870);
nor U1520 (N_1520,N_815,N_932);
and U1521 (N_1521,N_798,N_831);
and U1522 (N_1522,N_612,N_267);
nand U1523 (N_1523,N_98,N_940);
and U1524 (N_1524,N_925,N_697);
nand U1525 (N_1525,N_63,N_97);
and U1526 (N_1526,N_658,N_647);
or U1527 (N_1527,N_891,N_56);
nand U1528 (N_1528,N_545,N_602);
nor U1529 (N_1529,N_17,N_767);
nand U1530 (N_1530,N_497,N_739);
nand U1531 (N_1531,N_776,N_302);
or U1532 (N_1532,N_266,N_480);
nor U1533 (N_1533,N_461,N_542);
or U1534 (N_1534,N_326,N_970);
and U1535 (N_1535,N_443,N_43);
nand U1536 (N_1536,N_100,N_542);
or U1537 (N_1537,N_546,N_366);
and U1538 (N_1538,N_175,N_981);
or U1539 (N_1539,N_121,N_793);
and U1540 (N_1540,N_386,N_755);
and U1541 (N_1541,N_201,N_926);
or U1542 (N_1542,N_662,N_536);
nand U1543 (N_1543,N_281,N_855);
and U1544 (N_1544,N_310,N_170);
nor U1545 (N_1545,N_291,N_846);
nand U1546 (N_1546,N_102,N_764);
and U1547 (N_1547,N_487,N_662);
and U1548 (N_1548,N_307,N_131);
nand U1549 (N_1549,N_469,N_705);
nor U1550 (N_1550,N_537,N_360);
and U1551 (N_1551,N_705,N_66);
nor U1552 (N_1552,N_790,N_439);
nand U1553 (N_1553,N_452,N_422);
nor U1554 (N_1554,N_953,N_881);
and U1555 (N_1555,N_860,N_943);
or U1556 (N_1556,N_883,N_723);
xor U1557 (N_1557,N_394,N_422);
or U1558 (N_1558,N_883,N_143);
nand U1559 (N_1559,N_57,N_402);
nor U1560 (N_1560,N_754,N_798);
nor U1561 (N_1561,N_452,N_612);
nor U1562 (N_1562,N_865,N_612);
nor U1563 (N_1563,N_207,N_903);
and U1564 (N_1564,N_674,N_255);
or U1565 (N_1565,N_919,N_295);
nor U1566 (N_1566,N_151,N_803);
and U1567 (N_1567,N_801,N_809);
and U1568 (N_1568,N_683,N_481);
xnor U1569 (N_1569,N_257,N_487);
nand U1570 (N_1570,N_638,N_165);
nor U1571 (N_1571,N_847,N_292);
nand U1572 (N_1572,N_663,N_821);
and U1573 (N_1573,N_346,N_557);
or U1574 (N_1574,N_340,N_704);
nand U1575 (N_1575,N_496,N_239);
and U1576 (N_1576,N_935,N_377);
or U1577 (N_1577,N_993,N_689);
and U1578 (N_1578,N_279,N_457);
nor U1579 (N_1579,N_697,N_12);
nor U1580 (N_1580,N_44,N_431);
and U1581 (N_1581,N_899,N_142);
and U1582 (N_1582,N_848,N_381);
nand U1583 (N_1583,N_417,N_626);
nor U1584 (N_1584,N_478,N_955);
and U1585 (N_1585,N_789,N_223);
xor U1586 (N_1586,N_374,N_738);
nand U1587 (N_1587,N_699,N_751);
and U1588 (N_1588,N_929,N_391);
and U1589 (N_1589,N_408,N_394);
nand U1590 (N_1590,N_30,N_415);
nor U1591 (N_1591,N_396,N_584);
nor U1592 (N_1592,N_13,N_351);
or U1593 (N_1593,N_300,N_417);
or U1594 (N_1594,N_240,N_492);
or U1595 (N_1595,N_837,N_54);
and U1596 (N_1596,N_182,N_449);
or U1597 (N_1597,N_634,N_756);
or U1598 (N_1598,N_542,N_587);
and U1599 (N_1599,N_661,N_664);
nand U1600 (N_1600,N_932,N_575);
and U1601 (N_1601,N_816,N_288);
nand U1602 (N_1602,N_47,N_734);
and U1603 (N_1603,N_399,N_245);
or U1604 (N_1604,N_139,N_257);
nand U1605 (N_1605,N_430,N_316);
and U1606 (N_1606,N_557,N_443);
nor U1607 (N_1607,N_822,N_184);
or U1608 (N_1608,N_584,N_353);
nor U1609 (N_1609,N_108,N_805);
or U1610 (N_1610,N_460,N_900);
nor U1611 (N_1611,N_893,N_70);
or U1612 (N_1612,N_720,N_146);
nand U1613 (N_1613,N_603,N_961);
or U1614 (N_1614,N_395,N_733);
nand U1615 (N_1615,N_799,N_378);
or U1616 (N_1616,N_979,N_424);
and U1617 (N_1617,N_463,N_419);
nand U1618 (N_1618,N_421,N_275);
and U1619 (N_1619,N_874,N_818);
nor U1620 (N_1620,N_483,N_327);
nor U1621 (N_1621,N_135,N_371);
nand U1622 (N_1622,N_571,N_760);
nor U1623 (N_1623,N_389,N_685);
nor U1624 (N_1624,N_572,N_166);
nand U1625 (N_1625,N_121,N_488);
nor U1626 (N_1626,N_193,N_410);
nor U1627 (N_1627,N_955,N_438);
nor U1628 (N_1628,N_386,N_779);
or U1629 (N_1629,N_183,N_629);
nand U1630 (N_1630,N_569,N_167);
or U1631 (N_1631,N_570,N_836);
and U1632 (N_1632,N_780,N_745);
xnor U1633 (N_1633,N_519,N_218);
nand U1634 (N_1634,N_750,N_674);
nor U1635 (N_1635,N_825,N_527);
nor U1636 (N_1636,N_818,N_250);
nand U1637 (N_1637,N_511,N_743);
or U1638 (N_1638,N_471,N_71);
or U1639 (N_1639,N_403,N_526);
and U1640 (N_1640,N_164,N_324);
and U1641 (N_1641,N_617,N_751);
xnor U1642 (N_1642,N_461,N_427);
and U1643 (N_1643,N_507,N_958);
and U1644 (N_1644,N_59,N_300);
nand U1645 (N_1645,N_702,N_998);
nand U1646 (N_1646,N_818,N_220);
or U1647 (N_1647,N_333,N_395);
and U1648 (N_1648,N_961,N_256);
nand U1649 (N_1649,N_900,N_535);
and U1650 (N_1650,N_149,N_325);
and U1651 (N_1651,N_350,N_235);
or U1652 (N_1652,N_651,N_929);
nand U1653 (N_1653,N_445,N_78);
and U1654 (N_1654,N_461,N_800);
and U1655 (N_1655,N_759,N_382);
nor U1656 (N_1656,N_532,N_48);
nor U1657 (N_1657,N_322,N_887);
and U1658 (N_1658,N_957,N_431);
nor U1659 (N_1659,N_973,N_512);
nor U1660 (N_1660,N_139,N_0);
xor U1661 (N_1661,N_58,N_120);
and U1662 (N_1662,N_576,N_577);
or U1663 (N_1663,N_509,N_269);
or U1664 (N_1664,N_90,N_232);
or U1665 (N_1665,N_621,N_682);
nand U1666 (N_1666,N_768,N_761);
nor U1667 (N_1667,N_77,N_622);
or U1668 (N_1668,N_636,N_844);
xnor U1669 (N_1669,N_680,N_361);
nor U1670 (N_1670,N_720,N_151);
and U1671 (N_1671,N_419,N_354);
nor U1672 (N_1672,N_673,N_714);
and U1673 (N_1673,N_864,N_263);
nor U1674 (N_1674,N_829,N_850);
nor U1675 (N_1675,N_22,N_375);
and U1676 (N_1676,N_128,N_508);
nor U1677 (N_1677,N_523,N_188);
or U1678 (N_1678,N_739,N_249);
and U1679 (N_1679,N_636,N_787);
nand U1680 (N_1680,N_888,N_992);
nand U1681 (N_1681,N_938,N_506);
or U1682 (N_1682,N_937,N_584);
and U1683 (N_1683,N_701,N_347);
or U1684 (N_1684,N_883,N_655);
nand U1685 (N_1685,N_607,N_80);
or U1686 (N_1686,N_694,N_314);
nor U1687 (N_1687,N_339,N_817);
and U1688 (N_1688,N_215,N_720);
or U1689 (N_1689,N_722,N_538);
and U1690 (N_1690,N_240,N_259);
or U1691 (N_1691,N_982,N_545);
nor U1692 (N_1692,N_72,N_582);
nor U1693 (N_1693,N_527,N_113);
or U1694 (N_1694,N_5,N_84);
or U1695 (N_1695,N_847,N_686);
and U1696 (N_1696,N_198,N_738);
or U1697 (N_1697,N_116,N_132);
nand U1698 (N_1698,N_301,N_263);
nor U1699 (N_1699,N_425,N_545);
and U1700 (N_1700,N_539,N_371);
nor U1701 (N_1701,N_605,N_428);
and U1702 (N_1702,N_917,N_902);
nand U1703 (N_1703,N_817,N_942);
nor U1704 (N_1704,N_959,N_638);
and U1705 (N_1705,N_454,N_990);
nor U1706 (N_1706,N_622,N_710);
nor U1707 (N_1707,N_645,N_629);
nor U1708 (N_1708,N_707,N_552);
or U1709 (N_1709,N_905,N_657);
xnor U1710 (N_1710,N_503,N_10);
nor U1711 (N_1711,N_120,N_729);
and U1712 (N_1712,N_164,N_911);
and U1713 (N_1713,N_894,N_334);
nor U1714 (N_1714,N_281,N_694);
or U1715 (N_1715,N_42,N_611);
nand U1716 (N_1716,N_783,N_849);
nand U1717 (N_1717,N_721,N_702);
nor U1718 (N_1718,N_675,N_594);
nand U1719 (N_1719,N_140,N_646);
or U1720 (N_1720,N_810,N_5);
nor U1721 (N_1721,N_35,N_487);
nand U1722 (N_1722,N_661,N_13);
nand U1723 (N_1723,N_389,N_808);
nand U1724 (N_1724,N_151,N_718);
nand U1725 (N_1725,N_709,N_473);
or U1726 (N_1726,N_365,N_343);
and U1727 (N_1727,N_701,N_722);
nor U1728 (N_1728,N_25,N_740);
or U1729 (N_1729,N_32,N_729);
and U1730 (N_1730,N_322,N_911);
and U1731 (N_1731,N_328,N_73);
nand U1732 (N_1732,N_95,N_381);
nand U1733 (N_1733,N_945,N_361);
and U1734 (N_1734,N_636,N_304);
nand U1735 (N_1735,N_200,N_299);
and U1736 (N_1736,N_305,N_977);
nor U1737 (N_1737,N_651,N_706);
or U1738 (N_1738,N_618,N_518);
nor U1739 (N_1739,N_849,N_183);
xnor U1740 (N_1740,N_468,N_135);
or U1741 (N_1741,N_810,N_884);
and U1742 (N_1742,N_270,N_598);
nor U1743 (N_1743,N_285,N_733);
or U1744 (N_1744,N_589,N_557);
nor U1745 (N_1745,N_740,N_601);
and U1746 (N_1746,N_157,N_317);
nor U1747 (N_1747,N_541,N_594);
or U1748 (N_1748,N_799,N_830);
and U1749 (N_1749,N_237,N_946);
nand U1750 (N_1750,N_539,N_185);
or U1751 (N_1751,N_510,N_4);
nand U1752 (N_1752,N_834,N_858);
and U1753 (N_1753,N_553,N_819);
and U1754 (N_1754,N_698,N_69);
or U1755 (N_1755,N_671,N_192);
or U1756 (N_1756,N_559,N_290);
and U1757 (N_1757,N_940,N_300);
nor U1758 (N_1758,N_146,N_939);
nand U1759 (N_1759,N_70,N_529);
nor U1760 (N_1760,N_241,N_915);
and U1761 (N_1761,N_652,N_57);
nand U1762 (N_1762,N_709,N_968);
or U1763 (N_1763,N_42,N_986);
xor U1764 (N_1764,N_448,N_210);
and U1765 (N_1765,N_417,N_9);
nor U1766 (N_1766,N_907,N_700);
or U1767 (N_1767,N_111,N_55);
or U1768 (N_1768,N_88,N_592);
xor U1769 (N_1769,N_312,N_14);
or U1770 (N_1770,N_467,N_636);
nand U1771 (N_1771,N_147,N_237);
or U1772 (N_1772,N_985,N_157);
nor U1773 (N_1773,N_761,N_778);
nand U1774 (N_1774,N_794,N_731);
and U1775 (N_1775,N_886,N_873);
or U1776 (N_1776,N_110,N_372);
and U1777 (N_1777,N_357,N_773);
or U1778 (N_1778,N_206,N_445);
nand U1779 (N_1779,N_122,N_454);
nor U1780 (N_1780,N_38,N_690);
nor U1781 (N_1781,N_872,N_735);
or U1782 (N_1782,N_694,N_557);
and U1783 (N_1783,N_151,N_23);
nor U1784 (N_1784,N_571,N_243);
and U1785 (N_1785,N_608,N_143);
nor U1786 (N_1786,N_18,N_415);
and U1787 (N_1787,N_91,N_483);
or U1788 (N_1788,N_353,N_432);
or U1789 (N_1789,N_581,N_762);
or U1790 (N_1790,N_186,N_236);
or U1791 (N_1791,N_348,N_240);
nor U1792 (N_1792,N_786,N_40);
and U1793 (N_1793,N_666,N_954);
or U1794 (N_1794,N_940,N_864);
and U1795 (N_1795,N_200,N_637);
and U1796 (N_1796,N_649,N_255);
and U1797 (N_1797,N_169,N_13);
nor U1798 (N_1798,N_487,N_892);
or U1799 (N_1799,N_213,N_82);
and U1800 (N_1800,N_102,N_242);
or U1801 (N_1801,N_153,N_715);
nor U1802 (N_1802,N_55,N_17);
nor U1803 (N_1803,N_840,N_423);
nor U1804 (N_1804,N_274,N_994);
nor U1805 (N_1805,N_909,N_335);
and U1806 (N_1806,N_27,N_425);
nand U1807 (N_1807,N_20,N_757);
nor U1808 (N_1808,N_443,N_460);
nand U1809 (N_1809,N_345,N_500);
or U1810 (N_1810,N_336,N_278);
and U1811 (N_1811,N_800,N_225);
nor U1812 (N_1812,N_30,N_684);
and U1813 (N_1813,N_668,N_720);
or U1814 (N_1814,N_190,N_200);
and U1815 (N_1815,N_667,N_149);
nor U1816 (N_1816,N_915,N_361);
and U1817 (N_1817,N_796,N_711);
or U1818 (N_1818,N_377,N_372);
or U1819 (N_1819,N_301,N_812);
and U1820 (N_1820,N_765,N_159);
or U1821 (N_1821,N_984,N_894);
or U1822 (N_1822,N_483,N_738);
or U1823 (N_1823,N_780,N_982);
or U1824 (N_1824,N_212,N_390);
or U1825 (N_1825,N_500,N_606);
nand U1826 (N_1826,N_627,N_200);
or U1827 (N_1827,N_508,N_222);
and U1828 (N_1828,N_841,N_842);
nand U1829 (N_1829,N_559,N_820);
and U1830 (N_1830,N_200,N_993);
and U1831 (N_1831,N_749,N_281);
nor U1832 (N_1832,N_436,N_997);
or U1833 (N_1833,N_191,N_160);
nor U1834 (N_1834,N_232,N_975);
or U1835 (N_1835,N_442,N_858);
or U1836 (N_1836,N_380,N_638);
and U1837 (N_1837,N_66,N_375);
or U1838 (N_1838,N_239,N_597);
and U1839 (N_1839,N_798,N_62);
nand U1840 (N_1840,N_408,N_445);
or U1841 (N_1841,N_443,N_990);
or U1842 (N_1842,N_249,N_986);
nor U1843 (N_1843,N_855,N_954);
nor U1844 (N_1844,N_749,N_544);
nand U1845 (N_1845,N_667,N_727);
or U1846 (N_1846,N_581,N_318);
nor U1847 (N_1847,N_466,N_899);
nor U1848 (N_1848,N_584,N_910);
xnor U1849 (N_1849,N_358,N_517);
nor U1850 (N_1850,N_141,N_419);
and U1851 (N_1851,N_995,N_550);
nand U1852 (N_1852,N_134,N_449);
nand U1853 (N_1853,N_216,N_766);
nor U1854 (N_1854,N_950,N_587);
nand U1855 (N_1855,N_316,N_846);
and U1856 (N_1856,N_229,N_406);
nor U1857 (N_1857,N_695,N_796);
nand U1858 (N_1858,N_778,N_862);
or U1859 (N_1859,N_331,N_244);
and U1860 (N_1860,N_814,N_511);
nor U1861 (N_1861,N_540,N_935);
and U1862 (N_1862,N_498,N_638);
nor U1863 (N_1863,N_703,N_546);
nand U1864 (N_1864,N_340,N_655);
or U1865 (N_1865,N_548,N_543);
and U1866 (N_1866,N_555,N_377);
nand U1867 (N_1867,N_827,N_164);
nand U1868 (N_1868,N_380,N_387);
or U1869 (N_1869,N_599,N_81);
nor U1870 (N_1870,N_977,N_711);
xnor U1871 (N_1871,N_838,N_546);
nand U1872 (N_1872,N_616,N_331);
nor U1873 (N_1873,N_671,N_200);
nor U1874 (N_1874,N_690,N_471);
or U1875 (N_1875,N_784,N_96);
or U1876 (N_1876,N_584,N_425);
and U1877 (N_1877,N_90,N_916);
and U1878 (N_1878,N_847,N_7);
xor U1879 (N_1879,N_17,N_980);
nand U1880 (N_1880,N_548,N_836);
and U1881 (N_1881,N_48,N_584);
and U1882 (N_1882,N_117,N_50);
nor U1883 (N_1883,N_903,N_20);
nand U1884 (N_1884,N_43,N_750);
and U1885 (N_1885,N_828,N_53);
and U1886 (N_1886,N_836,N_987);
and U1887 (N_1887,N_876,N_357);
nand U1888 (N_1888,N_292,N_593);
nand U1889 (N_1889,N_288,N_199);
nor U1890 (N_1890,N_146,N_991);
and U1891 (N_1891,N_625,N_523);
and U1892 (N_1892,N_59,N_684);
and U1893 (N_1893,N_424,N_476);
or U1894 (N_1894,N_163,N_328);
nor U1895 (N_1895,N_995,N_245);
nand U1896 (N_1896,N_774,N_116);
nor U1897 (N_1897,N_342,N_660);
or U1898 (N_1898,N_537,N_691);
nand U1899 (N_1899,N_729,N_827);
or U1900 (N_1900,N_903,N_445);
nor U1901 (N_1901,N_19,N_929);
and U1902 (N_1902,N_343,N_215);
nand U1903 (N_1903,N_530,N_128);
or U1904 (N_1904,N_141,N_438);
nand U1905 (N_1905,N_20,N_373);
and U1906 (N_1906,N_672,N_970);
and U1907 (N_1907,N_464,N_61);
and U1908 (N_1908,N_566,N_307);
or U1909 (N_1909,N_107,N_965);
nor U1910 (N_1910,N_922,N_193);
or U1911 (N_1911,N_125,N_367);
nor U1912 (N_1912,N_26,N_355);
nor U1913 (N_1913,N_953,N_709);
nand U1914 (N_1914,N_807,N_155);
nand U1915 (N_1915,N_136,N_644);
or U1916 (N_1916,N_709,N_29);
nand U1917 (N_1917,N_990,N_347);
nor U1918 (N_1918,N_334,N_762);
nand U1919 (N_1919,N_404,N_799);
nand U1920 (N_1920,N_765,N_223);
nor U1921 (N_1921,N_897,N_332);
nor U1922 (N_1922,N_598,N_396);
and U1923 (N_1923,N_479,N_606);
and U1924 (N_1924,N_822,N_482);
and U1925 (N_1925,N_772,N_699);
nor U1926 (N_1926,N_816,N_562);
nor U1927 (N_1927,N_621,N_469);
nand U1928 (N_1928,N_933,N_507);
nor U1929 (N_1929,N_867,N_130);
nor U1930 (N_1930,N_185,N_833);
and U1931 (N_1931,N_678,N_481);
nor U1932 (N_1932,N_935,N_632);
and U1933 (N_1933,N_470,N_392);
and U1934 (N_1934,N_138,N_458);
nand U1935 (N_1935,N_631,N_436);
or U1936 (N_1936,N_760,N_957);
nor U1937 (N_1937,N_420,N_972);
and U1938 (N_1938,N_421,N_856);
and U1939 (N_1939,N_179,N_757);
nor U1940 (N_1940,N_557,N_485);
and U1941 (N_1941,N_313,N_429);
and U1942 (N_1942,N_424,N_926);
nor U1943 (N_1943,N_929,N_258);
nand U1944 (N_1944,N_219,N_863);
or U1945 (N_1945,N_358,N_142);
and U1946 (N_1946,N_247,N_170);
nand U1947 (N_1947,N_917,N_767);
and U1948 (N_1948,N_773,N_904);
nor U1949 (N_1949,N_158,N_11);
xnor U1950 (N_1950,N_840,N_843);
nor U1951 (N_1951,N_116,N_35);
nand U1952 (N_1952,N_797,N_745);
or U1953 (N_1953,N_959,N_1);
and U1954 (N_1954,N_619,N_785);
nand U1955 (N_1955,N_884,N_907);
and U1956 (N_1956,N_427,N_876);
nand U1957 (N_1957,N_872,N_581);
and U1958 (N_1958,N_899,N_411);
nor U1959 (N_1959,N_723,N_99);
nor U1960 (N_1960,N_773,N_8);
and U1961 (N_1961,N_834,N_957);
nand U1962 (N_1962,N_231,N_451);
nand U1963 (N_1963,N_199,N_652);
or U1964 (N_1964,N_652,N_989);
or U1965 (N_1965,N_91,N_721);
nor U1966 (N_1966,N_365,N_93);
and U1967 (N_1967,N_224,N_891);
or U1968 (N_1968,N_328,N_609);
and U1969 (N_1969,N_216,N_666);
nand U1970 (N_1970,N_852,N_29);
nand U1971 (N_1971,N_111,N_607);
nand U1972 (N_1972,N_586,N_948);
nor U1973 (N_1973,N_669,N_436);
nor U1974 (N_1974,N_672,N_236);
or U1975 (N_1975,N_297,N_915);
nor U1976 (N_1976,N_467,N_628);
and U1977 (N_1977,N_801,N_311);
xnor U1978 (N_1978,N_557,N_409);
nor U1979 (N_1979,N_871,N_590);
or U1980 (N_1980,N_402,N_325);
and U1981 (N_1981,N_397,N_254);
nor U1982 (N_1982,N_879,N_28);
and U1983 (N_1983,N_828,N_2);
and U1984 (N_1984,N_792,N_980);
and U1985 (N_1985,N_125,N_715);
nor U1986 (N_1986,N_476,N_312);
nand U1987 (N_1987,N_282,N_894);
nor U1988 (N_1988,N_270,N_160);
and U1989 (N_1989,N_761,N_552);
or U1990 (N_1990,N_513,N_929);
nor U1991 (N_1991,N_384,N_974);
nand U1992 (N_1992,N_987,N_507);
nor U1993 (N_1993,N_311,N_98);
nor U1994 (N_1994,N_369,N_439);
nor U1995 (N_1995,N_533,N_706);
nor U1996 (N_1996,N_455,N_602);
nor U1997 (N_1997,N_729,N_200);
nand U1998 (N_1998,N_527,N_419);
or U1999 (N_1999,N_251,N_765);
xor U2000 (N_2000,N_1524,N_1428);
or U2001 (N_2001,N_1075,N_1648);
xnor U2002 (N_2002,N_1223,N_1722);
nor U2003 (N_2003,N_1485,N_1758);
nor U2004 (N_2004,N_1477,N_1625);
nand U2005 (N_2005,N_1965,N_1955);
or U2006 (N_2006,N_1580,N_1816);
nand U2007 (N_2007,N_1669,N_1231);
nor U2008 (N_2008,N_1261,N_1717);
or U2009 (N_2009,N_1459,N_1576);
nand U2010 (N_2010,N_1643,N_1316);
and U2011 (N_2011,N_1448,N_1679);
or U2012 (N_2012,N_1694,N_1764);
and U2013 (N_2013,N_1315,N_1196);
xor U2014 (N_2014,N_1769,N_1107);
or U2015 (N_2015,N_1760,N_1345);
nand U2016 (N_2016,N_1569,N_1218);
nor U2017 (N_2017,N_1918,N_1403);
and U2018 (N_2018,N_1372,N_1960);
nor U2019 (N_2019,N_1347,N_1521);
nor U2020 (N_2020,N_1424,N_1386);
or U2021 (N_2021,N_1962,N_1629);
nand U2022 (N_2022,N_1836,N_1137);
nand U2023 (N_2023,N_1886,N_1048);
and U2024 (N_2024,N_1635,N_1684);
nand U2025 (N_2025,N_1865,N_1209);
nand U2026 (N_2026,N_1968,N_1890);
nor U2027 (N_2027,N_1479,N_1368);
nor U2028 (N_2028,N_1799,N_1365);
nand U2029 (N_2029,N_1084,N_1068);
nor U2030 (N_2030,N_1932,N_1011);
nor U2031 (N_2031,N_1681,N_1638);
nor U2032 (N_2032,N_1740,N_1162);
or U2033 (N_2033,N_1037,N_1619);
or U2034 (N_2034,N_1839,N_1237);
nand U2035 (N_2035,N_1626,N_1391);
nor U2036 (N_2036,N_1259,N_1299);
nor U2037 (N_2037,N_1054,N_1471);
nor U2038 (N_2038,N_1605,N_1375);
and U2039 (N_2039,N_1260,N_1108);
nand U2040 (N_2040,N_1660,N_1346);
or U2041 (N_2041,N_1041,N_1359);
nand U2042 (N_2042,N_1480,N_1438);
and U2043 (N_2043,N_1122,N_1465);
nand U2044 (N_2044,N_1138,N_1535);
and U2045 (N_2045,N_1744,N_1161);
or U2046 (N_2046,N_1541,N_1060);
or U2047 (N_2047,N_1321,N_1361);
or U2048 (N_2048,N_1667,N_1856);
and U2049 (N_2049,N_1814,N_1500);
and U2050 (N_2050,N_1227,N_1398);
nand U2051 (N_2051,N_1967,N_1492);
and U2052 (N_2052,N_1363,N_1022);
nand U2053 (N_2053,N_1826,N_1631);
nand U2054 (N_2054,N_1604,N_1240);
nand U2055 (N_2055,N_1077,N_1001);
and U2056 (N_2056,N_1936,N_1741);
nor U2057 (N_2057,N_1919,N_1730);
or U2058 (N_2058,N_1591,N_1080);
nand U2059 (N_2059,N_1297,N_1832);
and U2060 (N_2060,N_1466,N_1738);
nor U2061 (N_2061,N_1874,N_1169);
nor U2062 (N_2062,N_1731,N_1497);
nor U2063 (N_2063,N_1934,N_1053);
nand U2064 (N_2064,N_1817,N_1385);
nor U2065 (N_2065,N_1410,N_1892);
and U2066 (N_2066,N_1654,N_1776);
nor U2067 (N_2067,N_1951,N_1462);
and U2068 (N_2068,N_1376,N_1644);
nand U2069 (N_2069,N_1247,N_1748);
or U2070 (N_2070,N_1467,N_1783);
and U2071 (N_2071,N_1258,N_1241);
nor U2072 (N_2072,N_1308,N_1505);
nand U2073 (N_2073,N_1045,N_1334);
and U2074 (N_2074,N_1422,N_1763);
and U2075 (N_2075,N_1458,N_1507);
or U2076 (N_2076,N_1439,N_1300);
and U2077 (N_2077,N_1163,N_1049);
nor U2078 (N_2078,N_1494,N_1910);
nor U2079 (N_2079,N_1743,N_1303);
nand U2080 (N_2080,N_1562,N_1245);
or U2081 (N_2081,N_1533,N_1559);
and U2082 (N_2082,N_1124,N_1073);
nand U2083 (N_2083,N_1703,N_1502);
nand U2084 (N_2084,N_1343,N_1578);
and U2085 (N_2085,N_1849,N_1794);
nand U2086 (N_2086,N_1652,N_1349);
nor U2087 (N_2087,N_1023,N_1283);
nand U2088 (N_2088,N_1013,N_1174);
nor U2089 (N_2089,N_1057,N_1802);
or U2090 (N_2090,N_1618,N_1607);
and U2091 (N_2091,N_1036,N_1553);
and U2092 (N_2092,N_1104,N_1370);
nor U2093 (N_2093,N_1336,N_1145);
or U2094 (N_2094,N_1859,N_1225);
or U2095 (N_2095,N_1809,N_1118);
or U2096 (N_2096,N_1351,N_1751);
or U2097 (N_2097,N_1229,N_1517);
or U2098 (N_2098,N_1020,N_1728);
nor U2099 (N_2099,N_1242,N_1340);
nor U2100 (N_2100,N_1811,N_1292);
nor U2101 (N_2101,N_1499,N_1705);
nor U2102 (N_2102,N_1687,N_1949);
nand U2103 (N_2103,N_1094,N_1305);
or U2104 (N_2104,N_1434,N_1288);
and U2105 (N_2105,N_1083,N_1676);
nand U2106 (N_2106,N_1690,N_1989);
and U2107 (N_2107,N_1530,N_1510);
nor U2108 (N_2108,N_1573,N_1854);
or U2109 (N_2109,N_1926,N_1615);
nand U2110 (N_2110,N_1437,N_1662);
xnor U2111 (N_2111,N_1018,N_1713);
nor U2112 (N_2112,N_1254,N_1537);
nand U2113 (N_2113,N_1608,N_1423);
nor U2114 (N_2114,N_1482,N_1357);
or U2115 (N_2115,N_1866,N_1561);
and U2116 (N_2116,N_1790,N_1895);
nand U2117 (N_2117,N_1050,N_1983);
and U2118 (N_2118,N_1975,N_1944);
or U2119 (N_2119,N_1238,N_1992);
or U2120 (N_2120,N_1101,N_1824);
or U2121 (N_2121,N_1312,N_1204);
or U2122 (N_2122,N_1445,N_1613);
nor U2123 (N_2123,N_1233,N_1538);
nor U2124 (N_2124,N_1055,N_1228);
or U2125 (N_2125,N_1021,N_1767);
nor U2126 (N_2126,N_1313,N_1915);
nand U2127 (N_2127,N_1364,N_1394);
and U2128 (N_2128,N_1747,N_1270);
and U2129 (N_2129,N_1078,N_1175);
or U2130 (N_2130,N_1151,N_1838);
nand U2131 (N_2131,N_1449,N_1454);
or U2132 (N_2132,N_1444,N_1870);
or U2133 (N_2133,N_1686,N_1600);
nor U2134 (N_2134,N_1883,N_1426);
or U2135 (N_2135,N_1456,N_1503);
and U2136 (N_2136,N_1433,N_1056);
nand U2137 (N_2137,N_1765,N_1256);
or U2138 (N_2138,N_1081,N_1855);
or U2139 (N_2139,N_1211,N_1296);
nand U2140 (N_2140,N_1851,N_1215);
nand U2141 (N_2141,N_1501,N_1447);
nor U2142 (N_2142,N_1588,N_1985);
and U2143 (N_2143,N_1198,N_1806);
nor U2144 (N_2144,N_1294,N_1655);
and U2145 (N_2145,N_1033,N_1082);
nor U2146 (N_2146,N_1621,N_1155);
nand U2147 (N_2147,N_1925,N_1134);
and U2148 (N_2148,N_1401,N_1250);
nand U2149 (N_2149,N_1555,N_1478);
or U2150 (N_2150,N_1189,N_1724);
or U2151 (N_2151,N_1495,N_1773);
nor U2152 (N_2152,N_1243,N_1729);
nand U2153 (N_2153,N_1328,N_1322);
or U2154 (N_2154,N_1360,N_1484);
nand U2155 (N_2155,N_1947,N_1582);
and U2156 (N_2156,N_1476,N_1689);
and U2157 (N_2157,N_1795,N_1620);
and U2158 (N_2158,N_1788,N_1121);
nand U2159 (N_2159,N_1006,N_1413);
nand U2160 (N_2160,N_1611,N_1031);
nor U2161 (N_2161,N_1812,N_1771);
nor U2162 (N_2162,N_1852,N_1047);
or U2163 (N_2163,N_1831,N_1651);
and U2164 (N_2164,N_1143,N_1818);
and U2165 (N_2165,N_1040,N_1111);
or U2166 (N_2166,N_1381,N_1861);
nand U2167 (N_2167,N_1550,N_1072);
and U2168 (N_2168,N_1164,N_1863);
or U2169 (N_2169,N_1692,N_1335);
nand U2170 (N_2170,N_1374,N_1711);
and U2171 (N_2171,N_1441,N_1969);
nor U2172 (N_2172,N_1453,N_1583);
nor U2173 (N_2173,N_1793,N_1419);
and U2174 (N_2174,N_1131,N_1825);
nor U2175 (N_2175,N_1903,N_1027);
nand U2176 (N_2176,N_1026,N_1464);
nor U2177 (N_2177,N_1924,N_1596);
and U2178 (N_2178,N_1366,N_1805);
nor U2179 (N_2179,N_1125,N_1834);
nor U2180 (N_2180,N_1123,N_1481);
and U2181 (N_2181,N_1570,N_1135);
nand U2182 (N_2182,N_1086,N_1864);
and U2183 (N_2183,N_1871,N_1180);
nor U2184 (N_2184,N_1668,N_1509);
and U2185 (N_2185,N_1791,N_1956);
or U2186 (N_2186,N_1592,N_1688);
and U2187 (N_2187,N_1289,N_1603);
nand U2188 (N_2188,N_1102,N_1945);
or U2189 (N_2189,N_1064,N_1405);
or U2190 (N_2190,N_1429,N_1115);
nand U2191 (N_2191,N_1267,N_1496);
nand U2192 (N_2192,N_1848,N_1797);
nor U2193 (N_2193,N_1337,N_1130);
nor U2194 (N_2194,N_1837,N_1062);
nand U2195 (N_2195,N_1217,N_1264);
or U2196 (N_2196,N_1165,N_1113);
nand U2197 (N_2197,N_1966,N_1586);
and U2198 (N_2198,N_1845,N_1276);
xor U2199 (N_2199,N_1046,N_1132);
nand U2200 (N_2200,N_1443,N_1732);
nand U2201 (N_2201,N_1220,N_1158);
nand U2202 (N_2202,N_1407,N_1762);
nor U2203 (N_2203,N_1725,N_1558);
nand U2204 (N_2204,N_1133,N_1539);
or U2205 (N_2205,N_1272,N_1534);
nor U2206 (N_2206,N_1532,N_1324);
and U2207 (N_2207,N_1330,N_1599);
or U2208 (N_2208,N_1772,N_1959);
nor U2209 (N_2209,N_1787,N_1786);
or U2210 (N_2210,N_1880,N_1885);
nand U2211 (N_2211,N_1455,N_1784);
or U2212 (N_2212,N_1397,N_1602);
xnor U2213 (N_2213,N_1002,N_1896);
nor U2214 (N_2214,N_1207,N_1030);
nand U2215 (N_2215,N_1263,N_1379);
nand U2216 (N_2216,N_1986,N_1905);
or U2217 (N_2217,N_1768,N_1981);
and U2218 (N_2218,N_1007,N_1167);
and U2219 (N_2219,N_1700,N_1339);
and U2220 (N_2220,N_1702,N_1319);
nand U2221 (N_2221,N_1511,N_1636);
nand U2222 (N_2222,N_1554,N_1257);
and U2223 (N_2223,N_1807,N_1003);
or U2224 (N_2224,N_1995,N_1005);
and U2225 (N_2225,N_1286,N_1803);
nand U2226 (N_2226,N_1377,N_1043);
nor U2227 (N_2227,N_1493,N_1187);
and U2228 (N_2228,N_1463,N_1352);
and U2229 (N_2229,N_1311,N_1927);
and U2230 (N_2230,N_1513,N_1416);
and U2231 (N_2231,N_1674,N_1536);
and U2232 (N_2232,N_1156,N_1516);
nand U2233 (N_2233,N_1984,N_1693);
nor U2234 (N_2234,N_1733,N_1159);
nand U2235 (N_2235,N_1012,N_1344);
nor U2236 (N_2236,N_1815,N_1295);
nand U2237 (N_2237,N_1109,N_1899);
nor U2238 (N_2238,N_1982,N_1551);
nand U2239 (N_2239,N_1753,N_1672);
and U2240 (N_2240,N_1774,N_1819);
or U2241 (N_2241,N_1746,N_1194);
and U2242 (N_2242,N_1565,N_1285);
and U2243 (N_2243,N_1846,N_1408);
and U2244 (N_2244,N_1004,N_1875);
and U2245 (N_2245,N_1182,N_1172);
or U2246 (N_2246,N_1901,N_1110);
and U2247 (N_2247,N_1181,N_1757);
nor U2248 (N_2248,N_1879,N_1572);
nor U2249 (N_2249,N_1902,N_1504);
nor U2250 (N_2250,N_1099,N_1628);
nor U2251 (N_2251,N_1010,N_1869);
or U2252 (N_2252,N_1898,N_1318);
nor U2253 (N_2253,N_1548,N_1140);
nand U2254 (N_2254,N_1683,N_1279);
or U2255 (N_2255,N_1146,N_1273);
nor U2256 (N_2256,N_1190,N_1128);
nand U2257 (N_2257,N_1446,N_1092);
nor U2258 (N_2258,N_1239,N_1704);
or U2259 (N_2259,N_1076,N_1844);
nand U2260 (N_2260,N_1106,N_1601);
nand U2261 (N_2261,N_1673,N_1469);
nand U2262 (N_2262,N_1634,N_1939);
and U2263 (N_2263,N_1878,N_1251);
or U2264 (N_2264,N_1293,N_1906);
or U2265 (N_2265,N_1515,N_1008);
nand U2266 (N_2266,N_1800,N_1282);
and U2267 (N_2267,N_1390,N_1396);
and U2268 (N_2268,N_1953,N_1656);
nor U2269 (N_2269,N_1201,N_1275);
or U2270 (N_2270,N_1997,N_1659);
nor U2271 (N_2271,N_1320,N_1544);
nor U2272 (N_2272,N_1640,N_1540);
nor U2273 (N_2273,N_1206,N_1468);
and U2274 (N_2274,N_1088,N_1119);
and U2275 (N_2275,N_1828,N_1627);
and U2276 (N_2276,N_1853,N_1435);
nor U2277 (N_2277,N_1265,N_1563);
and U2278 (N_2278,N_1298,N_1095);
or U2279 (N_2279,N_1779,N_1042);
nor U2280 (N_2280,N_1577,N_1759);
xor U2281 (N_2281,N_1900,N_1677);
and U2282 (N_2282,N_1742,N_1508);
or U2283 (N_2283,N_1029,N_1928);
or U2284 (N_2284,N_1059,N_1362);
nor U2285 (N_2285,N_1754,N_1523);
and U2286 (N_2286,N_1105,N_1808);
nand U2287 (N_2287,N_1058,N_1149);
nor U2288 (N_2288,N_1658,N_1281);
nand U2289 (N_2289,N_1709,N_1547);
nor U2290 (N_2290,N_1192,N_1016);
and U2291 (N_2291,N_1144,N_1671);
nand U2292 (N_2292,N_1922,N_1665);
or U2293 (N_2293,N_1796,N_1150);
or U2294 (N_2294,N_1933,N_1996);
nor U2295 (N_2295,N_1065,N_1929);
nor U2296 (N_2296,N_1317,N_1527);
nor U2297 (N_2297,N_1789,N_1695);
and U2298 (N_2298,N_1531,N_1979);
xor U2299 (N_2299,N_1399,N_1798);
or U2300 (N_2300,N_1560,N_1326);
and U2301 (N_2301,N_1378,N_1205);
nand U2302 (N_2302,N_1472,N_1813);
or U2303 (N_2303,N_1197,N_1761);
or U2304 (N_2304,N_1063,N_1931);
xor U2305 (N_2305,N_1735,N_1810);
and U2306 (N_2306,N_1066,N_1830);
or U2307 (N_2307,N_1451,N_1486);
or U2308 (N_2308,N_1858,N_1384);
nor U2309 (N_2309,N_1100,N_1680);
nor U2310 (N_2310,N_1913,N_1184);
or U2311 (N_2311,N_1157,N_1999);
and U2312 (N_2312,N_1745,N_1701);
or U2313 (N_2313,N_1781,N_1622);
or U2314 (N_2314,N_1714,N_1567);
or U2315 (N_2315,N_1706,N_1718);
xnor U2316 (N_2316,N_1202,N_1338);
nand U2317 (N_2317,N_1017,N_1406);
nand U2318 (N_2318,N_1179,N_1470);
nor U2319 (N_2319,N_1208,N_1009);
and U2320 (N_2320,N_1970,N_1921);
nor U2321 (N_2321,N_1222,N_1142);
nor U2322 (N_2322,N_1766,N_1860);
nand U2323 (N_2323,N_1052,N_1061);
nand U2324 (N_2324,N_1176,N_1200);
and U2325 (N_2325,N_1327,N_1543);
or U2326 (N_2326,N_1804,N_1420);
nand U2327 (N_2327,N_1498,N_1888);
xnor U2328 (N_2328,N_1612,N_1715);
and U2329 (N_2329,N_1051,N_1290);
and U2330 (N_2330,N_1873,N_1675);
and U2331 (N_2331,N_1409,N_1226);
and U2332 (N_2332,N_1342,N_1015);
nand U2333 (N_2333,N_1964,N_1038);
or U2334 (N_2334,N_1912,N_1727);
nor U2335 (N_2335,N_1475,N_1987);
nor U2336 (N_2336,N_1801,N_1019);
nor U2337 (N_2337,N_1958,N_1483);
xnor U2338 (N_2338,N_1224,N_1302);
and U2339 (N_2339,N_1822,N_1387);
nor U2340 (N_2340,N_1721,N_1957);
or U2341 (N_2341,N_1598,N_1942);
and U2342 (N_2342,N_1884,N_1737);
nor U2343 (N_2343,N_1491,N_1271);
xor U2344 (N_2344,N_1332,N_1199);
nor U2345 (N_2345,N_1993,N_1734);
nand U2346 (N_2346,N_1545,N_1350);
nor U2347 (N_2347,N_1400,N_1230);
and U2348 (N_2348,N_1353,N_1976);
nand U2349 (N_2349,N_1606,N_1177);
nor U2350 (N_2350,N_1623,N_1193);
or U2351 (N_2351,N_1307,N_1526);
nand U2352 (N_2352,N_1367,N_1421);
nor U2353 (N_2353,N_1909,N_1708);
and U2354 (N_2354,N_1440,N_1699);
or U2355 (N_2355,N_1147,N_1395);
or U2356 (N_2356,N_1488,N_1388);
nand U2357 (N_2357,N_1840,N_1028);
or U2358 (N_2358,N_1266,N_1430);
and U2359 (N_2359,N_1542,N_1487);
and U2360 (N_2360,N_1522,N_1219);
nand U2361 (N_2361,N_1961,N_1373);
or U2362 (N_2362,N_1452,N_1000);
or U2363 (N_2363,N_1232,N_1249);
and U2364 (N_2364,N_1114,N_1436);
or U2365 (N_2365,N_1685,N_1418);
or U2366 (N_2366,N_1358,N_1647);
xor U2367 (N_2367,N_1571,N_1946);
or U2368 (N_2368,N_1633,N_1097);
or U2369 (N_2369,N_1291,N_1940);
nand U2370 (N_2370,N_1093,N_1720);
or U2371 (N_2371,N_1331,N_1032);
nand U2372 (N_2372,N_1382,N_1750);
nor U2373 (N_2373,N_1557,N_1268);
nor U2374 (N_2374,N_1564,N_1739);
nor U2375 (N_2375,N_1126,N_1262);
and U2376 (N_2376,N_1777,N_1624);
and U2377 (N_2377,N_1723,N_1988);
nor U2378 (N_2378,N_1617,N_1461);
or U2379 (N_2379,N_1014,N_1719);
nor U2380 (N_2380,N_1183,N_1841);
nand U2381 (N_2381,N_1907,N_1402);
and U2382 (N_2382,N_1248,N_1597);
and U2383 (N_2383,N_1255,N_1178);
or U2384 (N_2384,N_1314,N_1891);
or U2385 (N_2385,N_1998,N_1712);
or U2386 (N_2386,N_1820,N_1881);
nand U2387 (N_2387,N_1425,N_1978);
or U2388 (N_2388,N_1756,N_1411);
nor U2389 (N_2389,N_1380,N_1404);
and U2390 (N_2390,N_1389,N_1442);
or U2391 (N_2391,N_1707,N_1657);
nand U2392 (N_2392,N_1923,N_1914);
nand U2393 (N_2393,N_1069,N_1460);
or U2394 (N_2394,N_1857,N_1792);
nor U2395 (N_2395,N_1710,N_1512);
nor U2396 (N_2396,N_1920,N_1129);
and U2397 (N_2397,N_1637,N_1089);
and U2398 (N_2398,N_1775,N_1185);
nor U2399 (N_2399,N_1221,N_1917);
nand U2400 (N_2400,N_1614,N_1876);
and U2401 (N_2401,N_1616,N_1417);
or U2402 (N_2402,N_1642,N_1091);
nand U2403 (N_2403,N_1749,N_1235);
or U2404 (N_2404,N_1116,N_1044);
and U2405 (N_2405,N_1974,N_1490);
xnor U2406 (N_2406,N_1034,N_1590);
or U2407 (N_2407,N_1392,N_1186);
nor U2408 (N_2408,N_1348,N_1593);
nand U2409 (N_2409,N_1284,N_1904);
nand U2410 (N_2410,N_1663,N_1148);
nand U2411 (N_2411,N_1666,N_1519);
or U2412 (N_2412,N_1214,N_1549);
nor U2413 (N_2413,N_1589,N_1941);
nor U2414 (N_2414,N_1195,N_1943);
nor U2415 (N_2415,N_1244,N_1872);
nand U2416 (N_2416,N_1278,N_1584);
nand U2417 (N_2417,N_1234,N_1520);
nand U2418 (N_2418,N_1323,N_1277);
xor U2419 (N_2419,N_1782,N_1972);
nand U2420 (N_2420,N_1780,N_1246);
nor U2421 (N_2421,N_1039,N_1457);
nand U2422 (N_2422,N_1645,N_1938);
nand U2423 (N_2423,N_1641,N_1369);
or U2424 (N_2424,N_1341,N_1168);
nand U2425 (N_2425,N_1153,N_1994);
nor U2426 (N_2426,N_1894,N_1575);
and U2427 (N_2427,N_1973,N_1670);
nand U2428 (N_2428,N_1356,N_1025);
and U2429 (N_2429,N_1897,N_1170);
nor U2430 (N_2430,N_1916,N_1306);
and U2431 (N_2431,N_1574,N_1253);
and U2432 (N_2432,N_1024,N_1098);
nor U2433 (N_2433,N_1096,N_1887);
and U2434 (N_2434,N_1304,N_1074);
or U2435 (N_2435,N_1889,N_1166);
and U2436 (N_2436,N_1977,N_1212);
or U2437 (N_2437,N_1847,N_1908);
nand U2438 (N_2438,N_1835,N_1661);
and U2439 (N_2439,N_1120,N_1329);
or U2440 (N_2440,N_1450,N_1103);
or U2441 (N_2441,N_1070,N_1829);
and U2442 (N_2442,N_1649,N_1691);
nor U2443 (N_2443,N_1546,N_1154);
and U2444 (N_2444,N_1210,N_1568);
or U2445 (N_2445,N_1432,N_1843);
nand U2446 (N_2446,N_1071,N_1087);
or U2447 (N_2447,N_1867,N_1112);
or U2448 (N_2448,N_1287,N_1833);
and U2449 (N_2449,N_1139,N_1950);
or U2450 (N_2450,N_1518,N_1141);
and U2451 (N_2451,N_1393,N_1354);
or U2452 (N_2452,N_1770,N_1587);
nand U2453 (N_2453,N_1188,N_1785);
nor U2454 (N_2454,N_1333,N_1823);
nand U2455 (N_2455,N_1877,N_1595);
or U2456 (N_2456,N_1990,N_1152);
nand U2457 (N_2457,N_1609,N_1698);
and U2458 (N_2458,N_1431,N_1216);
nand U2459 (N_2459,N_1203,N_1882);
nand U2460 (N_2460,N_1821,N_1252);
nand U2461 (N_2461,N_1274,N_1954);
nor U2462 (N_2462,N_1755,N_1678);
nand U2463 (N_2463,N_1474,N_1414);
or U2464 (N_2464,N_1213,N_1269);
or U2465 (N_2465,N_1716,N_1594);
nor U2466 (N_2466,N_1415,N_1650);
and U2467 (N_2467,N_1778,N_1581);
and U2468 (N_2468,N_1991,N_1696);
nor U2469 (N_2469,N_1736,N_1646);
or U2470 (N_2470,N_1355,N_1850);
nor U2471 (N_2471,N_1325,N_1971);
nor U2472 (N_2472,N_1930,N_1085);
nand U2473 (N_2473,N_1236,N_1566);
xnor U2474 (N_2474,N_1525,N_1632);
nand U2475 (N_2475,N_1136,N_1937);
nand U2476 (N_2476,N_1529,N_1579);
or U2477 (N_2477,N_1980,N_1489);
or U2478 (N_2478,N_1090,N_1552);
nand U2479 (N_2479,N_1842,N_1952);
or U2480 (N_2480,N_1630,N_1653);
nand U2481 (N_2481,N_1427,N_1948);
or U2482 (N_2482,N_1726,N_1171);
nand U2483 (N_2483,N_1682,N_1067);
xnor U2484 (N_2484,N_1506,N_1310);
nand U2485 (N_2485,N_1117,N_1639);
nand U2486 (N_2486,N_1862,N_1585);
and U2487 (N_2487,N_1697,N_1514);
and U2488 (N_2488,N_1371,N_1191);
nand U2489 (N_2489,N_1664,N_1528);
nor U2490 (N_2490,N_1412,N_1280);
or U2491 (N_2491,N_1309,N_1383);
nand U2492 (N_2492,N_1556,N_1173);
and U2493 (N_2493,N_1301,N_1752);
nand U2494 (N_2494,N_1893,N_1827);
nand U2495 (N_2495,N_1035,N_1473);
nor U2496 (N_2496,N_1610,N_1868);
or U2497 (N_2497,N_1160,N_1911);
or U2498 (N_2498,N_1963,N_1079);
or U2499 (N_2499,N_1127,N_1935);
nor U2500 (N_2500,N_1768,N_1369);
and U2501 (N_2501,N_1549,N_1120);
and U2502 (N_2502,N_1618,N_1944);
nor U2503 (N_2503,N_1641,N_1565);
or U2504 (N_2504,N_1798,N_1018);
nor U2505 (N_2505,N_1824,N_1678);
or U2506 (N_2506,N_1018,N_1231);
nand U2507 (N_2507,N_1693,N_1803);
nand U2508 (N_2508,N_1635,N_1244);
and U2509 (N_2509,N_1824,N_1302);
or U2510 (N_2510,N_1466,N_1115);
nand U2511 (N_2511,N_1757,N_1646);
nand U2512 (N_2512,N_1870,N_1653);
or U2513 (N_2513,N_1045,N_1927);
and U2514 (N_2514,N_1462,N_1652);
or U2515 (N_2515,N_1736,N_1406);
nand U2516 (N_2516,N_1018,N_1825);
and U2517 (N_2517,N_1731,N_1050);
or U2518 (N_2518,N_1472,N_1173);
nand U2519 (N_2519,N_1752,N_1031);
or U2520 (N_2520,N_1880,N_1636);
nand U2521 (N_2521,N_1117,N_1244);
nand U2522 (N_2522,N_1520,N_1095);
nor U2523 (N_2523,N_1354,N_1905);
or U2524 (N_2524,N_1470,N_1371);
nor U2525 (N_2525,N_1330,N_1004);
nor U2526 (N_2526,N_1166,N_1410);
nand U2527 (N_2527,N_1642,N_1269);
or U2528 (N_2528,N_1522,N_1454);
nor U2529 (N_2529,N_1164,N_1495);
nor U2530 (N_2530,N_1377,N_1597);
nor U2531 (N_2531,N_1062,N_1518);
and U2532 (N_2532,N_1092,N_1931);
nand U2533 (N_2533,N_1219,N_1553);
or U2534 (N_2534,N_1088,N_1186);
nor U2535 (N_2535,N_1479,N_1634);
nor U2536 (N_2536,N_1730,N_1127);
nor U2537 (N_2537,N_1297,N_1438);
nor U2538 (N_2538,N_1587,N_1387);
nor U2539 (N_2539,N_1164,N_1959);
and U2540 (N_2540,N_1984,N_1120);
nor U2541 (N_2541,N_1131,N_1463);
and U2542 (N_2542,N_1725,N_1406);
nand U2543 (N_2543,N_1241,N_1198);
nor U2544 (N_2544,N_1377,N_1314);
nor U2545 (N_2545,N_1829,N_1763);
or U2546 (N_2546,N_1772,N_1575);
nor U2547 (N_2547,N_1713,N_1085);
or U2548 (N_2548,N_1955,N_1394);
and U2549 (N_2549,N_1620,N_1894);
nor U2550 (N_2550,N_1052,N_1194);
and U2551 (N_2551,N_1373,N_1001);
and U2552 (N_2552,N_1724,N_1772);
or U2553 (N_2553,N_1960,N_1139);
and U2554 (N_2554,N_1755,N_1717);
or U2555 (N_2555,N_1377,N_1301);
nand U2556 (N_2556,N_1543,N_1608);
nor U2557 (N_2557,N_1425,N_1617);
or U2558 (N_2558,N_1030,N_1588);
and U2559 (N_2559,N_1886,N_1422);
or U2560 (N_2560,N_1908,N_1315);
nor U2561 (N_2561,N_1441,N_1182);
or U2562 (N_2562,N_1245,N_1709);
xor U2563 (N_2563,N_1166,N_1734);
xor U2564 (N_2564,N_1455,N_1699);
or U2565 (N_2565,N_1828,N_1341);
or U2566 (N_2566,N_1560,N_1317);
or U2567 (N_2567,N_1578,N_1166);
nor U2568 (N_2568,N_1092,N_1953);
or U2569 (N_2569,N_1685,N_1501);
nand U2570 (N_2570,N_1942,N_1282);
and U2571 (N_2571,N_1946,N_1011);
or U2572 (N_2572,N_1377,N_1063);
nor U2573 (N_2573,N_1445,N_1903);
nor U2574 (N_2574,N_1246,N_1590);
nand U2575 (N_2575,N_1709,N_1057);
nand U2576 (N_2576,N_1374,N_1545);
nor U2577 (N_2577,N_1540,N_1013);
and U2578 (N_2578,N_1313,N_1316);
or U2579 (N_2579,N_1371,N_1823);
or U2580 (N_2580,N_1503,N_1188);
and U2581 (N_2581,N_1309,N_1856);
and U2582 (N_2582,N_1013,N_1853);
or U2583 (N_2583,N_1374,N_1416);
nand U2584 (N_2584,N_1118,N_1329);
and U2585 (N_2585,N_1447,N_1503);
and U2586 (N_2586,N_1367,N_1747);
or U2587 (N_2587,N_1241,N_1260);
or U2588 (N_2588,N_1979,N_1714);
and U2589 (N_2589,N_1740,N_1972);
nand U2590 (N_2590,N_1222,N_1199);
nand U2591 (N_2591,N_1400,N_1013);
nor U2592 (N_2592,N_1705,N_1628);
nor U2593 (N_2593,N_1316,N_1479);
nor U2594 (N_2594,N_1386,N_1900);
nand U2595 (N_2595,N_1346,N_1162);
nand U2596 (N_2596,N_1261,N_1487);
nor U2597 (N_2597,N_1239,N_1250);
nor U2598 (N_2598,N_1881,N_1475);
nor U2599 (N_2599,N_1510,N_1346);
or U2600 (N_2600,N_1115,N_1780);
or U2601 (N_2601,N_1331,N_1703);
xor U2602 (N_2602,N_1696,N_1174);
nor U2603 (N_2603,N_1551,N_1782);
and U2604 (N_2604,N_1773,N_1786);
or U2605 (N_2605,N_1968,N_1956);
xnor U2606 (N_2606,N_1433,N_1320);
and U2607 (N_2607,N_1032,N_1214);
nor U2608 (N_2608,N_1762,N_1142);
or U2609 (N_2609,N_1109,N_1005);
or U2610 (N_2610,N_1685,N_1740);
or U2611 (N_2611,N_1141,N_1644);
and U2612 (N_2612,N_1210,N_1771);
nand U2613 (N_2613,N_1026,N_1851);
and U2614 (N_2614,N_1793,N_1816);
or U2615 (N_2615,N_1028,N_1886);
nor U2616 (N_2616,N_1937,N_1585);
nand U2617 (N_2617,N_1764,N_1464);
nand U2618 (N_2618,N_1123,N_1302);
and U2619 (N_2619,N_1527,N_1854);
nor U2620 (N_2620,N_1274,N_1664);
or U2621 (N_2621,N_1151,N_1137);
nand U2622 (N_2622,N_1798,N_1787);
and U2623 (N_2623,N_1147,N_1578);
and U2624 (N_2624,N_1561,N_1710);
nand U2625 (N_2625,N_1105,N_1082);
nand U2626 (N_2626,N_1347,N_1314);
nand U2627 (N_2627,N_1293,N_1210);
nand U2628 (N_2628,N_1864,N_1884);
nor U2629 (N_2629,N_1943,N_1159);
nor U2630 (N_2630,N_1150,N_1403);
nor U2631 (N_2631,N_1261,N_1145);
nor U2632 (N_2632,N_1475,N_1788);
and U2633 (N_2633,N_1094,N_1349);
nor U2634 (N_2634,N_1250,N_1182);
or U2635 (N_2635,N_1311,N_1619);
and U2636 (N_2636,N_1250,N_1287);
or U2637 (N_2637,N_1018,N_1096);
or U2638 (N_2638,N_1367,N_1679);
and U2639 (N_2639,N_1456,N_1867);
nand U2640 (N_2640,N_1888,N_1081);
or U2641 (N_2641,N_1516,N_1262);
and U2642 (N_2642,N_1939,N_1292);
nor U2643 (N_2643,N_1023,N_1050);
xnor U2644 (N_2644,N_1627,N_1331);
and U2645 (N_2645,N_1376,N_1044);
or U2646 (N_2646,N_1414,N_1440);
or U2647 (N_2647,N_1935,N_1432);
nand U2648 (N_2648,N_1105,N_1582);
and U2649 (N_2649,N_1638,N_1450);
nor U2650 (N_2650,N_1888,N_1066);
and U2651 (N_2651,N_1979,N_1184);
and U2652 (N_2652,N_1413,N_1904);
nor U2653 (N_2653,N_1847,N_1950);
nand U2654 (N_2654,N_1687,N_1095);
or U2655 (N_2655,N_1446,N_1015);
and U2656 (N_2656,N_1148,N_1311);
nand U2657 (N_2657,N_1321,N_1087);
nor U2658 (N_2658,N_1065,N_1149);
nor U2659 (N_2659,N_1266,N_1316);
and U2660 (N_2660,N_1374,N_1120);
and U2661 (N_2661,N_1954,N_1464);
nor U2662 (N_2662,N_1622,N_1343);
nand U2663 (N_2663,N_1360,N_1126);
nand U2664 (N_2664,N_1339,N_1617);
and U2665 (N_2665,N_1403,N_1564);
and U2666 (N_2666,N_1840,N_1297);
nor U2667 (N_2667,N_1950,N_1111);
nor U2668 (N_2668,N_1641,N_1228);
or U2669 (N_2669,N_1232,N_1743);
nand U2670 (N_2670,N_1090,N_1061);
or U2671 (N_2671,N_1035,N_1614);
or U2672 (N_2672,N_1460,N_1026);
nor U2673 (N_2673,N_1974,N_1619);
xor U2674 (N_2674,N_1697,N_1267);
and U2675 (N_2675,N_1628,N_1466);
nand U2676 (N_2676,N_1812,N_1602);
nor U2677 (N_2677,N_1774,N_1998);
and U2678 (N_2678,N_1261,N_1984);
nor U2679 (N_2679,N_1154,N_1568);
or U2680 (N_2680,N_1265,N_1918);
or U2681 (N_2681,N_1408,N_1483);
and U2682 (N_2682,N_1426,N_1576);
and U2683 (N_2683,N_1857,N_1477);
nor U2684 (N_2684,N_1923,N_1148);
and U2685 (N_2685,N_1252,N_1428);
and U2686 (N_2686,N_1533,N_1979);
xor U2687 (N_2687,N_1576,N_1341);
nor U2688 (N_2688,N_1629,N_1344);
or U2689 (N_2689,N_1054,N_1675);
and U2690 (N_2690,N_1551,N_1346);
and U2691 (N_2691,N_1328,N_1045);
nand U2692 (N_2692,N_1086,N_1334);
nand U2693 (N_2693,N_1158,N_1967);
nor U2694 (N_2694,N_1817,N_1297);
nor U2695 (N_2695,N_1459,N_1615);
nand U2696 (N_2696,N_1253,N_1383);
and U2697 (N_2697,N_1636,N_1191);
nand U2698 (N_2698,N_1478,N_1772);
nor U2699 (N_2699,N_1095,N_1323);
nand U2700 (N_2700,N_1688,N_1845);
and U2701 (N_2701,N_1729,N_1837);
nor U2702 (N_2702,N_1259,N_1113);
or U2703 (N_2703,N_1043,N_1136);
or U2704 (N_2704,N_1683,N_1251);
nor U2705 (N_2705,N_1855,N_1966);
nor U2706 (N_2706,N_1267,N_1477);
nand U2707 (N_2707,N_1656,N_1043);
and U2708 (N_2708,N_1155,N_1727);
and U2709 (N_2709,N_1753,N_1613);
nand U2710 (N_2710,N_1599,N_1042);
nor U2711 (N_2711,N_1878,N_1529);
and U2712 (N_2712,N_1694,N_1002);
nand U2713 (N_2713,N_1647,N_1507);
and U2714 (N_2714,N_1837,N_1053);
nand U2715 (N_2715,N_1762,N_1340);
or U2716 (N_2716,N_1849,N_1612);
nor U2717 (N_2717,N_1016,N_1571);
nand U2718 (N_2718,N_1709,N_1745);
nand U2719 (N_2719,N_1974,N_1870);
nand U2720 (N_2720,N_1984,N_1461);
and U2721 (N_2721,N_1847,N_1194);
nor U2722 (N_2722,N_1790,N_1234);
and U2723 (N_2723,N_1528,N_1125);
nor U2724 (N_2724,N_1584,N_1489);
and U2725 (N_2725,N_1763,N_1069);
nand U2726 (N_2726,N_1006,N_1485);
and U2727 (N_2727,N_1772,N_1128);
or U2728 (N_2728,N_1560,N_1454);
nor U2729 (N_2729,N_1491,N_1415);
or U2730 (N_2730,N_1359,N_1702);
nand U2731 (N_2731,N_1694,N_1081);
or U2732 (N_2732,N_1055,N_1563);
nor U2733 (N_2733,N_1610,N_1747);
nand U2734 (N_2734,N_1558,N_1220);
and U2735 (N_2735,N_1719,N_1698);
nor U2736 (N_2736,N_1242,N_1483);
nand U2737 (N_2737,N_1516,N_1953);
nor U2738 (N_2738,N_1728,N_1543);
nor U2739 (N_2739,N_1158,N_1724);
nor U2740 (N_2740,N_1337,N_1945);
nand U2741 (N_2741,N_1060,N_1289);
and U2742 (N_2742,N_1617,N_1436);
nor U2743 (N_2743,N_1696,N_1049);
nor U2744 (N_2744,N_1466,N_1787);
and U2745 (N_2745,N_1716,N_1086);
or U2746 (N_2746,N_1272,N_1379);
nor U2747 (N_2747,N_1893,N_1455);
or U2748 (N_2748,N_1187,N_1617);
nor U2749 (N_2749,N_1163,N_1835);
and U2750 (N_2750,N_1104,N_1607);
or U2751 (N_2751,N_1331,N_1458);
nand U2752 (N_2752,N_1492,N_1206);
and U2753 (N_2753,N_1646,N_1829);
or U2754 (N_2754,N_1255,N_1763);
nor U2755 (N_2755,N_1136,N_1851);
or U2756 (N_2756,N_1511,N_1519);
nor U2757 (N_2757,N_1439,N_1634);
or U2758 (N_2758,N_1897,N_1732);
nand U2759 (N_2759,N_1866,N_1687);
and U2760 (N_2760,N_1856,N_1707);
nand U2761 (N_2761,N_1659,N_1968);
or U2762 (N_2762,N_1668,N_1308);
nand U2763 (N_2763,N_1821,N_1774);
nand U2764 (N_2764,N_1541,N_1197);
xor U2765 (N_2765,N_1450,N_1117);
xnor U2766 (N_2766,N_1168,N_1555);
and U2767 (N_2767,N_1189,N_1588);
nand U2768 (N_2768,N_1862,N_1509);
and U2769 (N_2769,N_1788,N_1694);
nand U2770 (N_2770,N_1544,N_1689);
or U2771 (N_2771,N_1622,N_1991);
and U2772 (N_2772,N_1602,N_1127);
nand U2773 (N_2773,N_1755,N_1170);
and U2774 (N_2774,N_1240,N_1511);
nand U2775 (N_2775,N_1859,N_1985);
nand U2776 (N_2776,N_1918,N_1365);
nor U2777 (N_2777,N_1417,N_1520);
nand U2778 (N_2778,N_1864,N_1702);
nor U2779 (N_2779,N_1041,N_1896);
and U2780 (N_2780,N_1787,N_1337);
or U2781 (N_2781,N_1510,N_1084);
and U2782 (N_2782,N_1582,N_1329);
nor U2783 (N_2783,N_1405,N_1623);
nand U2784 (N_2784,N_1569,N_1965);
and U2785 (N_2785,N_1123,N_1942);
or U2786 (N_2786,N_1879,N_1752);
and U2787 (N_2787,N_1233,N_1292);
and U2788 (N_2788,N_1619,N_1739);
and U2789 (N_2789,N_1706,N_1556);
nor U2790 (N_2790,N_1365,N_1716);
or U2791 (N_2791,N_1995,N_1025);
nor U2792 (N_2792,N_1559,N_1993);
or U2793 (N_2793,N_1928,N_1349);
nand U2794 (N_2794,N_1201,N_1710);
and U2795 (N_2795,N_1574,N_1616);
and U2796 (N_2796,N_1368,N_1344);
or U2797 (N_2797,N_1548,N_1267);
xnor U2798 (N_2798,N_1761,N_1614);
nand U2799 (N_2799,N_1394,N_1148);
and U2800 (N_2800,N_1961,N_1583);
nor U2801 (N_2801,N_1226,N_1713);
nor U2802 (N_2802,N_1148,N_1383);
nand U2803 (N_2803,N_1107,N_1613);
and U2804 (N_2804,N_1417,N_1008);
nor U2805 (N_2805,N_1897,N_1935);
and U2806 (N_2806,N_1970,N_1796);
or U2807 (N_2807,N_1529,N_1320);
or U2808 (N_2808,N_1219,N_1745);
nand U2809 (N_2809,N_1130,N_1632);
nor U2810 (N_2810,N_1909,N_1214);
and U2811 (N_2811,N_1716,N_1771);
and U2812 (N_2812,N_1220,N_1160);
nor U2813 (N_2813,N_1925,N_1547);
and U2814 (N_2814,N_1771,N_1945);
nand U2815 (N_2815,N_1143,N_1133);
and U2816 (N_2816,N_1505,N_1336);
and U2817 (N_2817,N_1206,N_1509);
xnor U2818 (N_2818,N_1665,N_1442);
nor U2819 (N_2819,N_1146,N_1221);
nand U2820 (N_2820,N_1542,N_1218);
or U2821 (N_2821,N_1483,N_1328);
or U2822 (N_2822,N_1892,N_1024);
or U2823 (N_2823,N_1639,N_1871);
nand U2824 (N_2824,N_1104,N_1999);
nor U2825 (N_2825,N_1789,N_1644);
or U2826 (N_2826,N_1116,N_1081);
xnor U2827 (N_2827,N_1366,N_1839);
nand U2828 (N_2828,N_1229,N_1545);
and U2829 (N_2829,N_1441,N_1688);
nand U2830 (N_2830,N_1196,N_1190);
and U2831 (N_2831,N_1006,N_1453);
or U2832 (N_2832,N_1780,N_1569);
nand U2833 (N_2833,N_1020,N_1417);
or U2834 (N_2834,N_1223,N_1394);
or U2835 (N_2835,N_1973,N_1301);
and U2836 (N_2836,N_1012,N_1109);
nor U2837 (N_2837,N_1292,N_1183);
and U2838 (N_2838,N_1790,N_1958);
or U2839 (N_2839,N_1152,N_1262);
and U2840 (N_2840,N_1265,N_1435);
xnor U2841 (N_2841,N_1741,N_1603);
and U2842 (N_2842,N_1121,N_1334);
and U2843 (N_2843,N_1560,N_1110);
and U2844 (N_2844,N_1302,N_1129);
and U2845 (N_2845,N_1102,N_1490);
or U2846 (N_2846,N_1641,N_1811);
or U2847 (N_2847,N_1483,N_1170);
nor U2848 (N_2848,N_1757,N_1072);
or U2849 (N_2849,N_1111,N_1604);
or U2850 (N_2850,N_1149,N_1610);
nand U2851 (N_2851,N_1308,N_1151);
nor U2852 (N_2852,N_1946,N_1671);
nor U2853 (N_2853,N_1955,N_1609);
nor U2854 (N_2854,N_1033,N_1294);
and U2855 (N_2855,N_1725,N_1872);
nor U2856 (N_2856,N_1389,N_1853);
and U2857 (N_2857,N_1018,N_1261);
or U2858 (N_2858,N_1395,N_1189);
nor U2859 (N_2859,N_1037,N_1239);
xor U2860 (N_2860,N_1153,N_1596);
or U2861 (N_2861,N_1343,N_1088);
or U2862 (N_2862,N_1183,N_1783);
and U2863 (N_2863,N_1234,N_1050);
nand U2864 (N_2864,N_1840,N_1514);
nand U2865 (N_2865,N_1338,N_1765);
or U2866 (N_2866,N_1510,N_1225);
and U2867 (N_2867,N_1878,N_1428);
and U2868 (N_2868,N_1919,N_1989);
or U2869 (N_2869,N_1982,N_1066);
and U2870 (N_2870,N_1079,N_1259);
nor U2871 (N_2871,N_1609,N_1944);
xnor U2872 (N_2872,N_1171,N_1096);
or U2873 (N_2873,N_1330,N_1768);
nor U2874 (N_2874,N_1291,N_1435);
and U2875 (N_2875,N_1748,N_1400);
nand U2876 (N_2876,N_1069,N_1624);
xor U2877 (N_2877,N_1753,N_1917);
and U2878 (N_2878,N_1315,N_1820);
and U2879 (N_2879,N_1225,N_1520);
or U2880 (N_2880,N_1813,N_1076);
nand U2881 (N_2881,N_1134,N_1898);
nand U2882 (N_2882,N_1195,N_1121);
nor U2883 (N_2883,N_1709,N_1632);
xor U2884 (N_2884,N_1725,N_1716);
nor U2885 (N_2885,N_1654,N_1074);
and U2886 (N_2886,N_1985,N_1788);
nand U2887 (N_2887,N_1897,N_1305);
nor U2888 (N_2888,N_1243,N_1692);
nor U2889 (N_2889,N_1757,N_1770);
nand U2890 (N_2890,N_1610,N_1722);
and U2891 (N_2891,N_1536,N_1262);
or U2892 (N_2892,N_1443,N_1041);
xor U2893 (N_2893,N_1949,N_1741);
and U2894 (N_2894,N_1388,N_1503);
xor U2895 (N_2895,N_1155,N_1715);
xnor U2896 (N_2896,N_1926,N_1010);
nor U2897 (N_2897,N_1131,N_1087);
and U2898 (N_2898,N_1386,N_1752);
nor U2899 (N_2899,N_1718,N_1418);
and U2900 (N_2900,N_1172,N_1112);
nand U2901 (N_2901,N_1085,N_1192);
nor U2902 (N_2902,N_1396,N_1374);
xor U2903 (N_2903,N_1938,N_1420);
or U2904 (N_2904,N_1944,N_1546);
nor U2905 (N_2905,N_1579,N_1791);
nand U2906 (N_2906,N_1692,N_1340);
nor U2907 (N_2907,N_1440,N_1321);
or U2908 (N_2908,N_1947,N_1008);
and U2909 (N_2909,N_1501,N_1703);
and U2910 (N_2910,N_1208,N_1074);
or U2911 (N_2911,N_1631,N_1832);
or U2912 (N_2912,N_1209,N_1201);
nor U2913 (N_2913,N_1603,N_1891);
or U2914 (N_2914,N_1902,N_1046);
nand U2915 (N_2915,N_1059,N_1296);
nand U2916 (N_2916,N_1913,N_1226);
nor U2917 (N_2917,N_1078,N_1152);
nor U2918 (N_2918,N_1490,N_1576);
or U2919 (N_2919,N_1457,N_1515);
nand U2920 (N_2920,N_1926,N_1114);
or U2921 (N_2921,N_1428,N_1068);
nand U2922 (N_2922,N_1589,N_1842);
xor U2923 (N_2923,N_1574,N_1056);
or U2924 (N_2924,N_1117,N_1805);
nand U2925 (N_2925,N_1124,N_1072);
nor U2926 (N_2926,N_1862,N_1617);
nand U2927 (N_2927,N_1801,N_1537);
and U2928 (N_2928,N_1148,N_1735);
nor U2929 (N_2929,N_1170,N_1271);
nand U2930 (N_2930,N_1066,N_1962);
and U2931 (N_2931,N_1480,N_1339);
nor U2932 (N_2932,N_1130,N_1496);
nor U2933 (N_2933,N_1743,N_1529);
nor U2934 (N_2934,N_1675,N_1284);
nand U2935 (N_2935,N_1934,N_1487);
nand U2936 (N_2936,N_1806,N_1974);
nor U2937 (N_2937,N_1057,N_1965);
nor U2938 (N_2938,N_1853,N_1647);
or U2939 (N_2939,N_1610,N_1621);
or U2940 (N_2940,N_1413,N_1908);
nand U2941 (N_2941,N_1662,N_1725);
or U2942 (N_2942,N_1571,N_1974);
nor U2943 (N_2943,N_1026,N_1459);
nor U2944 (N_2944,N_1814,N_1987);
or U2945 (N_2945,N_1677,N_1948);
or U2946 (N_2946,N_1819,N_1369);
or U2947 (N_2947,N_1150,N_1638);
nand U2948 (N_2948,N_1097,N_1339);
nand U2949 (N_2949,N_1090,N_1257);
nand U2950 (N_2950,N_1296,N_1958);
or U2951 (N_2951,N_1026,N_1797);
or U2952 (N_2952,N_1459,N_1239);
nor U2953 (N_2953,N_1808,N_1863);
and U2954 (N_2954,N_1305,N_1881);
nand U2955 (N_2955,N_1616,N_1132);
and U2956 (N_2956,N_1702,N_1745);
or U2957 (N_2957,N_1807,N_1085);
and U2958 (N_2958,N_1730,N_1010);
or U2959 (N_2959,N_1552,N_1246);
or U2960 (N_2960,N_1782,N_1639);
or U2961 (N_2961,N_1416,N_1038);
or U2962 (N_2962,N_1865,N_1614);
and U2963 (N_2963,N_1255,N_1044);
nand U2964 (N_2964,N_1590,N_1573);
and U2965 (N_2965,N_1953,N_1439);
nor U2966 (N_2966,N_1192,N_1264);
or U2967 (N_2967,N_1356,N_1744);
nand U2968 (N_2968,N_1550,N_1191);
and U2969 (N_2969,N_1168,N_1207);
and U2970 (N_2970,N_1655,N_1028);
and U2971 (N_2971,N_1296,N_1928);
nand U2972 (N_2972,N_1513,N_1002);
or U2973 (N_2973,N_1626,N_1725);
nand U2974 (N_2974,N_1962,N_1565);
nor U2975 (N_2975,N_1064,N_1685);
nor U2976 (N_2976,N_1924,N_1575);
and U2977 (N_2977,N_1881,N_1240);
nand U2978 (N_2978,N_1228,N_1986);
nor U2979 (N_2979,N_1097,N_1839);
and U2980 (N_2980,N_1156,N_1403);
and U2981 (N_2981,N_1125,N_1266);
nand U2982 (N_2982,N_1487,N_1016);
nand U2983 (N_2983,N_1992,N_1285);
nor U2984 (N_2984,N_1082,N_1325);
and U2985 (N_2985,N_1277,N_1935);
and U2986 (N_2986,N_1211,N_1155);
and U2987 (N_2987,N_1097,N_1391);
nand U2988 (N_2988,N_1407,N_1444);
nand U2989 (N_2989,N_1474,N_1030);
nand U2990 (N_2990,N_1487,N_1792);
and U2991 (N_2991,N_1937,N_1299);
or U2992 (N_2992,N_1870,N_1795);
nor U2993 (N_2993,N_1131,N_1629);
nand U2994 (N_2994,N_1257,N_1001);
nand U2995 (N_2995,N_1546,N_1658);
or U2996 (N_2996,N_1788,N_1206);
nor U2997 (N_2997,N_1425,N_1535);
nand U2998 (N_2998,N_1245,N_1024);
and U2999 (N_2999,N_1444,N_1278);
or U3000 (N_3000,N_2010,N_2623);
nand U3001 (N_3001,N_2272,N_2622);
and U3002 (N_3002,N_2288,N_2447);
and U3003 (N_3003,N_2459,N_2082);
nor U3004 (N_3004,N_2433,N_2872);
and U3005 (N_3005,N_2657,N_2890);
and U3006 (N_3006,N_2231,N_2265);
nand U3007 (N_3007,N_2561,N_2660);
nor U3008 (N_3008,N_2531,N_2384);
nand U3009 (N_3009,N_2391,N_2085);
and U3010 (N_3010,N_2939,N_2744);
and U3011 (N_3011,N_2119,N_2441);
nor U3012 (N_3012,N_2113,N_2118);
or U3013 (N_3013,N_2729,N_2403);
nor U3014 (N_3014,N_2855,N_2399);
nand U3015 (N_3015,N_2086,N_2696);
nor U3016 (N_3016,N_2960,N_2739);
or U3017 (N_3017,N_2785,N_2619);
nor U3018 (N_3018,N_2332,N_2347);
or U3019 (N_3019,N_2478,N_2810);
or U3020 (N_3020,N_2471,N_2873);
or U3021 (N_3021,N_2976,N_2148);
nand U3022 (N_3022,N_2781,N_2618);
or U3023 (N_3023,N_2450,N_2899);
and U3024 (N_3024,N_2383,N_2610);
nand U3025 (N_3025,N_2421,N_2259);
and U3026 (N_3026,N_2922,N_2166);
nand U3027 (N_3027,N_2732,N_2343);
and U3028 (N_3028,N_2613,N_2581);
nor U3029 (N_3029,N_2766,N_2539);
nor U3030 (N_3030,N_2263,N_2392);
nand U3031 (N_3031,N_2591,N_2200);
and U3032 (N_3032,N_2755,N_2134);
nand U3033 (N_3033,N_2205,N_2625);
or U3034 (N_3034,N_2714,N_2888);
and U3035 (N_3035,N_2730,N_2754);
and U3036 (N_3036,N_2507,N_2606);
nor U3037 (N_3037,N_2098,N_2629);
and U3038 (N_3038,N_2838,N_2595);
nor U3039 (N_3039,N_2004,N_2209);
and U3040 (N_3040,N_2814,N_2449);
and U3041 (N_3041,N_2327,N_2645);
nand U3042 (N_3042,N_2779,N_2084);
or U3043 (N_3043,N_2269,N_2175);
or U3044 (N_3044,N_2844,N_2602);
or U3045 (N_3045,N_2470,N_2163);
nand U3046 (N_3046,N_2499,N_2656);
and U3047 (N_3047,N_2527,N_2079);
nand U3048 (N_3048,N_2789,N_2135);
nor U3049 (N_3049,N_2128,N_2117);
or U3050 (N_3050,N_2364,N_2847);
and U3051 (N_3051,N_2481,N_2062);
or U3052 (N_3052,N_2544,N_2593);
nor U3053 (N_3053,N_2219,N_2199);
and U3054 (N_3054,N_2044,N_2035);
nand U3055 (N_3055,N_2815,N_2165);
nor U3056 (N_3056,N_2159,N_2257);
nand U3057 (N_3057,N_2483,N_2579);
or U3058 (N_3058,N_2260,N_2253);
and U3059 (N_3059,N_2412,N_2647);
or U3060 (N_3060,N_2115,N_2549);
nand U3061 (N_3061,N_2637,N_2167);
or U3062 (N_3062,N_2715,N_2464);
nor U3063 (N_3063,N_2140,N_2106);
nand U3064 (N_3064,N_2210,N_2051);
and U3065 (N_3065,N_2748,N_2190);
xnor U3066 (N_3066,N_2952,N_2609);
or U3067 (N_3067,N_2168,N_2104);
and U3068 (N_3068,N_2643,N_2331);
and U3069 (N_3069,N_2792,N_2676);
or U3070 (N_3070,N_2054,N_2057);
nand U3071 (N_3071,N_2768,N_2000);
or U3072 (N_3072,N_2102,N_2221);
nor U3073 (N_3073,N_2813,N_2359);
nor U3074 (N_3074,N_2979,N_2823);
or U3075 (N_3075,N_2353,N_2654);
nand U3076 (N_3076,N_2801,N_2500);
and U3077 (N_3077,N_2662,N_2493);
xnor U3078 (N_3078,N_2928,N_2162);
nor U3079 (N_3079,N_2911,N_2039);
or U3080 (N_3080,N_2719,N_2131);
and U3081 (N_3081,N_2154,N_2315);
and U3082 (N_3082,N_2338,N_2805);
or U3083 (N_3083,N_2965,N_2892);
or U3084 (N_3084,N_2711,N_2868);
or U3085 (N_3085,N_2408,N_2157);
or U3086 (N_3086,N_2372,N_2191);
and U3087 (N_3087,N_2524,N_2120);
nor U3088 (N_3088,N_2870,N_2519);
or U3089 (N_3089,N_2809,N_2393);
and U3090 (N_3090,N_2281,N_2211);
nor U3091 (N_3091,N_2405,N_2895);
and U3092 (N_3092,N_2149,N_2698);
or U3093 (N_3093,N_2664,N_2759);
or U3094 (N_3094,N_2103,N_2428);
nand U3095 (N_3095,N_2126,N_2017);
and U3096 (N_3096,N_2420,N_2280);
nand U3097 (N_3097,N_2093,N_2087);
nor U3098 (N_3098,N_2440,N_2073);
or U3099 (N_3099,N_2316,N_2632);
nor U3100 (N_3100,N_2816,N_2058);
nor U3101 (N_3101,N_2189,N_2943);
and U3102 (N_3102,N_2742,N_2097);
and U3103 (N_3103,N_2068,N_2827);
or U3104 (N_3104,N_2592,N_2217);
and U3105 (N_3105,N_2278,N_2357);
or U3106 (N_3106,N_2456,N_2641);
nand U3107 (N_3107,N_2290,N_2497);
nor U3108 (N_3108,N_2794,N_2757);
nor U3109 (N_3109,N_2961,N_2566);
nor U3110 (N_3110,N_2871,N_2516);
nor U3111 (N_3111,N_2758,N_2704);
or U3112 (N_3112,N_2036,N_2308);
or U3113 (N_3113,N_2249,N_2633);
nor U3114 (N_3114,N_2434,N_2027);
nor U3115 (N_3115,N_2917,N_2957);
nand U3116 (N_3116,N_2089,N_2514);
nand U3117 (N_3117,N_2614,N_2997);
and U3118 (N_3118,N_2038,N_2802);
nand U3119 (N_3119,N_2110,N_2448);
nand U3120 (N_3120,N_2473,N_2174);
and U3121 (N_3121,N_2684,N_2671);
or U3122 (N_3122,N_2046,N_2026);
nand U3123 (N_3123,N_2438,N_2831);
nand U3124 (N_3124,N_2621,N_2246);
or U3125 (N_3125,N_2092,N_2562);
or U3126 (N_3126,N_2548,N_2612);
or U3127 (N_3127,N_2072,N_2414);
or U3128 (N_3128,N_2993,N_2385);
nor U3129 (N_3129,N_2750,N_2243);
nand U3130 (N_3130,N_2371,N_2983);
nor U3131 (N_3131,N_2956,N_2208);
or U3132 (N_3132,N_2430,N_2193);
and U3133 (N_3133,N_2691,N_2611);
nor U3134 (N_3134,N_2410,N_2419);
or U3135 (N_3135,N_2505,N_2032);
or U3136 (N_3136,N_2161,N_2709);
nor U3137 (N_3137,N_2491,N_2821);
and U3138 (N_3138,N_2362,N_2699);
and U3139 (N_3139,N_2342,N_2649);
or U3140 (N_3140,N_2793,N_2913);
and U3141 (N_3141,N_2902,N_2651);
or U3142 (N_3142,N_2881,N_2920);
or U3143 (N_3143,N_2096,N_2713);
nand U3144 (N_3144,N_2731,N_2803);
and U3145 (N_3145,N_2452,N_2587);
nand U3146 (N_3146,N_2953,N_2176);
nor U3147 (N_3147,N_2261,N_2749);
and U3148 (N_3148,N_2417,N_2415);
nor U3149 (N_3149,N_2250,N_2294);
or U3150 (N_3150,N_2884,N_2880);
nor U3151 (N_3151,N_2553,N_2934);
nor U3152 (N_3152,N_2672,N_2791);
and U3153 (N_3153,N_2885,N_2277);
nor U3154 (N_3154,N_2747,N_2558);
nor U3155 (N_3155,N_2511,N_2689);
nor U3156 (N_3156,N_2559,N_2639);
nand U3157 (N_3157,N_2429,N_2297);
nand U3158 (N_3158,N_2404,N_2963);
and U3159 (N_3159,N_2107,N_2770);
and U3160 (N_3160,N_2454,N_2906);
and U3161 (N_3161,N_2774,N_2738);
or U3162 (N_3162,N_2045,N_2274);
nor U3163 (N_3163,N_2775,N_2160);
or U3164 (N_3164,N_2151,N_2066);
nor U3165 (N_3165,N_2653,N_2582);
and U3166 (N_3166,N_2155,N_2981);
and U3167 (N_3167,N_2427,N_2998);
nor U3168 (N_3168,N_2903,N_2285);
or U3169 (N_3169,N_2053,N_2893);
nor U3170 (N_3170,N_2508,N_2933);
nor U3171 (N_3171,N_2977,N_2318);
and U3172 (N_3172,N_2122,N_2786);
nand U3173 (N_3173,N_2145,N_2652);
nand U3174 (N_3174,N_2735,N_2503);
nand U3175 (N_3175,N_2520,N_2487);
or U3176 (N_3176,N_2179,N_2075);
or U3177 (N_3177,N_2863,N_2728);
nor U3178 (N_3178,N_2406,N_2212);
and U3179 (N_3179,N_2848,N_2631);
and U3180 (N_3180,N_2368,N_2918);
or U3181 (N_3181,N_2169,N_2170);
and U3182 (N_3182,N_2829,N_2576);
or U3183 (N_3183,N_2437,N_2279);
and U3184 (N_3184,N_2239,N_2509);
nor U3185 (N_3185,N_2330,N_2736);
or U3186 (N_3186,N_2528,N_2356);
and U3187 (N_3187,N_2047,N_2552);
nor U3188 (N_3188,N_2756,N_2289);
and U3189 (N_3189,N_2780,N_2258);
and U3190 (N_3190,N_2457,N_2948);
nand U3191 (N_3191,N_2144,N_2230);
and U3192 (N_3192,N_2186,N_2195);
nand U3193 (N_3193,N_2254,N_2530);
or U3194 (N_3194,N_2101,N_2642);
nand U3195 (N_3195,N_2008,N_2301);
and U3196 (N_3196,N_2620,N_2306);
nor U3197 (N_3197,N_2941,N_2557);
or U3198 (N_3198,N_2986,N_2206);
or U3199 (N_3199,N_2182,N_2034);
and U3200 (N_3200,N_2108,N_2143);
nand U3201 (N_3201,N_2773,N_2512);
and U3202 (N_3202,N_2705,N_2442);
and U3203 (N_3203,N_2864,N_2325);
or U3204 (N_3204,N_2019,N_2382);
nand U3205 (N_3205,N_2152,N_2266);
and U3206 (N_3206,N_2198,N_2924);
nor U3207 (N_3207,N_2575,N_2129);
nor U3208 (N_3208,N_2726,N_2894);
and U3209 (N_3209,N_2865,N_2379);
or U3210 (N_3210,N_2495,N_2146);
nor U3211 (N_3211,N_2300,N_2605);
xor U3212 (N_3212,N_2799,N_2866);
nor U3213 (N_3213,N_2255,N_2349);
and U3214 (N_3214,N_2822,N_2475);
or U3215 (N_3215,N_2589,N_2954);
and U3216 (N_3216,N_2373,N_2929);
and U3217 (N_3217,N_2227,N_2094);
nor U3218 (N_3218,N_2431,N_2076);
nand U3219 (N_3219,N_2282,N_2071);
nor U3220 (N_3220,N_2234,N_2365);
and U3221 (N_3221,N_2564,N_2955);
nand U3222 (N_3222,N_2188,N_2172);
nor U3223 (N_3223,N_2295,N_2029);
or U3224 (N_3224,N_2334,N_2240);
and U3225 (N_3225,N_2882,N_2387);
nand U3226 (N_3226,N_2667,N_2411);
or U3227 (N_3227,N_2467,N_2818);
nor U3228 (N_3228,N_2059,N_2262);
nand U3229 (N_3229,N_2970,N_2740);
and U3230 (N_3230,N_2974,N_2538);
and U3231 (N_3231,N_2237,N_2064);
or U3232 (N_3232,N_2042,N_2617);
nor U3233 (N_3233,N_2665,N_2769);
and U3234 (N_3234,N_2626,N_2795);
and U3235 (N_3235,N_2400,N_2139);
nand U3236 (N_3236,N_2533,N_2241);
and U3237 (N_3237,N_2762,N_2099);
nor U3238 (N_3238,N_2367,N_2876);
or U3239 (N_3239,N_2247,N_2028);
or U3240 (N_3240,N_2796,N_2753);
nand U3241 (N_3241,N_2883,N_2572);
nor U3242 (N_3242,N_2994,N_2291);
nor U3243 (N_3243,N_2472,N_2666);
nor U3244 (N_3244,N_2127,N_2628);
nor U3245 (N_3245,N_2225,N_2462);
or U3246 (N_3246,N_2095,N_2123);
or U3247 (N_3247,N_2350,N_2687);
nor U3248 (N_3248,N_2321,N_2307);
nor U3249 (N_3249,N_2634,N_2023);
nand U3250 (N_3250,N_2710,N_2063);
nor U3251 (N_3251,N_2150,N_2694);
or U3252 (N_3252,N_2927,N_2223);
nor U3253 (N_3253,N_2005,N_2601);
and U3254 (N_3254,N_2422,N_2109);
or U3255 (N_3255,N_2568,N_2987);
and U3256 (N_3256,N_2015,N_2771);
nor U3257 (N_3257,N_2320,N_2783);
nor U3258 (N_3258,N_2192,N_2184);
and U3259 (N_3259,N_2502,N_2078);
nand U3260 (N_3260,N_2743,N_2070);
or U3261 (N_3261,N_2337,N_2604);
xnor U3262 (N_3262,N_2366,N_2418);
nor U3263 (N_3263,N_2849,N_2389);
or U3264 (N_3264,N_2011,N_2455);
nand U3265 (N_3265,N_2837,N_2721);
and U3266 (N_3266,N_2242,N_2854);
or U3267 (N_3267,N_2940,N_2080);
nand U3268 (N_3268,N_2469,N_2302);
and U3269 (N_3269,N_2580,N_2340);
xnor U3270 (N_3270,N_2790,N_2835);
nand U3271 (N_3271,N_2286,N_2287);
nor U3272 (N_3272,N_2964,N_2658);
or U3273 (N_3273,N_2850,N_2820);
nand U3274 (N_3274,N_2485,N_2222);
nor U3275 (N_3275,N_2708,N_2048);
nor U3276 (N_3276,N_2788,N_2466);
and U3277 (N_3277,N_2886,N_2323);
or U3278 (N_3278,N_2703,N_2173);
nor U3279 (N_3279,N_2949,N_2857);
and U3280 (N_3280,N_2311,N_2583);
nand U3281 (N_3281,N_2624,N_2040);
nor U3282 (N_3282,N_2958,N_2663);
nor U3283 (N_3283,N_2930,N_2608);
and U3284 (N_3284,N_2014,N_2130);
and U3285 (N_3285,N_2482,N_2989);
or U3286 (N_3286,N_2644,N_2599);
or U3287 (N_3287,N_2317,N_2712);
or U3288 (N_3288,N_2183,N_2697);
and U3289 (N_3289,N_2985,N_2369);
nor U3290 (N_3290,N_2245,N_2980);
xor U3291 (N_3291,N_2322,N_2492);
or U3292 (N_3292,N_2007,N_2819);
and U3293 (N_3293,N_2846,N_2396);
nor U3294 (N_3294,N_2695,N_2951);
nor U3295 (N_3295,N_2778,N_2012);
and U3296 (N_3296,N_2121,N_2545);
and U3297 (N_3297,N_2006,N_2061);
nor U3298 (N_3298,N_2304,N_2377);
nand U3299 (N_3299,N_2640,N_2669);
or U3300 (N_3300,N_2830,N_2506);
nor U3301 (N_3301,N_2596,N_2706);
and U3302 (N_3302,N_2513,N_2213);
or U3303 (N_3303,N_2984,N_2378);
nand U3304 (N_3304,N_2547,N_2901);
nand U3305 (N_3305,N_2734,N_2532);
nor U3306 (N_3306,N_2180,N_2990);
nand U3307 (N_3307,N_2273,N_2767);
nand U3308 (N_3308,N_2800,N_2153);
or U3309 (N_3309,N_2563,N_2537);
nand U3310 (N_3310,N_2523,N_2238);
nor U3311 (N_3311,N_2220,N_2878);
and U3312 (N_3312,N_2555,N_2959);
nor U3313 (N_3313,N_2124,N_2588);
nand U3314 (N_3314,N_2425,N_2867);
and U3315 (N_3315,N_2171,N_2594);
nor U3316 (N_3316,N_2187,N_2394);
nor U3317 (N_3317,N_2765,N_2013);
nand U3318 (N_3318,N_2907,N_2584);
or U3319 (N_3319,N_2479,N_2312);
nor U3320 (N_3320,N_2975,N_2616);
or U3321 (N_3321,N_2016,N_2853);
or U3322 (N_3322,N_2002,N_2443);
nand U3323 (N_3323,N_2522,N_2218);
nand U3324 (N_3324,N_2201,N_2060);
nand U3325 (N_3325,N_2668,N_2484);
nand U3326 (N_3326,N_2271,N_2248);
nand U3327 (N_3327,N_2825,N_2275);
nor U3328 (N_3328,N_2679,N_2090);
or U3329 (N_3329,N_2310,N_2670);
and U3330 (N_3330,N_2486,N_2069);
nor U3331 (N_3331,N_2682,N_2091);
nand U3332 (N_3332,N_2900,N_2797);
or U3333 (N_3333,N_2116,N_2707);
or U3334 (N_3334,N_2615,N_2374);
nand U3335 (N_3335,N_2398,N_2474);
xnor U3336 (N_3336,N_2125,N_2686);
nor U3337 (N_3337,N_2501,N_2363);
or U3338 (N_3338,N_2834,N_2083);
nor U3339 (N_3339,N_2891,N_2270);
nand U3340 (N_3340,N_2158,N_2214);
or U3341 (N_3341,N_2590,N_2752);
or U3342 (N_3342,N_2808,N_2718);
and U3343 (N_3343,N_2496,N_2636);
and U3344 (N_3344,N_2515,N_2675);
nand U3345 (N_3345,N_2650,N_2760);
nor U3346 (N_3346,N_2833,N_2529);
and U3347 (N_3347,N_2946,N_2982);
nor U3348 (N_3348,N_2020,N_2388);
nor U3349 (N_3349,N_2862,N_2842);
nor U3350 (N_3350,N_2784,N_2635);
and U3351 (N_3351,N_2426,N_2973);
or U3352 (N_3352,N_2390,N_2877);
xor U3353 (N_3353,N_2723,N_2298);
and U3354 (N_3354,N_2551,N_2185);
nor U3355 (N_3355,N_2256,N_2251);
nand U3356 (N_3356,N_2879,N_2009);
nor U3357 (N_3357,N_2296,N_2041);
and U3358 (N_3358,N_2305,N_2937);
nor U3359 (N_3359,N_2380,N_2510);
and U3360 (N_3360,N_2137,N_2832);
and U3361 (N_3361,N_2971,N_2232);
or U3362 (N_3362,N_2197,N_2352);
and U3363 (N_3363,N_2646,N_2692);
nand U3364 (N_3364,N_2114,N_2319);
nor U3365 (N_3365,N_2859,N_2910);
or U3366 (N_3366,N_2578,N_2284);
nand U3367 (N_3367,N_2680,N_2346);
nor U3368 (N_3368,N_2283,N_2926);
or U3369 (N_3369,N_2550,N_2534);
and U3370 (N_3370,N_2490,N_2517);
or U3371 (N_3371,N_2567,N_2276);
and U3372 (N_3372,N_2717,N_2025);
nand U3373 (N_3373,N_2228,N_2416);
or U3374 (N_3374,N_2932,N_2055);
nand U3375 (N_3375,N_2461,N_2860);
nor U3376 (N_3376,N_2224,N_2465);
nand U3377 (N_3377,N_2498,N_2494);
and U3378 (N_3378,N_2351,N_2648);
nand U3379 (N_3379,N_2313,N_2861);
xnor U3380 (N_3380,N_2370,N_2142);
and U3381 (N_3381,N_2138,N_2683);
nor U3382 (N_3382,N_2630,N_2674);
nand U3383 (N_3383,N_2655,N_2702);
nor U3384 (N_3384,N_2056,N_2100);
nand U3385 (N_3385,N_2541,N_2701);
nor U3386 (N_3386,N_2423,N_2360);
and U3387 (N_3387,N_2194,N_2908);
nor U3388 (N_3388,N_2915,N_2972);
or U3389 (N_3389,N_2329,N_2341);
nand U3390 (N_3390,N_2081,N_2887);
nor U3391 (N_3391,N_2598,N_2571);
or U3392 (N_3392,N_2777,N_2996);
nor U3393 (N_3393,N_2141,N_2476);
and U3394 (N_3394,N_2931,N_2458);
or U3395 (N_3395,N_2968,N_2905);
nand U3396 (N_3396,N_2874,N_2573);
nor U3397 (N_3397,N_2181,N_2381);
nand U3398 (N_3398,N_2746,N_2178);
and U3399 (N_3399,N_2216,N_2597);
and U3400 (N_3400,N_2067,N_2944);
or U3401 (N_3401,N_2489,N_2435);
or U3402 (N_3402,N_2737,N_2204);
nor U3403 (N_3403,N_2309,N_2335);
nor U3404 (N_3404,N_2049,N_2022);
nor U3405 (N_3405,N_2542,N_2088);
nor U3406 (N_3406,N_2741,N_2812);
xor U3407 (N_3407,N_2999,N_2586);
nor U3408 (N_3408,N_2807,N_2386);
or U3409 (N_3409,N_2839,N_2772);
and U3410 (N_3410,N_2339,N_2824);
nand U3411 (N_3411,N_2003,N_2600);
nand U3412 (N_3412,N_2518,N_2836);
and U3413 (N_3413,N_2681,N_2546);
and U3414 (N_3414,N_2852,N_2751);
and U3415 (N_3415,N_2858,N_2397);
and U3416 (N_3416,N_2402,N_2111);
or U3417 (N_3417,N_2875,N_2348);
nor U3418 (N_3418,N_2303,N_2811);
or U3419 (N_3419,N_2226,N_2207);
or U3420 (N_3420,N_2543,N_2806);
and U3421 (N_3421,N_2413,N_2925);
or U3422 (N_3422,N_2764,N_2947);
nand U3423 (N_3423,N_2700,N_2292);
or U3424 (N_3424,N_2244,N_2525);
and U3425 (N_3425,N_2690,N_2024);
or U3426 (N_3426,N_2962,N_2988);
or U3427 (N_3427,N_2156,N_2432);
and U3428 (N_3428,N_2229,N_2074);
nand U3429 (N_3429,N_2354,N_2904);
xor U3430 (N_3430,N_2336,N_2912);
or U3431 (N_3431,N_2361,N_2897);
nand U3432 (N_3432,N_2560,N_2856);
and U3433 (N_3433,N_2202,N_2607);
or U3434 (N_3434,N_2776,N_2935);
nor U3435 (N_3435,N_2050,N_2661);
xnor U3436 (N_3436,N_2136,N_2798);
nand U3437 (N_3437,N_2898,N_2215);
nor U3438 (N_3438,N_2488,N_2031);
or U3439 (N_3439,N_2293,N_2536);
and U3440 (N_3440,N_2376,N_2978);
or U3441 (N_3441,N_2540,N_2132);
nor U3442 (N_3442,N_2203,N_2569);
nand U3443 (N_3443,N_2177,N_2919);
or U3444 (N_3444,N_2299,N_2914);
or U3445 (N_3445,N_2451,N_2233);
and U3446 (N_3446,N_2077,N_2720);
or U3447 (N_3447,N_2535,N_2724);
nand U3448 (N_3448,N_2196,N_2030);
nand U3449 (N_3449,N_2565,N_2685);
nor U3450 (N_3450,N_2577,N_2424);
nor U3451 (N_3451,N_2267,N_2043);
nor U3452 (N_3452,N_2804,N_2722);
and U3453 (N_3453,N_2328,N_2733);
nor U3454 (N_3454,N_2052,N_2936);
nor U3455 (N_3455,N_2782,N_2570);
nand U3456 (N_3456,N_2314,N_2763);
or U3457 (N_3457,N_2966,N_2401);
nor U3458 (N_3458,N_2333,N_2843);
or U3459 (N_3459,N_2727,N_2826);
nor U3460 (N_3460,N_2745,N_2869);
or U3461 (N_3461,N_2638,N_2147);
nor U3462 (N_3462,N_2678,N_2923);
xnor U3463 (N_3463,N_2112,N_2845);
nand U3464 (N_3464,N_2574,N_2252);
nor U3465 (N_3465,N_2521,N_2995);
nor U3466 (N_3466,N_2446,N_2851);
nand U3467 (N_3467,N_2018,N_2817);
and U3468 (N_3468,N_2969,N_2264);
and U3469 (N_3469,N_2673,N_2001);
or U3470 (N_3470,N_2345,N_2460);
nand U3471 (N_3471,N_2407,N_2236);
nor U3472 (N_3472,N_2344,N_2409);
and U3473 (N_3473,N_2268,N_2659);
nor U3474 (N_3474,N_2375,N_2504);
and U3475 (N_3475,N_2453,N_2326);
nand U3476 (N_3476,N_2688,N_2889);
or U3477 (N_3477,N_2942,N_2693);
or U3478 (N_3478,N_2554,N_2358);
nand U3479 (N_3479,N_2037,N_2463);
or U3480 (N_3480,N_2627,N_2105);
nand U3481 (N_3481,N_2725,N_2991);
and U3482 (N_3482,N_2585,N_2556);
nand U3483 (N_3483,N_2021,N_2945);
nand U3484 (N_3484,N_2716,N_2324);
and U3485 (N_3485,N_2896,N_2164);
nor U3486 (N_3486,N_2468,N_2841);
or U3487 (N_3487,N_2828,N_2909);
or U3488 (N_3488,N_2439,N_2921);
or U3489 (N_3489,N_2235,N_2992);
nand U3490 (N_3490,N_2444,N_2677);
nor U3491 (N_3491,N_2603,N_2477);
and U3492 (N_3492,N_2916,N_2938);
and U3493 (N_3493,N_2436,N_2967);
and U3494 (N_3494,N_2033,N_2480);
nand U3495 (N_3495,N_2133,N_2065);
nand U3496 (N_3496,N_2526,N_2840);
or U3497 (N_3497,N_2787,N_2355);
and U3498 (N_3498,N_2761,N_2395);
nor U3499 (N_3499,N_2445,N_2950);
nor U3500 (N_3500,N_2247,N_2040);
and U3501 (N_3501,N_2128,N_2512);
or U3502 (N_3502,N_2911,N_2603);
xor U3503 (N_3503,N_2621,N_2877);
nor U3504 (N_3504,N_2311,N_2088);
nor U3505 (N_3505,N_2665,N_2772);
nor U3506 (N_3506,N_2156,N_2574);
and U3507 (N_3507,N_2934,N_2810);
or U3508 (N_3508,N_2495,N_2637);
nor U3509 (N_3509,N_2171,N_2114);
or U3510 (N_3510,N_2044,N_2326);
nor U3511 (N_3511,N_2781,N_2505);
or U3512 (N_3512,N_2333,N_2144);
nand U3513 (N_3513,N_2394,N_2698);
nand U3514 (N_3514,N_2281,N_2887);
nor U3515 (N_3515,N_2904,N_2783);
nor U3516 (N_3516,N_2373,N_2925);
nor U3517 (N_3517,N_2604,N_2021);
or U3518 (N_3518,N_2474,N_2324);
and U3519 (N_3519,N_2830,N_2908);
or U3520 (N_3520,N_2713,N_2306);
nand U3521 (N_3521,N_2432,N_2453);
and U3522 (N_3522,N_2263,N_2954);
or U3523 (N_3523,N_2650,N_2143);
or U3524 (N_3524,N_2311,N_2333);
or U3525 (N_3525,N_2995,N_2780);
or U3526 (N_3526,N_2026,N_2547);
nand U3527 (N_3527,N_2874,N_2144);
or U3528 (N_3528,N_2476,N_2700);
and U3529 (N_3529,N_2127,N_2631);
and U3530 (N_3530,N_2363,N_2587);
or U3531 (N_3531,N_2131,N_2208);
and U3532 (N_3532,N_2929,N_2449);
and U3533 (N_3533,N_2226,N_2975);
or U3534 (N_3534,N_2405,N_2966);
or U3535 (N_3535,N_2553,N_2664);
nor U3536 (N_3536,N_2881,N_2299);
or U3537 (N_3537,N_2156,N_2203);
nand U3538 (N_3538,N_2474,N_2825);
nand U3539 (N_3539,N_2044,N_2150);
and U3540 (N_3540,N_2549,N_2057);
nor U3541 (N_3541,N_2122,N_2346);
or U3542 (N_3542,N_2631,N_2960);
and U3543 (N_3543,N_2789,N_2776);
nor U3544 (N_3544,N_2975,N_2372);
and U3545 (N_3545,N_2762,N_2553);
and U3546 (N_3546,N_2386,N_2273);
and U3547 (N_3547,N_2754,N_2198);
and U3548 (N_3548,N_2827,N_2586);
or U3549 (N_3549,N_2566,N_2499);
nor U3550 (N_3550,N_2323,N_2893);
nor U3551 (N_3551,N_2191,N_2928);
or U3552 (N_3552,N_2855,N_2286);
nand U3553 (N_3553,N_2522,N_2429);
or U3554 (N_3554,N_2382,N_2083);
nand U3555 (N_3555,N_2375,N_2413);
and U3556 (N_3556,N_2070,N_2397);
nor U3557 (N_3557,N_2673,N_2411);
or U3558 (N_3558,N_2690,N_2835);
and U3559 (N_3559,N_2324,N_2672);
and U3560 (N_3560,N_2206,N_2130);
and U3561 (N_3561,N_2005,N_2063);
or U3562 (N_3562,N_2130,N_2873);
and U3563 (N_3563,N_2167,N_2250);
nand U3564 (N_3564,N_2727,N_2908);
and U3565 (N_3565,N_2162,N_2187);
nor U3566 (N_3566,N_2492,N_2726);
xor U3567 (N_3567,N_2809,N_2617);
or U3568 (N_3568,N_2703,N_2993);
nand U3569 (N_3569,N_2773,N_2630);
nand U3570 (N_3570,N_2005,N_2831);
nand U3571 (N_3571,N_2097,N_2160);
nand U3572 (N_3572,N_2290,N_2787);
or U3573 (N_3573,N_2608,N_2649);
or U3574 (N_3574,N_2421,N_2638);
nand U3575 (N_3575,N_2892,N_2754);
nor U3576 (N_3576,N_2874,N_2563);
and U3577 (N_3577,N_2994,N_2945);
or U3578 (N_3578,N_2951,N_2067);
nand U3579 (N_3579,N_2816,N_2797);
nor U3580 (N_3580,N_2806,N_2630);
or U3581 (N_3581,N_2527,N_2734);
or U3582 (N_3582,N_2205,N_2473);
or U3583 (N_3583,N_2706,N_2462);
and U3584 (N_3584,N_2540,N_2151);
and U3585 (N_3585,N_2188,N_2656);
nand U3586 (N_3586,N_2128,N_2847);
nor U3587 (N_3587,N_2336,N_2712);
nand U3588 (N_3588,N_2700,N_2051);
and U3589 (N_3589,N_2161,N_2289);
or U3590 (N_3590,N_2629,N_2685);
xor U3591 (N_3591,N_2919,N_2505);
and U3592 (N_3592,N_2475,N_2814);
nand U3593 (N_3593,N_2130,N_2911);
xor U3594 (N_3594,N_2129,N_2290);
nand U3595 (N_3595,N_2729,N_2641);
nor U3596 (N_3596,N_2170,N_2916);
nand U3597 (N_3597,N_2943,N_2919);
xor U3598 (N_3598,N_2198,N_2582);
or U3599 (N_3599,N_2619,N_2729);
xor U3600 (N_3600,N_2999,N_2405);
xor U3601 (N_3601,N_2905,N_2195);
or U3602 (N_3602,N_2907,N_2695);
and U3603 (N_3603,N_2208,N_2166);
or U3604 (N_3604,N_2380,N_2978);
nand U3605 (N_3605,N_2982,N_2581);
nand U3606 (N_3606,N_2279,N_2801);
nor U3607 (N_3607,N_2817,N_2496);
nor U3608 (N_3608,N_2092,N_2862);
or U3609 (N_3609,N_2489,N_2305);
or U3610 (N_3610,N_2816,N_2076);
nor U3611 (N_3611,N_2929,N_2321);
nand U3612 (N_3612,N_2261,N_2791);
nand U3613 (N_3613,N_2677,N_2618);
nor U3614 (N_3614,N_2142,N_2374);
nand U3615 (N_3615,N_2039,N_2208);
and U3616 (N_3616,N_2520,N_2358);
or U3617 (N_3617,N_2569,N_2973);
and U3618 (N_3618,N_2786,N_2825);
nand U3619 (N_3619,N_2159,N_2997);
or U3620 (N_3620,N_2733,N_2179);
and U3621 (N_3621,N_2349,N_2835);
xnor U3622 (N_3622,N_2989,N_2533);
nor U3623 (N_3623,N_2920,N_2666);
and U3624 (N_3624,N_2521,N_2767);
and U3625 (N_3625,N_2696,N_2592);
nand U3626 (N_3626,N_2394,N_2673);
and U3627 (N_3627,N_2612,N_2839);
nand U3628 (N_3628,N_2818,N_2313);
or U3629 (N_3629,N_2079,N_2351);
nor U3630 (N_3630,N_2098,N_2592);
nand U3631 (N_3631,N_2639,N_2457);
or U3632 (N_3632,N_2254,N_2810);
or U3633 (N_3633,N_2213,N_2477);
nor U3634 (N_3634,N_2035,N_2780);
or U3635 (N_3635,N_2137,N_2239);
nor U3636 (N_3636,N_2001,N_2024);
nor U3637 (N_3637,N_2422,N_2761);
and U3638 (N_3638,N_2956,N_2993);
nand U3639 (N_3639,N_2035,N_2625);
nand U3640 (N_3640,N_2349,N_2507);
nor U3641 (N_3641,N_2322,N_2120);
nor U3642 (N_3642,N_2113,N_2680);
or U3643 (N_3643,N_2262,N_2129);
xor U3644 (N_3644,N_2729,N_2413);
nor U3645 (N_3645,N_2467,N_2494);
and U3646 (N_3646,N_2761,N_2042);
or U3647 (N_3647,N_2059,N_2424);
or U3648 (N_3648,N_2697,N_2480);
nand U3649 (N_3649,N_2830,N_2657);
nand U3650 (N_3650,N_2525,N_2774);
nor U3651 (N_3651,N_2395,N_2644);
or U3652 (N_3652,N_2326,N_2400);
or U3653 (N_3653,N_2600,N_2191);
nand U3654 (N_3654,N_2039,N_2843);
and U3655 (N_3655,N_2709,N_2604);
or U3656 (N_3656,N_2131,N_2429);
and U3657 (N_3657,N_2802,N_2235);
or U3658 (N_3658,N_2136,N_2260);
and U3659 (N_3659,N_2697,N_2119);
and U3660 (N_3660,N_2269,N_2712);
and U3661 (N_3661,N_2726,N_2644);
or U3662 (N_3662,N_2011,N_2353);
or U3663 (N_3663,N_2716,N_2759);
or U3664 (N_3664,N_2517,N_2516);
nand U3665 (N_3665,N_2728,N_2283);
and U3666 (N_3666,N_2757,N_2114);
nand U3667 (N_3667,N_2809,N_2371);
or U3668 (N_3668,N_2453,N_2876);
and U3669 (N_3669,N_2711,N_2808);
nor U3670 (N_3670,N_2259,N_2540);
and U3671 (N_3671,N_2914,N_2772);
and U3672 (N_3672,N_2112,N_2717);
or U3673 (N_3673,N_2681,N_2750);
nand U3674 (N_3674,N_2904,N_2740);
and U3675 (N_3675,N_2222,N_2724);
and U3676 (N_3676,N_2105,N_2434);
nand U3677 (N_3677,N_2944,N_2939);
or U3678 (N_3678,N_2628,N_2204);
nand U3679 (N_3679,N_2423,N_2262);
nand U3680 (N_3680,N_2326,N_2714);
or U3681 (N_3681,N_2707,N_2491);
nand U3682 (N_3682,N_2404,N_2782);
and U3683 (N_3683,N_2241,N_2330);
or U3684 (N_3684,N_2731,N_2738);
nor U3685 (N_3685,N_2566,N_2134);
nor U3686 (N_3686,N_2056,N_2838);
and U3687 (N_3687,N_2214,N_2696);
and U3688 (N_3688,N_2814,N_2296);
and U3689 (N_3689,N_2383,N_2866);
and U3690 (N_3690,N_2471,N_2934);
nand U3691 (N_3691,N_2965,N_2861);
or U3692 (N_3692,N_2703,N_2402);
or U3693 (N_3693,N_2167,N_2105);
nor U3694 (N_3694,N_2345,N_2462);
and U3695 (N_3695,N_2646,N_2021);
nor U3696 (N_3696,N_2287,N_2356);
xor U3697 (N_3697,N_2954,N_2052);
nor U3698 (N_3698,N_2545,N_2536);
nor U3699 (N_3699,N_2713,N_2883);
or U3700 (N_3700,N_2243,N_2268);
and U3701 (N_3701,N_2390,N_2049);
and U3702 (N_3702,N_2703,N_2507);
nor U3703 (N_3703,N_2426,N_2071);
nor U3704 (N_3704,N_2160,N_2042);
or U3705 (N_3705,N_2033,N_2503);
nor U3706 (N_3706,N_2798,N_2565);
nand U3707 (N_3707,N_2458,N_2659);
and U3708 (N_3708,N_2438,N_2165);
nor U3709 (N_3709,N_2688,N_2651);
nand U3710 (N_3710,N_2076,N_2365);
nand U3711 (N_3711,N_2301,N_2054);
or U3712 (N_3712,N_2819,N_2885);
or U3713 (N_3713,N_2814,N_2194);
and U3714 (N_3714,N_2401,N_2815);
nand U3715 (N_3715,N_2115,N_2044);
and U3716 (N_3716,N_2747,N_2358);
or U3717 (N_3717,N_2591,N_2954);
nor U3718 (N_3718,N_2321,N_2873);
and U3719 (N_3719,N_2095,N_2071);
nor U3720 (N_3720,N_2836,N_2150);
nor U3721 (N_3721,N_2301,N_2728);
nand U3722 (N_3722,N_2526,N_2914);
nor U3723 (N_3723,N_2729,N_2163);
nor U3724 (N_3724,N_2336,N_2532);
nand U3725 (N_3725,N_2180,N_2688);
and U3726 (N_3726,N_2328,N_2743);
nand U3727 (N_3727,N_2363,N_2644);
or U3728 (N_3728,N_2501,N_2469);
nor U3729 (N_3729,N_2042,N_2000);
and U3730 (N_3730,N_2046,N_2528);
nand U3731 (N_3731,N_2307,N_2631);
or U3732 (N_3732,N_2246,N_2639);
nand U3733 (N_3733,N_2486,N_2861);
nor U3734 (N_3734,N_2420,N_2032);
nand U3735 (N_3735,N_2535,N_2141);
xor U3736 (N_3736,N_2430,N_2673);
nor U3737 (N_3737,N_2034,N_2331);
nor U3738 (N_3738,N_2188,N_2611);
and U3739 (N_3739,N_2115,N_2129);
or U3740 (N_3740,N_2021,N_2425);
nor U3741 (N_3741,N_2334,N_2804);
or U3742 (N_3742,N_2046,N_2960);
or U3743 (N_3743,N_2549,N_2898);
nor U3744 (N_3744,N_2620,N_2895);
and U3745 (N_3745,N_2709,N_2324);
and U3746 (N_3746,N_2613,N_2679);
nor U3747 (N_3747,N_2894,N_2780);
nor U3748 (N_3748,N_2763,N_2217);
nand U3749 (N_3749,N_2925,N_2859);
and U3750 (N_3750,N_2626,N_2842);
nand U3751 (N_3751,N_2275,N_2602);
nor U3752 (N_3752,N_2484,N_2621);
nand U3753 (N_3753,N_2258,N_2720);
and U3754 (N_3754,N_2320,N_2623);
and U3755 (N_3755,N_2538,N_2623);
or U3756 (N_3756,N_2334,N_2499);
or U3757 (N_3757,N_2809,N_2785);
and U3758 (N_3758,N_2216,N_2779);
and U3759 (N_3759,N_2536,N_2119);
nand U3760 (N_3760,N_2341,N_2633);
and U3761 (N_3761,N_2361,N_2854);
or U3762 (N_3762,N_2538,N_2743);
xnor U3763 (N_3763,N_2459,N_2687);
and U3764 (N_3764,N_2504,N_2542);
nor U3765 (N_3765,N_2571,N_2936);
nand U3766 (N_3766,N_2913,N_2719);
or U3767 (N_3767,N_2116,N_2595);
nand U3768 (N_3768,N_2874,N_2322);
and U3769 (N_3769,N_2119,N_2131);
nor U3770 (N_3770,N_2946,N_2703);
or U3771 (N_3771,N_2590,N_2627);
nor U3772 (N_3772,N_2704,N_2630);
nand U3773 (N_3773,N_2360,N_2091);
or U3774 (N_3774,N_2035,N_2634);
nor U3775 (N_3775,N_2950,N_2632);
nor U3776 (N_3776,N_2430,N_2862);
and U3777 (N_3777,N_2386,N_2110);
nand U3778 (N_3778,N_2295,N_2583);
nand U3779 (N_3779,N_2859,N_2523);
nand U3780 (N_3780,N_2857,N_2191);
and U3781 (N_3781,N_2333,N_2017);
or U3782 (N_3782,N_2920,N_2089);
nor U3783 (N_3783,N_2345,N_2905);
nor U3784 (N_3784,N_2313,N_2496);
and U3785 (N_3785,N_2129,N_2440);
nor U3786 (N_3786,N_2574,N_2963);
or U3787 (N_3787,N_2618,N_2814);
or U3788 (N_3788,N_2348,N_2136);
or U3789 (N_3789,N_2260,N_2081);
and U3790 (N_3790,N_2651,N_2513);
nor U3791 (N_3791,N_2707,N_2139);
or U3792 (N_3792,N_2388,N_2850);
nand U3793 (N_3793,N_2567,N_2335);
nand U3794 (N_3794,N_2653,N_2444);
nor U3795 (N_3795,N_2079,N_2221);
or U3796 (N_3796,N_2809,N_2567);
xor U3797 (N_3797,N_2979,N_2897);
nor U3798 (N_3798,N_2064,N_2215);
or U3799 (N_3799,N_2486,N_2409);
nor U3800 (N_3800,N_2659,N_2181);
nor U3801 (N_3801,N_2290,N_2547);
xor U3802 (N_3802,N_2745,N_2352);
nand U3803 (N_3803,N_2523,N_2623);
nor U3804 (N_3804,N_2029,N_2078);
and U3805 (N_3805,N_2889,N_2551);
nor U3806 (N_3806,N_2861,N_2543);
and U3807 (N_3807,N_2239,N_2908);
and U3808 (N_3808,N_2367,N_2927);
and U3809 (N_3809,N_2767,N_2984);
nand U3810 (N_3810,N_2653,N_2390);
xor U3811 (N_3811,N_2651,N_2200);
or U3812 (N_3812,N_2661,N_2420);
and U3813 (N_3813,N_2912,N_2605);
xnor U3814 (N_3814,N_2027,N_2211);
nand U3815 (N_3815,N_2789,N_2095);
nor U3816 (N_3816,N_2744,N_2044);
or U3817 (N_3817,N_2953,N_2990);
xnor U3818 (N_3818,N_2932,N_2497);
nor U3819 (N_3819,N_2168,N_2880);
nor U3820 (N_3820,N_2235,N_2041);
and U3821 (N_3821,N_2983,N_2966);
and U3822 (N_3822,N_2059,N_2670);
and U3823 (N_3823,N_2303,N_2469);
nor U3824 (N_3824,N_2082,N_2424);
nand U3825 (N_3825,N_2363,N_2721);
nand U3826 (N_3826,N_2202,N_2445);
nand U3827 (N_3827,N_2873,N_2158);
and U3828 (N_3828,N_2621,N_2244);
nor U3829 (N_3829,N_2005,N_2585);
and U3830 (N_3830,N_2245,N_2499);
and U3831 (N_3831,N_2137,N_2085);
or U3832 (N_3832,N_2826,N_2311);
and U3833 (N_3833,N_2968,N_2936);
or U3834 (N_3834,N_2372,N_2732);
xnor U3835 (N_3835,N_2059,N_2789);
nand U3836 (N_3836,N_2194,N_2024);
nor U3837 (N_3837,N_2452,N_2563);
xor U3838 (N_3838,N_2563,N_2441);
nor U3839 (N_3839,N_2178,N_2037);
nor U3840 (N_3840,N_2424,N_2323);
and U3841 (N_3841,N_2628,N_2424);
or U3842 (N_3842,N_2766,N_2518);
and U3843 (N_3843,N_2747,N_2569);
or U3844 (N_3844,N_2942,N_2716);
nand U3845 (N_3845,N_2548,N_2300);
nor U3846 (N_3846,N_2224,N_2493);
nor U3847 (N_3847,N_2564,N_2327);
and U3848 (N_3848,N_2624,N_2053);
and U3849 (N_3849,N_2726,N_2506);
or U3850 (N_3850,N_2537,N_2454);
nor U3851 (N_3851,N_2701,N_2604);
and U3852 (N_3852,N_2347,N_2945);
and U3853 (N_3853,N_2180,N_2955);
nor U3854 (N_3854,N_2999,N_2653);
or U3855 (N_3855,N_2724,N_2677);
and U3856 (N_3856,N_2082,N_2164);
and U3857 (N_3857,N_2193,N_2771);
and U3858 (N_3858,N_2973,N_2170);
or U3859 (N_3859,N_2350,N_2865);
and U3860 (N_3860,N_2051,N_2171);
and U3861 (N_3861,N_2634,N_2321);
nor U3862 (N_3862,N_2377,N_2425);
nand U3863 (N_3863,N_2565,N_2432);
nand U3864 (N_3864,N_2093,N_2515);
nand U3865 (N_3865,N_2355,N_2804);
nand U3866 (N_3866,N_2987,N_2529);
and U3867 (N_3867,N_2766,N_2209);
or U3868 (N_3868,N_2599,N_2491);
nor U3869 (N_3869,N_2976,N_2554);
or U3870 (N_3870,N_2325,N_2896);
nand U3871 (N_3871,N_2879,N_2496);
or U3872 (N_3872,N_2611,N_2516);
and U3873 (N_3873,N_2390,N_2275);
and U3874 (N_3874,N_2238,N_2132);
or U3875 (N_3875,N_2823,N_2680);
nand U3876 (N_3876,N_2858,N_2236);
or U3877 (N_3877,N_2424,N_2592);
and U3878 (N_3878,N_2745,N_2822);
nor U3879 (N_3879,N_2565,N_2095);
nand U3880 (N_3880,N_2669,N_2042);
or U3881 (N_3881,N_2506,N_2017);
nand U3882 (N_3882,N_2596,N_2711);
or U3883 (N_3883,N_2357,N_2854);
xor U3884 (N_3884,N_2746,N_2324);
xnor U3885 (N_3885,N_2413,N_2486);
or U3886 (N_3886,N_2930,N_2798);
or U3887 (N_3887,N_2338,N_2316);
and U3888 (N_3888,N_2936,N_2552);
or U3889 (N_3889,N_2316,N_2806);
or U3890 (N_3890,N_2367,N_2278);
nor U3891 (N_3891,N_2373,N_2778);
nor U3892 (N_3892,N_2765,N_2839);
and U3893 (N_3893,N_2926,N_2944);
nand U3894 (N_3894,N_2059,N_2832);
nor U3895 (N_3895,N_2984,N_2991);
nor U3896 (N_3896,N_2753,N_2941);
or U3897 (N_3897,N_2083,N_2377);
nor U3898 (N_3898,N_2659,N_2439);
xnor U3899 (N_3899,N_2281,N_2673);
nor U3900 (N_3900,N_2473,N_2193);
nor U3901 (N_3901,N_2456,N_2174);
nand U3902 (N_3902,N_2465,N_2351);
or U3903 (N_3903,N_2893,N_2574);
or U3904 (N_3904,N_2236,N_2567);
or U3905 (N_3905,N_2545,N_2970);
nand U3906 (N_3906,N_2578,N_2076);
nor U3907 (N_3907,N_2142,N_2418);
nor U3908 (N_3908,N_2737,N_2300);
nor U3909 (N_3909,N_2587,N_2665);
nand U3910 (N_3910,N_2091,N_2168);
or U3911 (N_3911,N_2792,N_2949);
or U3912 (N_3912,N_2424,N_2316);
and U3913 (N_3913,N_2008,N_2751);
and U3914 (N_3914,N_2774,N_2885);
nand U3915 (N_3915,N_2275,N_2751);
nor U3916 (N_3916,N_2406,N_2980);
nand U3917 (N_3917,N_2171,N_2693);
nand U3918 (N_3918,N_2537,N_2634);
and U3919 (N_3919,N_2889,N_2582);
nand U3920 (N_3920,N_2351,N_2238);
or U3921 (N_3921,N_2556,N_2392);
or U3922 (N_3922,N_2988,N_2003);
nand U3923 (N_3923,N_2254,N_2615);
xor U3924 (N_3924,N_2288,N_2165);
or U3925 (N_3925,N_2942,N_2781);
nor U3926 (N_3926,N_2663,N_2397);
or U3927 (N_3927,N_2484,N_2198);
nand U3928 (N_3928,N_2103,N_2954);
and U3929 (N_3929,N_2115,N_2541);
and U3930 (N_3930,N_2651,N_2809);
nand U3931 (N_3931,N_2861,N_2911);
nor U3932 (N_3932,N_2641,N_2887);
nand U3933 (N_3933,N_2698,N_2390);
and U3934 (N_3934,N_2418,N_2623);
nand U3935 (N_3935,N_2124,N_2804);
and U3936 (N_3936,N_2204,N_2179);
or U3937 (N_3937,N_2426,N_2433);
and U3938 (N_3938,N_2537,N_2826);
nor U3939 (N_3939,N_2904,N_2383);
and U3940 (N_3940,N_2259,N_2186);
nand U3941 (N_3941,N_2687,N_2490);
nor U3942 (N_3942,N_2861,N_2502);
and U3943 (N_3943,N_2275,N_2496);
and U3944 (N_3944,N_2152,N_2718);
nor U3945 (N_3945,N_2113,N_2949);
and U3946 (N_3946,N_2932,N_2778);
or U3947 (N_3947,N_2621,N_2365);
nor U3948 (N_3948,N_2327,N_2251);
nor U3949 (N_3949,N_2713,N_2619);
nor U3950 (N_3950,N_2141,N_2851);
nor U3951 (N_3951,N_2107,N_2545);
or U3952 (N_3952,N_2994,N_2433);
nor U3953 (N_3953,N_2588,N_2438);
nor U3954 (N_3954,N_2775,N_2118);
and U3955 (N_3955,N_2163,N_2235);
or U3956 (N_3956,N_2193,N_2508);
nand U3957 (N_3957,N_2007,N_2229);
or U3958 (N_3958,N_2198,N_2354);
or U3959 (N_3959,N_2061,N_2495);
nand U3960 (N_3960,N_2535,N_2925);
and U3961 (N_3961,N_2581,N_2479);
nor U3962 (N_3962,N_2036,N_2232);
nand U3963 (N_3963,N_2570,N_2894);
and U3964 (N_3964,N_2223,N_2402);
and U3965 (N_3965,N_2444,N_2683);
or U3966 (N_3966,N_2723,N_2309);
nor U3967 (N_3967,N_2137,N_2604);
or U3968 (N_3968,N_2769,N_2176);
or U3969 (N_3969,N_2306,N_2867);
or U3970 (N_3970,N_2882,N_2057);
nor U3971 (N_3971,N_2700,N_2764);
or U3972 (N_3972,N_2438,N_2166);
nand U3973 (N_3973,N_2895,N_2245);
or U3974 (N_3974,N_2342,N_2590);
nand U3975 (N_3975,N_2211,N_2879);
nand U3976 (N_3976,N_2390,N_2145);
nor U3977 (N_3977,N_2121,N_2943);
and U3978 (N_3978,N_2108,N_2756);
and U3979 (N_3979,N_2199,N_2838);
or U3980 (N_3980,N_2013,N_2514);
nand U3981 (N_3981,N_2049,N_2359);
nor U3982 (N_3982,N_2573,N_2011);
or U3983 (N_3983,N_2816,N_2600);
nor U3984 (N_3984,N_2690,N_2989);
nor U3985 (N_3985,N_2386,N_2812);
nand U3986 (N_3986,N_2623,N_2151);
nand U3987 (N_3987,N_2207,N_2066);
nand U3988 (N_3988,N_2516,N_2393);
or U3989 (N_3989,N_2947,N_2777);
xor U3990 (N_3990,N_2699,N_2946);
or U3991 (N_3991,N_2789,N_2845);
nor U3992 (N_3992,N_2169,N_2398);
nor U3993 (N_3993,N_2778,N_2506);
xnor U3994 (N_3994,N_2550,N_2669);
nand U3995 (N_3995,N_2544,N_2152);
nand U3996 (N_3996,N_2307,N_2573);
nor U3997 (N_3997,N_2456,N_2343);
and U3998 (N_3998,N_2488,N_2419);
or U3999 (N_3999,N_2227,N_2130);
or U4000 (N_4000,N_3671,N_3007);
nor U4001 (N_4001,N_3070,N_3031);
and U4002 (N_4002,N_3491,N_3365);
nor U4003 (N_4003,N_3992,N_3417);
nor U4004 (N_4004,N_3743,N_3419);
or U4005 (N_4005,N_3896,N_3801);
nor U4006 (N_4006,N_3897,N_3162);
or U4007 (N_4007,N_3455,N_3648);
nor U4008 (N_4008,N_3503,N_3068);
nand U4009 (N_4009,N_3302,N_3326);
or U4010 (N_4010,N_3389,N_3614);
and U4011 (N_4011,N_3855,N_3608);
nor U4012 (N_4012,N_3809,N_3130);
nor U4013 (N_4013,N_3159,N_3645);
nor U4014 (N_4014,N_3144,N_3245);
or U4015 (N_4015,N_3913,N_3197);
nor U4016 (N_4016,N_3292,N_3796);
nand U4017 (N_4017,N_3836,N_3787);
nand U4018 (N_4018,N_3203,N_3370);
or U4019 (N_4019,N_3221,N_3028);
nand U4020 (N_4020,N_3841,N_3189);
and U4021 (N_4021,N_3572,N_3510);
nand U4022 (N_4022,N_3478,N_3595);
or U4023 (N_4023,N_3117,N_3766);
nand U4024 (N_4024,N_3348,N_3573);
or U4025 (N_4025,N_3006,N_3575);
or U4026 (N_4026,N_3439,N_3300);
nor U4027 (N_4027,N_3599,N_3377);
or U4028 (N_4028,N_3862,N_3630);
nor U4029 (N_4029,N_3333,N_3716);
nand U4030 (N_4030,N_3378,N_3301);
or U4031 (N_4031,N_3156,N_3810);
nand U4032 (N_4032,N_3825,N_3297);
or U4033 (N_4033,N_3066,N_3536);
nor U4034 (N_4034,N_3613,N_3314);
nand U4035 (N_4035,N_3205,N_3968);
nand U4036 (N_4036,N_3580,N_3705);
nand U4037 (N_4037,N_3084,N_3294);
nor U4038 (N_4038,N_3818,N_3228);
nor U4039 (N_4039,N_3384,N_3519);
and U4040 (N_4040,N_3547,N_3316);
and U4041 (N_4041,N_3385,N_3895);
and U4042 (N_4042,N_3103,N_3473);
and U4043 (N_4043,N_3190,N_3083);
or U4044 (N_4044,N_3606,N_3415);
nand U4045 (N_4045,N_3967,N_3753);
and U4046 (N_4046,N_3468,N_3017);
nor U4047 (N_4047,N_3647,N_3125);
and U4048 (N_4048,N_3128,N_3792);
or U4049 (N_4049,N_3701,N_3234);
and U4050 (N_4050,N_3984,N_3247);
or U4051 (N_4051,N_3578,N_3835);
and U4052 (N_4052,N_3461,N_3677);
or U4053 (N_4053,N_3436,N_3372);
nand U4054 (N_4054,N_3496,N_3443);
nand U4055 (N_4055,N_3271,N_3669);
and U4056 (N_4056,N_3770,N_3977);
nor U4057 (N_4057,N_3708,N_3155);
and U4058 (N_4058,N_3584,N_3898);
or U4059 (N_4059,N_3242,N_3783);
or U4060 (N_4060,N_3636,N_3675);
or U4061 (N_4061,N_3704,N_3448);
or U4062 (N_4062,N_3535,N_3874);
and U4063 (N_4063,N_3528,N_3408);
and U4064 (N_4064,N_3893,N_3938);
nand U4065 (N_4065,N_3941,N_3209);
nand U4066 (N_4066,N_3930,N_3298);
nor U4067 (N_4067,N_3505,N_3104);
or U4068 (N_4068,N_3587,N_3512);
or U4069 (N_4069,N_3692,N_3921);
or U4070 (N_4070,N_3576,N_3602);
nand U4071 (N_4071,N_3024,N_3808);
or U4072 (N_4072,N_3344,N_3140);
nor U4073 (N_4073,N_3023,N_3459);
nor U4074 (N_4074,N_3212,N_3986);
and U4075 (N_4075,N_3826,N_3904);
or U4076 (N_4076,N_3165,N_3313);
nand U4077 (N_4077,N_3661,N_3187);
nor U4078 (N_4078,N_3579,N_3619);
nand U4079 (N_4079,N_3356,N_3523);
and U4080 (N_4080,N_3935,N_3964);
nor U4081 (N_4081,N_3914,N_3983);
nor U4082 (N_4082,N_3269,N_3422);
nand U4083 (N_4083,N_3036,N_3252);
and U4084 (N_4084,N_3848,N_3942);
and U4085 (N_4085,N_3453,N_3413);
or U4086 (N_4086,N_3554,N_3956);
nand U4087 (N_4087,N_3639,N_3336);
and U4088 (N_4088,N_3108,N_3131);
nor U4089 (N_4089,N_3574,N_3264);
or U4090 (N_4090,N_3392,N_3851);
nand U4091 (N_4091,N_3978,N_3226);
or U4092 (N_4092,N_3831,N_3534);
nor U4093 (N_4093,N_3232,N_3526);
nand U4094 (N_4094,N_3114,N_3660);
and U4095 (N_4095,N_3172,N_3025);
or U4096 (N_4096,N_3849,N_3063);
or U4097 (N_4097,N_3041,N_3993);
and U4098 (N_4098,N_3988,N_3659);
nand U4099 (N_4099,N_3364,N_3633);
and U4100 (N_4100,N_3627,N_3488);
xor U4101 (N_4101,N_3320,N_3097);
nand U4102 (N_4102,N_3767,N_3759);
and U4103 (N_4103,N_3390,N_3664);
or U4104 (N_4104,N_3737,N_3498);
nand U4105 (N_4105,N_3532,N_3566);
or U4106 (N_4106,N_3147,N_3880);
nand U4107 (N_4107,N_3700,N_3021);
and U4108 (N_4108,N_3888,N_3092);
nand U4109 (N_4109,N_3975,N_3618);
or U4110 (N_4110,N_3736,N_3411);
nand U4111 (N_4111,N_3844,N_3065);
nor U4112 (N_4112,N_3583,N_3592);
or U4113 (N_4113,N_3431,N_3717);
nor U4114 (N_4114,N_3973,N_3728);
or U4115 (N_4115,N_3186,N_3343);
nor U4116 (N_4116,N_3892,N_3918);
or U4117 (N_4117,N_3980,N_3632);
or U4118 (N_4118,N_3662,N_3134);
nand U4119 (N_4119,N_3658,N_3082);
nor U4120 (N_4120,N_3873,N_3557);
nor U4121 (N_4121,N_3426,N_3291);
and U4122 (N_4122,N_3043,N_3279);
nand U4123 (N_4123,N_3544,N_3217);
or U4124 (N_4124,N_3119,N_3734);
nand U4125 (N_4125,N_3255,N_3460);
nand U4126 (N_4126,N_3502,N_3901);
or U4127 (N_4127,N_3121,N_3571);
or U4128 (N_4128,N_3037,N_3740);
nor U4129 (N_4129,N_3141,N_3257);
or U4130 (N_4130,N_3014,N_3427);
or U4131 (N_4131,N_3802,N_3093);
or U4132 (N_4132,N_3253,N_3804);
and U4133 (N_4133,N_3244,N_3341);
nor U4134 (N_4134,N_3946,N_3886);
and U4135 (N_4135,N_3620,N_3054);
nand U4136 (N_4136,N_3278,N_3754);
or U4137 (N_4137,N_3714,N_3756);
or U4138 (N_4138,N_3761,N_3843);
or U4139 (N_4139,N_3860,N_3883);
nor U4140 (N_4140,N_3338,N_3868);
or U4141 (N_4141,N_3444,N_3075);
and U4142 (N_4142,N_3456,N_3713);
nor U4143 (N_4143,N_3755,N_3570);
nand U4144 (N_4144,N_3838,N_3237);
nor U4145 (N_4145,N_3793,N_3170);
or U4146 (N_4146,N_3072,N_3040);
nand U4147 (N_4147,N_3612,N_3044);
or U4148 (N_4148,N_3865,N_3123);
or U4149 (N_4149,N_3605,N_3936);
or U4150 (N_4150,N_3911,N_3230);
nor U4151 (N_4151,N_3497,N_3350);
or U4152 (N_4152,N_3702,N_3349);
nand U4153 (N_4153,N_3568,N_3591);
nor U4154 (N_4154,N_3721,N_3567);
nand U4155 (N_4155,N_3288,N_3745);
and U4156 (N_4156,N_3687,N_3481);
or U4157 (N_4157,N_3691,N_3120);
or U4158 (N_4158,N_3345,N_3013);
and U4159 (N_4159,N_3863,N_3805);
and U4160 (N_4160,N_3061,N_3136);
xnor U4161 (N_4161,N_3323,N_3876);
nor U4162 (N_4162,N_3507,N_3052);
and U4163 (N_4163,N_3394,N_3916);
nor U4164 (N_4164,N_3951,N_3931);
and U4165 (N_4165,N_3823,N_3680);
nor U4166 (N_4166,N_3397,N_3582);
nand U4167 (N_4167,N_3981,N_3788);
nor U4168 (N_4168,N_3005,N_3404);
nor U4169 (N_4169,N_3012,N_3877);
nor U4170 (N_4170,N_3772,N_3723);
and U4171 (N_4171,N_3915,N_3281);
nor U4172 (N_4172,N_3903,N_3414);
nand U4173 (N_4173,N_3601,N_3208);
nand U4174 (N_4174,N_3145,N_3233);
nand U4175 (N_4175,N_3227,N_3666);
nor U4176 (N_4176,N_3046,N_3961);
or U4177 (N_4177,N_3039,N_3373);
or U4178 (N_4178,N_3520,N_3943);
nand U4179 (N_4179,N_3195,N_3077);
and U4180 (N_4180,N_3790,N_3261);
or U4181 (N_4181,N_3667,N_3907);
or U4182 (N_4182,N_3985,N_3506);
and U4183 (N_4183,N_3295,N_3029);
nand U4184 (N_4184,N_3132,N_3543);
nor U4185 (N_4185,N_3749,N_3925);
nor U4186 (N_4186,N_3138,N_3254);
nand U4187 (N_4187,N_3192,N_3989);
nor U4188 (N_4188,N_3421,N_3246);
nand U4189 (N_4189,N_3188,N_3990);
nand U4190 (N_4190,N_3486,N_3797);
or U4191 (N_4191,N_3183,N_3803);
nor U4192 (N_4192,N_3194,N_3908);
nand U4193 (N_4193,N_3330,N_3479);
nand U4194 (N_4194,N_3173,N_3214);
or U4195 (N_4195,N_3565,N_3598);
nor U4196 (N_4196,N_3080,N_3465);
or U4197 (N_4197,N_3731,N_3504);
and U4198 (N_4198,N_3861,N_3449);
and U4199 (N_4199,N_3629,N_3588);
nor U4200 (N_4200,N_3485,N_3199);
and U4201 (N_4201,N_3056,N_3672);
nand U4202 (N_4202,N_3905,N_3391);
nor U4203 (N_4203,N_3290,N_3213);
xor U4204 (N_4204,N_3018,N_3937);
and U4205 (N_4205,N_3732,N_3940);
and U4206 (N_4206,N_3603,N_3850);
nor U4207 (N_4207,N_3429,N_3376);
and U4208 (N_4208,N_3387,N_3076);
nor U4209 (N_4209,N_3000,N_3765);
nor U4210 (N_4210,N_3684,N_3073);
or U4211 (N_4211,N_3435,N_3610);
nor U4212 (N_4212,N_3438,N_3762);
or U4213 (N_4213,N_3078,N_3537);
and U4214 (N_4214,N_3824,N_3727);
nor U4215 (N_4215,N_3361,N_3777);
and U4216 (N_4216,N_3926,N_3178);
nand U4217 (N_4217,N_3858,N_3229);
nor U4218 (N_4218,N_3109,N_3501);
or U4219 (N_4219,N_3773,N_3064);
and U4220 (N_4220,N_3798,N_3270);
nor U4221 (N_4221,N_3871,N_3428);
nand U4222 (N_4222,N_3353,N_3458);
nor U4223 (N_4223,N_3321,N_3222);
nand U4224 (N_4224,N_3464,N_3176);
nand U4225 (N_4225,N_3154,N_3581);
or U4226 (N_4226,N_3492,N_3358);
nand U4227 (N_4227,N_3335,N_3655);
nand U4228 (N_4228,N_3181,N_3932);
nand U4229 (N_4229,N_3955,N_3126);
and U4230 (N_4230,N_3681,N_3106);
nor U4231 (N_4231,N_3626,N_3347);
or U4232 (N_4232,N_3719,N_3371);
nor U4233 (N_4233,N_3157,N_3207);
and U4234 (N_4234,N_3319,N_3407);
and U4235 (N_4235,N_3410,N_3726);
nor U4236 (N_4236,N_3034,N_3164);
nand U4237 (N_4237,N_3569,N_3529);
or U4238 (N_4238,N_3033,N_3463);
nor U4239 (N_4239,N_3718,N_3474);
nor U4240 (N_4240,N_3062,N_3081);
nor U4241 (N_4241,N_3098,N_3337);
and U4242 (N_4242,N_3275,N_3634);
or U4243 (N_4243,N_3146,N_3499);
or U4244 (N_4244,N_3651,N_3440);
and U4245 (N_4245,N_3418,N_3885);
nand U4246 (N_4246,N_3631,N_3711);
or U4247 (N_4247,N_3396,N_3894);
or U4248 (N_4248,N_3558,N_3060);
nor U4249 (N_4249,N_3971,N_3842);
nand U4250 (N_4250,N_3267,N_3225);
or U4251 (N_4251,N_3697,N_3806);
or U4252 (N_4252,N_3346,N_3739);
nand U4253 (N_4253,N_3948,N_3712);
or U4254 (N_4254,N_3003,N_3864);
and U4255 (N_4255,N_3306,N_3779);
or U4256 (N_4256,N_3022,N_3322);
nor U4257 (N_4257,N_3210,N_3287);
nand U4258 (N_4258,N_3293,N_3774);
or U4259 (N_4259,N_3265,N_3696);
or U4260 (N_4260,N_3059,N_3383);
and U4261 (N_4261,N_3266,N_3462);
or U4262 (N_4262,N_3891,N_3887);
and U4263 (N_4263,N_3611,N_3169);
nand U4264 (N_4264,N_3500,N_3457);
and U4265 (N_4265,N_3161,N_3251);
or U4266 (N_4266,N_3331,N_3870);
or U4267 (N_4267,N_3202,N_3091);
and U4268 (N_4268,N_3924,N_3540);
or U4269 (N_4269,N_3920,N_3048);
nor U4270 (N_4270,N_3476,N_3508);
or U4271 (N_4271,N_3483,N_3211);
nand U4272 (N_4272,N_3733,N_3878);
nor U4273 (N_4273,N_3339,N_3859);
or U4274 (N_4274,N_3374,N_3546);
nor U4275 (N_4275,N_3781,N_3089);
nor U4276 (N_4276,N_3263,N_3654);
nand U4277 (N_4277,N_3906,N_3856);
nor U4278 (N_4278,N_3118,N_3193);
or U4279 (N_4279,N_3405,N_3152);
nand U4280 (N_4280,N_3996,N_3305);
nand U4281 (N_4281,N_3142,N_3074);
or U4282 (N_4282,N_3609,N_3088);
nand U4283 (N_4283,N_3315,N_3682);
nand U4284 (N_4284,N_3057,N_3853);
nand U4285 (N_4285,N_3177,N_3239);
nor U4286 (N_4286,N_3747,N_3368);
nor U4287 (N_4287,N_3454,N_3148);
nor U4288 (N_4288,N_3451,N_3615);
nand U4289 (N_4289,N_3515,N_3852);
or U4290 (N_4290,N_3067,N_3800);
and U4291 (N_4291,N_3812,N_3289);
nor U4292 (N_4292,N_3775,N_3351);
or U4293 (N_4293,N_3703,N_3381);
or U4294 (N_4294,N_3725,N_3004);
nor U4295 (N_4295,N_3312,N_3122);
nand U4296 (N_4296,N_3815,N_3690);
nand U4297 (N_4297,N_3215,N_3099);
or U4298 (N_4298,N_3129,N_3741);
nand U4299 (N_4299,N_3757,N_3471);
nand U4300 (N_4300,N_3527,N_3730);
and U4301 (N_4301,N_3934,N_3828);
or U4302 (N_4302,N_3751,N_3735);
nand U4303 (N_4303,N_3693,N_3890);
or U4304 (N_4304,N_3845,N_3958);
and U4305 (N_4305,N_3469,N_3524);
and U4306 (N_4306,N_3668,N_3259);
and U4307 (N_4307,N_3676,N_3991);
nand U4308 (N_4308,N_3038,N_3273);
nor U4309 (N_4309,N_3685,N_3447);
and U4310 (N_4310,N_3564,N_3517);
nand U4311 (N_4311,N_3811,N_3280);
nand U4312 (N_4312,N_3002,N_3722);
and U4313 (N_4313,N_3284,N_3837);
or U4314 (N_4314,N_3160,N_3107);
nand U4315 (N_4315,N_3477,N_3947);
and U4316 (N_4316,N_3830,N_3560);
and U4317 (N_4317,N_3869,N_3105);
and U4318 (N_4318,N_3495,N_3521);
xor U4319 (N_4319,N_3635,N_3650);
and U4320 (N_4320,N_3102,N_3933);
and U4321 (N_4321,N_3113,N_3998);
and U4322 (N_4322,N_3450,N_3555);
nand U4323 (N_4323,N_3917,N_3966);
and U4324 (N_4324,N_3694,N_3406);
nand U4325 (N_4325,N_3559,N_3051);
or U4326 (N_4326,N_3541,N_3218);
nor U4327 (N_4327,N_3324,N_3729);
nor U4328 (N_4328,N_3982,N_3785);
nand U4329 (N_4329,N_3533,N_3184);
nand U4330 (N_4330,N_3179,N_3027);
nor U4331 (N_4331,N_3309,N_3231);
and U4332 (N_4332,N_3604,N_3282);
nor U4333 (N_4333,N_3709,N_3786);
and U4334 (N_4334,N_3764,N_3832);
and U4335 (N_4335,N_3328,N_3401);
or U4336 (N_4336,N_3020,N_3437);
or U4337 (N_4337,N_3516,N_3166);
nand U4338 (N_4338,N_3311,N_3545);
and U4339 (N_4339,N_3642,N_3769);
and U4340 (N_4340,N_3442,N_3472);
nand U4341 (N_4341,N_3673,N_3791);
nand U4342 (N_4342,N_3268,N_3032);
nand U4343 (N_4343,N_3399,N_3807);
nor U4344 (N_4344,N_3285,N_3402);
nand U4345 (N_4345,N_3386,N_3875);
and U4346 (N_4346,N_3359,N_3699);
nor U4347 (N_4347,N_3274,N_3008);
and U4348 (N_4348,N_3551,N_3416);
or U4349 (N_4349,N_3970,N_3596);
and U4350 (N_4350,N_3960,N_3763);
and U4351 (N_4351,N_3276,N_3016);
nand U4352 (N_4352,N_3683,N_3191);
nor U4353 (N_4353,N_3015,N_3949);
and U4354 (N_4354,N_3182,N_3899);
or U4355 (N_4355,N_3889,N_3799);
or U4356 (N_4356,N_3997,N_3538);
nor U4357 (N_4357,N_3927,N_3133);
nor U4358 (N_4358,N_3518,N_3782);
and U4359 (N_4359,N_3678,N_3665);
nor U4360 (N_4360,N_3026,N_3771);
nor U4361 (N_4361,N_3670,N_3393);
or U4362 (N_4362,N_3738,N_3623);
nand U4363 (N_4363,N_3094,N_3085);
and U4364 (N_4364,N_3480,N_3553);
or U4365 (N_4365,N_3640,N_3995);
nor U4366 (N_4366,N_3151,N_3047);
and U4367 (N_4367,N_3470,N_3742);
or U4368 (N_4368,N_3340,N_3299);
or U4369 (N_4369,N_3352,N_3168);
or U4370 (N_4370,N_3248,N_3467);
nand U4371 (N_4371,N_3962,N_3952);
or U4372 (N_4372,N_3434,N_3784);
nand U4373 (N_4373,N_3550,N_3303);
and U4374 (N_4374,N_3403,N_3332);
and U4375 (N_4375,N_3432,N_3748);
or U4376 (N_4376,N_3380,N_3216);
and U4377 (N_4377,N_3577,N_3674);
nor U4378 (N_4378,N_3260,N_3482);
nor U4379 (N_4379,N_3135,N_3220);
nand U4380 (N_4380,N_3957,N_3624);
and U4381 (N_4381,N_3539,N_3600);
xnor U4382 (N_4382,N_3819,N_3689);
nand U4383 (N_4383,N_3042,N_3101);
nor U4384 (N_4384,N_3446,N_3055);
and U4385 (N_4385,N_3643,N_3362);
and U4386 (N_4386,N_3760,N_3881);
nand U4387 (N_4387,N_3272,N_3433);
or U4388 (N_4388,N_3308,N_3929);
or U4389 (N_4389,N_3820,N_3912);
nor U4390 (N_4390,N_3706,N_3780);
xor U4391 (N_4391,N_3834,N_3549);
and U4392 (N_4392,N_3744,N_3010);
nand U4393 (N_4393,N_3637,N_3698);
nand U4394 (N_4394,N_3310,N_3096);
or U4395 (N_4395,N_3663,N_3750);
or U4396 (N_4396,N_3652,N_3412);
or U4397 (N_4397,N_3866,N_3695);
nand U4398 (N_4398,N_3079,N_3525);
nand U4399 (N_4399,N_3342,N_3827);
and U4400 (N_4400,N_3707,N_3965);
and U4401 (N_4401,N_3616,N_3163);
or U4402 (N_4402,N_3939,N_3425);
or U4403 (N_4403,N_3180,N_3286);
nand U4404 (N_4404,N_3867,N_3902);
or U4405 (N_4405,N_3149,N_3656);
and U4406 (N_4406,N_3009,N_3531);
or U4407 (N_4407,N_3019,N_3355);
nor U4408 (N_4408,N_3715,N_3087);
and U4409 (N_4409,N_3127,N_3090);
or U4410 (N_4410,N_3768,N_3489);
nand U4411 (N_4411,N_3882,N_3833);
and U4412 (N_4412,N_3919,N_3334);
nor U4413 (N_4413,N_3593,N_3112);
or U4414 (N_4414,N_3369,N_3175);
and U4415 (N_4415,N_3283,N_3950);
or U4416 (N_4416,N_3258,N_3277);
or U4417 (N_4417,N_3243,N_3360);
and U4418 (N_4418,N_3969,N_3240);
nor U4419 (N_4419,N_3910,N_3822);
nand U4420 (N_4420,N_3445,N_3909);
or U4421 (N_4421,N_3110,N_3649);
nor U4422 (N_4422,N_3999,N_3095);
or U4423 (N_4423,N_3688,N_3398);
nor U4424 (N_4424,N_3409,N_3111);
nand U4425 (N_4425,N_3625,N_3653);
or U4426 (N_4426,N_3366,N_3974);
and U4427 (N_4427,N_3900,N_3236);
and U4428 (N_4428,N_3847,N_3423);
nand U4429 (N_4429,N_3686,N_3475);
and U4430 (N_4430,N_3318,N_3628);
nand U4431 (N_4431,N_3622,N_3420);
nand U4432 (N_4432,N_3585,N_3879);
nor U4433 (N_4433,N_3382,N_3752);
and U4434 (N_4434,N_3388,N_3049);
or U4435 (N_4435,N_3794,N_3976);
nor U4436 (N_4436,N_3814,N_3710);
or U4437 (N_4437,N_3185,N_3354);
nand U4438 (N_4438,N_3100,N_3171);
nor U4439 (N_4439,N_3200,N_3466);
nand U4440 (N_4440,N_3137,N_3307);
nor U4441 (N_4441,N_3363,N_3045);
and U4442 (N_4442,N_3400,N_3329);
or U4443 (N_4443,N_3124,N_3795);
or U4444 (N_4444,N_3201,N_3679);
nand U4445 (N_4445,N_3789,N_3972);
xor U4446 (N_4446,N_3452,N_3235);
nor U4447 (N_4447,N_3561,N_3238);
or U4448 (N_4448,N_3327,N_3589);
nand U4449 (N_4449,N_3249,N_3562);
or U4450 (N_4450,N_3963,N_3953);
and U4451 (N_4451,N_3494,N_3641);
nor U4452 (N_4452,N_3646,N_3241);
nor U4453 (N_4453,N_3430,N_3617);
nor U4454 (N_4454,N_3821,N_3839);
or U4455 (N_4455,N_3817,N_3198);
or U4456 (N_4456,N_3840,N_3001);
or U4457 (N_4457,N_3857,N_3053);
xor U4458 (N_4458,N_3011,N_3071);
nand U4459 (N_4459,N_3317,N_3050);
nand U4460 (N_4460,N_3778,N_3223);
or U4461 (N_4461,N_3219,N_3514);
nor U4462 (N_4462,N_3923,N_3987);
or U4463 (N_4463,N_3484,N_3367);
and U4464 (N_4464,N_3493,N_3979);
or U4465 (N_4465,N_3621,N_3139);
nor U4466 (N_4466,N_3143,N_3776);
or U4467 (N_4467,N_3994,N_3954);
nor U4468 (N_4468,N_3959,N_3296);
nand U4469 (N_4469,N_3375,N_3115);
or U4470 (N_4470,N_3250,N_3158);
nand U4471 (N_4471,N_3490,N_3206);
nand U4472 (N_4472,N_3196,N_3086);
xnor U4473 (N_4473,N_3552,N_3816);
or U4474 (N_4474,N_3720,N_3542);
nor U4475 (N_4475,N_3607,N_3509);
or U4476 (N_4476,N_3597,N_3116);
nor U4477 (N_4477,N_3325,N_3644);
nand U4478 (N_4478,N_3922,N_3657);
or U4479 (N_4479,N_3556,N_3513);
or U4480 (N_4480,N_3357,N_3204);
nor U4481 (N_4481,N_3846,N_3522);
nor U4482 (N_4482,N_3424,N_3586);
and U4483 (N_4483,N_3872,N_3746);
nand U4484 (N_4484,N_3884,N_3548);
and U4485 (N_4485,N_3829,N_3638);
nand U4486 (N_4486,N_3945,N_3441);
or U4487 (N_4487,N_3854,N_3594);
nand U4488 (N_4488,N_3224,N_3035);
and U4489 (N_4489,N_3256,N_3379);
nor U4490 (N_4490,N_3395,N_3563);
and U4491 (N_4491,N_3150,N_3758);
and U4492 (N_4492,N_3590,N_3174);
and U4493 (N_4493,N_3030,N_3944);
or U4494 (N_4494,N_3153,N_3487);
nand U4495 (N_4495,N_3511,N_3304);
nor U4496 (N_4496,N_3167,N_3724);
or U4497 (N_4497,N_3530,N_3058);
nand U4498 (N_4498,N_3069,N_3813);
nand U4499 (N_4499,N_3928,N_3262);
xnor U4500 (N_4500,N_3217,N_3919);
nand U4501 (N_4501,N_3641,N_3897);
nand U4502 (N_4502,N_3900,N_3858);
nand U4503 (N_4503,N_3747,N_3212);
nor U4504 (N_4504,N_3106,N_3793);
xnor U4505 (N_4505,N_3609,N_3766);
nand U4506 (N_4506,N_3395,N_3425);
nand U4507 (N_4507,N_3587,N_3468);
nand U4508 (N_4508,N_3829,N_3025);
and U4509 (N_4509,N_3345,N_3870);
nand U4510 (N_4510,N_3043,N_3507);
nand U4511 (N_4511,N_3171,N_3556);
nor U4512 (N_4512,N_3853,N_3255);
nand U4513 (N_4513,N_3733,N_3599);
or U4514 (N_4514,N_3877,N_3863);
and U4515 (N_4515,N_3562,N_3508);
or U4516 (N_4516,N_3472,N_3065);
nor U4517 (N_4517,N_3001,N_3145);
and U4518 (N_4518,N_3670,N_3487);
or U4519 (N_4519,N_3921,N_3030);
nor U4520 (N_4520,N_3728,N_3972);
and U4521 (N_4521,N_3986,N_3084);
or U4522 (N_4522,N_3690,N_3139);
nand U4523 (N_4523,N_3465,N_3246);
and U4524 (N_4524,N_3994,N_3527);
nand U4525 (N_4525,N_3482,N_3098);
or U4526 (N_4526,N_3767,N_3318);
or U4527 (N_4527,N_3140,N_3709);
xnor U4528 (N_4528,N_3137,N_3848);
nor U4529 (N_4529,N_3845,N_3105);
or U4530 (N_4530,N_3893,N_3745);
and U4531 (N_4531,N_3625,N_3195);
nand U4532 (N_4532,N_3600,N_3044);
nor U4533 (N_4533,N_3763,N_3382);
nand U4534 (N_4534,N_3397,N_3318);
nand U4535 (N_4535,N_3675,N_3418);
nor U4536 (N_4536,N_3239,N_3320);
or U4537 (N_4537,N_3118,N_3653);
nor U4538 (N_4538,N_3804,N_3457);
nand U4539 (N_4539,N_3335,N_3649);
nor U4540 (N_4540,N_3847,N_3559);
or U4541 (N_4541,N_3295,N_3365);
nor U4542 (N_4542,N_3352,N_3222);
nor U4543 (N_4543,N_3171,N_3051);
nand U4544 (N_4544,N_3999,N_3641);
nor U4545 (N_4545,N_3786,N_3251);
nand U4546 (N_4546,N_3093,N_3341);
or U4547 (N_4547,N_3074,N_3159);
nor U4548 (N_4548,N_3046,N_3698);
nand U4549 (N_4549,N_3798,N_3990);
and U4550 (N_4550,N_3663,N_3373);
or U4551 (N_4551,N_3508,N_3209);
nand U4552 (N_4552,N_3486,N_3626);
nand U4553 (N_4553,N_3262,N_3705);
nand U4554 (N_4554,N_3517,N_3979);
and U4555 (N_4555,N_3652,N_3104);
nand U4556 (N_4556,N_3044,N_3268);
or U4557 (N_4557,N_3493,N_3525);
or U4558 (N_4558,N_3323,N_3745);
nand U4559 (N_4559,N_3614,N_3647);
and U4560 (N_4560,N_3972,N_3594);
nand U4561 (N_4561,N_3122,N_3650);
nor U4562 (N_4562,N_3060,N_3212);
and U4563 (N_4563,N_3171,N_3273);
nand U4564 (N_4564,N_3519,N_3590);
and U4565 (N_4565,N_3601,N_3345);
and U4566 (N_4566,N_3445,N_3388);
and U4567 (N_4567,N_3349,N_3757);
nand U4568 (N_4568,N_3637,N_3561);
nand U4569 (N_4569,N_3337,N_3633);
xor U4570 (N_4570,N_3154,N_3651);
nand U4571 (N_4571,N_3204,N_3032);
or U4572 (N_4572,N_3557,N_3172);
nand U4573 (N_4573,N_3085,N_3062);
nor U4574 (N_4574,N_3891,N_3622);
nand U4575 (N_4575,N_3707,N_3885);
or U4576 (N_4576,N_3096,N_3917);
nor U4577 (N_4577,N_3215,N_3859);
nand U4578 (N_4578,N_3111,N_3928);
nand U4579 (N_4579,N_3754,N_3374);
nand U4580 (N_4580,N_3634,N_3425);
nor U4581 (N_4581,N_3131,N_3481);
and U4582 (N_4582,N_3495,N_3509);
or U4583 (N_4583,N_3794,N_3330);
nand U4584 (N_4584,N_3146,N_3737);
nand U4585 (N_4585,N_3091,N_3203);
nor U4586 (N_4586,N_3184,N_3852);
and U4587 (N_4587,N_3124,N_3268);
nand U4588 (N_4588,N_3522,N_3436);
or U4589 (N_4589,N_3801,N_3711);
nor U4590 (N_4590,N_3635,N_3261);
or U4591 (N_4591,N_3448,N_3411);
nand U4592 (N_4592,N_3541,N_3998);
or U4593 (N_4593,N_3446,N_3353);
and U4594 (N_4594,N_3367,N_3835);
or U4595 (N_4595,N_3707,N_3963);
or U4596 (N_4596,N_3359,N_3725);
nand U4597 (N_4597,N_3764,N_3515);
xor U4598 (N_4598,N_3312,N_3836);
xor U4599 (N_4599,N_3319,N_3421);
nand U4600 (N_4600,N_3697,N_3185);
nor U4601 (N_4601,N_3921,N_3418);
nor U4602 (N_4602,N_3775,N_3774);
and U4603 (N_4603,N_3179,N_3143);
and U4604 (N_4604,N_3839,N_3443);
nor U4605 (N_4605,N_3645,N_3440);
nor U4606 (N_4606,N_3759,N_3664);
xnor U4607 (N_4607,N_3012,N_3802);
nand U4608 (N_4608,N_3393,N_3537);
nand U4609 (N_4609,N_3711,N_3718);
or U4610 (N_4610,N_3682,N_3744);
or U4611 (N_4611,N_3464,N_3931);
and U4612 (N_4612,N_3697,N_3355);
nor U4613 (N_4613,N_3954,N_3275);
nand U4614 (N_4614,N_3380,N_3680);
and U4615 (N_4615,N_3512,N_3030);
nand U4616 (N_4616,N_3319,N_3220);
nor U4617 (N_4617,N_3716,N_3754);
or U4618 (N_4618,N_3925,N_3433);
xnor U4619 (N_4619,N_3753,N_3900);
xnor U4620 (N_4620,N_3841,N_3068);
or U4621 (N_4621,N_3891,N_3763);
or U4622 (N_4622,N_3069,N_3820);
nor U4623 (N_4623,N_3569,N_3950);
nor U4624 (N_4624,N_3923,N_3197);
and U4625 (N_4625,N_3121,N_3850);
nand U4626 (N_4626,N_3833,N_3813);
nand U4627 (N_4627,N_3851,N_3450);
nor U4628 (N_4628,N_3316,N_3410);
and U4629 (N_4629,N_3789,N_3462);
or U4630 (N_4630,N_3237,N_3175);
and U4631 (N_4631,N_3920,N_3171);
nand U4632 (N_4632,N_3005,N_3473);
and U4633 (N_4633,N_3133,N_3066);
nor U4634 (N_4634,N_3359,N_3001);
and U4635 (N_4635,N_3057,N_3551);
nor U4636 (N_4636,N_3720,N_3514);
and U4637 (N_4637,N_3438,N_3444);
nor U4638 (N_4638,N_3493,N_3860);
or U4639 (N_4639,N_3235,N_3537);
nand U4640 (N_4640,N_3195,N_3058);
nor U4641 (N_4641,N_3774,N_3117);
and U4642 (N_4642,N_3202,N_3796);
and U4643 (N_4643,N_3252,N_3276);
and U4644 (N_4644,N_3355,N_3712);
and U4645 (N_4645,N_3141,N_3095);
or U4646 (N_4646,N_3579,N_3034);
and U4647 (N_4647,N_3827,N_3401);
nor U4648 (N_4648,N_3388,N_3231);
nand U4649 (N_4649,N_3672,N_3786);
and U4650 (N_4650,N_3034,N_3101);
or U4651 (N_4651,N_3587,N_3292);
or U4652 (N_4652,N_3304,N_3538);
nor U4653 (N_4653,N_3970,N_3576);
xor U4654 (N_4654,N_3753,N_3824);
and U4655 (N_4655,N_3980,N_3974);
nor U4656 (N_4656,N_3529,N_3740);
nor U4657 (N_4657,N_3587,N_3586);
and U4658 (N_4658,N_3312,N_3979);
and U4659 (N_4659,N_3579,N_3258);
nor U4660 (N_4660,N_3684,N_3732);
or U4661 (N_4661,N_3091,N_3948);
and U4662 (N_4662,N_3192,N_3069);
or U4663 (N_4663,N_3242,N_3988);
nor U4664 (N_4664,N_3406,N_3125);
and U4665 (N_4665,N_3242,N_3238);
or U4666 (N_4666,N_3180,N_3769);
nand U4667 (N_4667,N_3472,N_3238);
nand U4668 (N_4668,N_3604,N_3774);
nand U4669 (N_4669,N_3518,N_3706);
and U4670 (N_4670,N_3782,N_3405);
and U4671 (N_4671,N_3551,N_3660);
nand U4672 (N_4672,N_3082,N_3048);
nor U4673 (N_4673,N_3529,N_3098);
or U4674 (N_4674,N_3594,N_3777);
or U4675 (N_4675,N_3462,N_3143);
xnor U4676 (N_4676,N_3824,N_3379);
or U4677 (N_4677,N_3874,N_3274);
nand U4678 (N_4678,N_3107,N_3068);
nor U4679 (N_4679,N_3916,N_3492);
nand U4680 (N_4680,N_3281,N_3856);
and U4681 (N_4681,N_3914,N_3508);
and U4682 (N_4682,N_3556,N_3546);
or U4683 (N_4683,N_3146,N_3537);
or U4684 (N_4684,N_3121,N_3719);
or U4685 (N_4685,N_3492,N_3143);
nand U4686 (N_4686,N_3057,N_3777);
and U4687 (N_4687,N_3420,N_3864);
or U4688 (N_4688,N_3788,N_3747);
or U4689 (N_4689,N_3037,N_3610);
or U4690 (N_4690,N_3886,N_3044);
nand U4691 (N_4691,N_3009,N_3397);
nor U4692 (N_4692,N_3001,N_3259);
and U4693 (N_4693,N_3195,N_3403);
nor U4694 (N_4694,N_3661,N_3477);
nand U4695 (N_4695,N_3889,N_3510);
nor U4696 (N_4696,N_3552,N_3546);
and U4697 (N_4697,N_3638,N_3800);
or U4698 (N_4698,N_3255,N_3011);
nor U4699 (N_4699,N_3279,N_3275);
or U4700 (N_4700,N_3845,N_3338);
nor U4701 (N_4701,N_3476,N_3428);
nor U4702 (N_4702,N_3914,N_3434);
nand U4703 (N_4703,N_3849,N_3930);
nor U4704 (N_4704,N_3091,N_3035);
and U4705 (N_4705,N_3076,N_3098);
or U4706 (N_4706,N_3320,N_3911);
and U4707 (N_4707,N_3381,N_3607);
nor U4708 (N_4708,N_3759,N_3626);
and U4709 (N_4709,N_3049,N_3665);
nand U4710 (N_4710,N_3519,N_3286);
nor U4711 (N_4711,N_3196,N_3967);
and U4712 (N_4712,N_3560,N_3464);
nor U4713 (N_4713,N_3242,N_3860);
nand U4714 (N_4714,N_3203,N_3621);
nor U4715 (N_4715,N_3405,N_3065);
nor U4716 (N_4716,N_3658,N_3593);
xor U4717 (N_4717,N_3071,N_3782);
nor U4718 (N_4718,N_3198,N_3756);
nand U4719 (N_4719,N_3208,N_3868);
and U4720 (N_4720,N_3563,N_3725);
nor U4721 (N_4721,N_3592,N_3877);
and U4722 (N_4722,N_3296,N_3479);
nand U4723 (N_4723,N_3961,N_3950);
nor U4724 (N_4724,N_3386,N_3677);
nor U4725 (N_4725,N_3595,N_3269);
nand U4726 (N_4726,N_3585,N_3762);
nor U4727 (N_4727,N_3335,N_3163);
or U4728 (N_4728,N_3772,N_3803);
or U4729 (N_4729,N_3188,N_3531);
and U4730 (N_4730,N_3701,N_3735);
nand U4731 (N_4731,N_3061,N_3399);
and U4732 (N_4732,N_3462,N_3662);
nor U4733 (N_4733,N_3230,N_3952);
nand U4734 (N_4734,N_3859,N_3166);
and U4735 (N_4735,N_3881,N_3188);
nor U4736 (N_4736,N_3286,N_3490);
nor U4737 (N_4737,N_3533,N_3564);
nand U4738 (N_4738,N_3892,N_3895);
or U4739 (N_4739,N_3476,N_3300);
or U4740 (N_4740,N_3044,N_3741);
nand U4741 (N_4741,N_3601,N_3173);
nor U4742 (N_4742,N_3660,N_3101);
xor U4743 (N_4743,N_3569,N_3037);
or U4744 (N_4744,N_3687,N_3617);
and U4745 (N_4745,N_3453,N_3538);
nand U4746 (N_4746,N_3094,N_3884);
and U4747 (N_4747,N_3050,N_3886);
xor U4748 (N_4748,N_3242,N_3052);
or U4749 (N_4749,N_3245,N_3644);
nor U4750 (N_4750,N_3323,N_3201);
nor U4751 (N_4751,N_3820,N_3505);
or U4752 (N_4752,N_3843,N_3925);
nand U4753 (N_4753,N_3133,N_3436);
and U4754 (N_4754,N_3520,N_3332);
nor U4755 (N_4755,N_3209,N_3409);
or U4756 (N_4756,N_3451,N_3708);
and U4757 (N_4757,N_3986,N_3348);
and U4758 (N_4758,N_3733,N_3231);
or U4759 (N_4759,N_3222,N_3916);
and U4760 (N_4760,N_3781,N_3831);
or U4761 (N_4761,N_3738,N_3392);
and U4762 (N_4762,N_3524,N_3883);
or U4763 (N_4763,N_3052,N_3082);
nor U4764 (N_4764,N_3114,N_3491);
nand U4765 (N_4765,N_3861,N_3019);
and U4766 (N_4766,N_3013,N_3261);
or U4767 (N_4767,N_3056,N_3852);
nor U4768 (N_4768,N_3502,N_3123);
nor U4769 (N_4769,N_3616,N_3024);
nor U4770 (N_4770,N_3282,N_3956);
nor U4771 (N_4771,N_3090,N_3354);
and U4772 (N_4772,N_3942,N_3357);
nand U4773 (N_4773,N_3037,N_3169);
and U4774 (N_4774,N_3725,N_3287);
or U4775 (N_4775,N_3643,N_3810);
nor U4776 (N_4776,N_3022,N_3846);
and U4777 (N_4777,N_3474,N_3713);
nor U4778 (N_4778,N_3331,N_3509);
nand U4779 (N_4779,N_3820,N_3594);
and U4780 (N_4780,N_3810,N_3528);
nand U4781 (N_4781,N_3699,N_3146);
or U4782 (N_4782,N_3692,N_3132);
and U4783 (N_4783,N_3913,N_3982);
and U4784 (N_4784,N_3288,N_3378);
and U4785 (N_4785,N_3869,N_3635);
or U4786 (N_4786,N_3164,N_3339);
and U4787 (N_4787,N_3761,N_3149);
nand U4788 (N_4788,N_3090,N_3239);
nor U4789 (N_4789,N_3893,N_3062);
nand U4790 (N_4790,N_3363,N_3572);
nand U4791 (N_4791,N_3498,N_3681);
or U4792 (N_4792,N_3352,N_3929);
xor U4793 (N_4793,N_3546,N_3943);
nor U4794 (N_4794,N_3499,N_3196);
nor U4795 (N_4795,N_3736,N_3575);
and U4796 (N_4796,N_3477,N_3330);
nor U4797 (N_4797,N_3926,N_3196);
nor U4798 (N_4798,N_3060,N_3649);
or U4799 (N_4799,N_3402,N_3092);
nand U4800 (N_4800,N_3973,N_3339);
or U4801 (N_4801,N_3648,N_3222);
and U4802 (N_4802,N_3108,N_3725);
and U4803 (N_4803,N_3101,N_3613);
nor U4804 (N_4804,N_3849,N_3124);
nand U4805 (N_4805,N_3702,N_3972);
nand U4806 (N_4806,N_3138,N_3857);
nor U4807 (N_4807,N_3709,N_3645);
nor U4808 (N_4808,N_3610,N_3915);
nor U4809 (N_4809,N_3440,N_3093);
and U4810 (N_4810,N_3938,N_3066);
nand U4811 (N_4811,N_3189,N_3780);
or U4812 (N_4812,N_3320,N_3065);
nor U4813 (N_4813,N_3604,N_3069);
nor U4814 (N_4814,N_3847,N_3451);
or U4815 (N_4815,N_3638,N_3516);
or U4816 (N_4816,N_3994,N_3894);
nand U4817 (N_4817,N_3525,N_3546);
or U4818 (N_4818,N_3706,N_3858);
nand U4819 (N_4819,N_3403,N_3911);
nand U4820 (N_4820,N_3477,N_3919);
nor U4821 (N_4821,N_3018,N_3215);
or U4822 (N_4822,N_3355,N_3384);
xor U4823 (N_4823,N_3170,N_3805);
nor U4824 (N_4824,N_3756,N_3238);
and U4825 (N_4825,N_3383,N_3996);
or U4826 (N_4826,N_3488,N_3870);
nor U4827 (N_4827,N_3893,N_3378);
and U4828 (N_4828,N_3179,N_3556);
or U4829 (N_4829,N_3084,N_3440);
nand U4830 (N_4830,N_3641,N_3244);
or U4831 (N_4831,N_3365,N_3487);
nor U4832 (N_4832,N_3238,N_3877);
nor U4833 (N_4833,N_3321,N_3172);
or U4834 (N_4834,N_3447,N_3622);
and U4835 (N_4835,N_3604,N_3352);
or U4836 (N_4836,N_3265,N_3418);
or U4837 (N_4837,N_3495,N_3110);
nand U4838 (N_4838,N_3292,N_3711);
nor U4839 (N_4839,N_3472,N_3099);
and U4840 (N_4840,N_3774,N_3629);
nor U4841 (N_4841,N_3205,N_3278);
nor U4842 (N_4842,N_3034,N_3244);
xnor U4843 (N_4843,N_3908,N_3542);
or U4844 (N_4844,N_3570,N_3054);
and U4845 (N_4845,N_3755,N_3590);
or U4846 (N_4846,N_3935,N_3978);
nor U4847 (N_4847,N_3922,N_3196);
xnor U4848 (N_4848,N_3159,N_3906);
and U4849 (N_4849,N_3290,N_3074);
and U4850 (N_4850,N_3784,N_3667);
and U4851 (N_4851,N_3982,N_3256);
or U4852 (N_4852,N_3170,N_3491);
or U4853 (N_4853,N_3352,N_3149);
nand U4854 (N_4854,N_3286,N_3078);
nor U4855 (N_4855,N_3280,N_3770);
or U4856 (N_4856,N_3480,N_3777);
nand U4857 (N_4857,N_3992,N_3473);
xnor U4858 (N_4858,N_3134,N_3416);
or U4859 (N_4859,N_3784,N_3643);
and U4860 (N_4860,N_3876,N_3356);
or U4861 (N_4861,N_3180,N_3767);
or U4862 (N_4862,N_3796,N_3049);
nor U4863 (N_4863,N_3325,N_3327);
nor U4864 (N_4864,N_3748,N_3085);
and U4865 (N_4865,N_3612,N_3208);
nor U4866 (N_4866,N_3570,N_3816);
or U4867 (N_4867,N_3658,N_3441);
and U4868 (N_4868,N_3683,N_3387);
and U4869 (N_4869,N_3257,N_3527);
or U4870 (N_4870,N_3747,N_3706);
or U4871 (N_4871,N_3226,N_3539);
nand U4872 (N_4872,N_3751,N_3888);
and U4873 (N_4873,N_3955,N_3534);
nand U4874 (N_4874,N_3273,N_3195);
nor U4875 (N_4875,N_3124,N_3688);
or U4876 (N_4876,N_3816,N_3277);
and U4877 (N_4877,N_3386,N_3974);
nor U4878 (N_4878,N_3251,N_3124);
nor U4879 (N_4879,N_3331,N_3322);
nor U4880 (N_4880,N_3096,N_3671);
or U4881 (N_4881,N_3146,N_3654);
nor U4882 (N_4882,N_3732,N_3264);
or U4883 (N_4883,N_3721,N_3677);
nand U4884 (N_4884,N_3530,N_3861);
nor U4885 (N_4885,N_3940,N_3001);
nor U4886 (N_4886,N_3066,N_3285);
and U4887 (N_4887,N_3719,N_3672);
nor U4888 (N_4888,N_3317,N_3441);
or U4889 (N_4889,N_3722,N_3881);
or U4890 (N_4890,N_3208,N_3455);
nor U4891 (N_4891,N_3164,N_3858);
nor U4892 (N_4892,N_3808,N_3925);
or U4893 (N_4893,N_3004,N_3831);
and U4894 (N_4894,N_3761,N_3486);
and U4895 (N_4895,N_3456,N_3822);
or U4896 (N_4896,N_3605,N_3944);
or U4897 (N_4897,N_3565,N_3613);
nor U4898 (N_4898,N_3352,N_3240);
nand U4899 (N_4899,N_3189,N_3581);
nand U4900 (N_4900,N_3244,N_3215);
nor U4901 (N_4901,N_3516,N_3017);
nor U4902 (N_4902,N_3769,N_3039);
and U4903 (N_4903,N_3985,N_3277);
or U4904 (N_4904,N_3395,N_3587);
nand U4905 (N_4905,N_3506,N_3362);
nor U4906 (N_4906,N_3228,N_3962);
nand U4907 (N_4907,N_3476,N_3126);
nor U4908 (N_4908,N_3295,N_3815);
xor U4909 (N_4909,N_3616,N_3671);
nor U4910 (N_4910,N_3692,N_3512);
nor U4911 (N_4911,N_3027,N_3237);
nor U4912 (N_4912,N_3879,N_3660);
or U4913 (N_4913,N_3989,N_3850);
and U4914 (N_4914,N_3075,N_3151);
nand U4915 (N_4915,N_3060,N_3646);
nand U4916 (N_4916,N_3764,N_3976);
nand U4917 (N_4917,N_3282,N_3260);
or U4918 (N_4918,N_3277,N_3755);
and U4919 (N_4919,N_3595,N_3288);
nand U4920 (N_4920,N_3056,N_3978);
nor U4921 (N_4921,N_3044,N_3293);
or U4922 (N_4922,N_3796,N_3767);
xnor U4923 (N_4923,N_3609,N_3794);
nor U4924 (N_4924,N_3304,N_3889);
or U4925 (N_4925,N_3612,N_3135);
or U4926 (N_4926,N_3855,N_3371);
nor U4927 (N_4927,N_3820,N_3011);
nand U4928 (N_4928,N_3539,N_3013);
nand U4929 (N_4929,N_3901,N_3861);
and U4930 (N_4930,N_3633,N_3715);
and U4931 (N_4931,N_3225,N_3132);
and U4932 (N_4932,N_3093,N_3284);
nand U4933 (N_4933,N_3604,N_3568);
and U4934 (N_4934,N_3711,N_3502);
and U4935 (N_4935,N_3052,N_3857);
nor U4936 (N_4936,N_3657,N_3721);
and U4937 (N_4937,N_3299,N_3834);
nand U4938 (N_4938,N_3580,N_3283);
nor U4939 (N_4939,N_3695,N_3021);
and U4940 (N_4940,N_3987,N_3691);
xor U4941 (N_4941,N_3894,N_3890);
nand U4942 (N_4942,N_3737,N_3782);
or U4943 (N_4943,N_3332,N_3537);
nor U4944 (N_4944,N_3553,N_3377);
or U4945 (N_4945,N_3498,N_3701);
nor U4946 (N_4946,N_3468,N_3845);
and U4947 (N_4947,N_3703,N_3070);
nor U4948 (N_4948,N_3500,N_3838);
and U4949 (N_4949,N_3243,N_3849);
nand U4950 (N_4950,N_3401,N_3189);
nand U4951 (N_4951,N_3405,N_3881);
or U4952 (N_4952,N_3901,N_3060);
and U4953 (N_4953,N_3619,N_3196);
nand U4954 (N_4954,N_3558,N_3271);
and U4955 (N_4955,N_3115,N_3480);
nand U4956 (N_4956,N_3208,N_3905);
or U4957 (N_4957,N_3346,N_3119);
and U4958 (N_4958,N_3410,N_3413);
and U4959 (N_4959,N_3711,N_3614);
nor U4960 (N_4960,N_3465,N_3509);
or U4961 (N_4961,N_3075,N_3420);
xor U4962 (N_4962,N_3105,N_3617);
nand U4963 (N_4963,N_3767,N_3559);
or U4964 (N_4964,N_3720,N_3640);
nor U4965 (N_4965,N_3817,N_3320);
nand U4966 (N_4966,N_3333,N_3775);
or U4967 (N_4967,N_3609,N_3107);
nor U4968 (N_4968,N_3678,N_3547);
nand U4969 (N_4969,N_3966,N_3863);
or U4970 (N_4970,N_3046,N_3876);
nor U4971 (N_4971,N_3791,N_3129);
and U4972 (N_4972,N_3707,N_3299);
and U4973 (N_4973,N_3801,N_3399);
nor U4974 (N_4974,N_3135,N_3864);
and U4975 (N_4975,N_3435,N_3833);
xor U4976 (N_4976,N_3185,N_3227);
or U4977 (N_4977,N_3667,N_3374);
nand U4978 (N_4978,N_3689,N_3520);
and U4979 (N_4979,N_3001,N_3478);
nand U4980 (N_4980,N_3606,N_3005);
nand U4981 (N_4981,N_3845,N_3325);
or U4982 (N_4982,N_3196,N_3265);
and U4983 (N_4983,N_3939,N_3487);
and U4984 (N_4984,N_3688,N_3372);
nand U4985 (N_4985,N_3885,N_3900);
nand U4986 (N_4986,N_3456,N_3464);
nand U4987 (N_4987,N_3593,N_3415);
and U4988 (N_4988,N_3250,N_3387);
or U4989 (N_4989,N_3888,N_3698);
nor U4990 (N_4990,N_3835,N_3815);
nand U4991 (N_4991,N_3976,N_3107);
nand U4992 (N_4992,N_3740,N_3358);
and U4993 (N_4993,N_3332,N_3121);
or U4994 (N_4994,N_3402,N_3707);
and U4995 (N_4995,N_3104,N_3060);
nand U4996 (N_4996,N_3951,N_3053);
nand U4997 (N_4997,N_3393,N_3994);
nor U4998 (N_4998,N_3866,N_3253);
nor U4999 (N_4999,N_3180,N_3050);
and U5000 (N_5000,N_4033,N_4678);
nor U5001 (N_5001,N_4928,N_4924);
nor U5002 (N_5002,N_4329,N_4335);
and U5003 (N_5003,N_4691,N_4814);
nand U5004 (N_5004,N_4470,N_4762);
and U5005 (N_5005,N_4885,N_4829);
nand U5006 (N_5006,N_4643,N_4874);
nand U5007 (N_5007,N_4913,N_4644);
nand U5008 (N_5008,N_4901,N_4249);
nor U5009 (N_5009,N_4992,N_4245);
nand U5010 (N_5010,N_4319,N_4324);
or U5011 (N_5011,N_4039,N_4440);
nand U5012 (N_5012,N_4174,N_4226);
and U5013 (N_5013,N_4731,N_4742);
nand U5014 (N_5014,N_4070,N_4252);
or U5015 (N_5015,N_4612,N_4600);
nor U5016 (N_5016,N_4301,N_4472);
or U5017 (N_5017,N_4498,N_4950);
and U5018 (N_5018,N_4476,N_4930);
xor U5019 (N_5019,N_4149,N_4812);
or U5020 (N_5020,N_4591,N_4859);
and U5021 (N_5021,N_4135,N_4271);
or U5022 (N_5022,N_4671,N_4881);
and U5023 (N_5023,N_4598,N_4270);
and U5024 (N_5024,N_4703,N_4247);
nand U5025 (N_5025,N_4791,N_4720);
nor U5026 (N_5026,N_4755,N_4892);
and U5027 (N_5027,N_4768,N_4403);
and U5028 (N_5028,N_4852,N_4743);
nor U5029 (N_5029,N_4434,N_4680);
nor U5030 (N_5030,N_4348,N_4134);
nor U5031 (N_5031,N_4053,N_4546);
and U5032 (N_5032,N_4845,N_4758);
xor U5033 (N_5033,N_4137,N_4839);
nor U5034 (N_5034,N_4266,N_4543);
nand U5035 (N_5035,N_4296,N_4336);
or U5036 (N_5036,N_4002,N_4902);
and U5037 (N_5037,N_4347,N_4798);
and U5038 (N_5038,N_4565,N_4869);
nand U5039 (N_5039,N_4450,N_4047);
and U5040 (N_5040,N_4352,N_4147);
or U5041 (N_5041,N_4970,N_4382);
nand U5042 (N_5042,N_4710,N_4824);
nor U5043 (N_5043,N_4133,N_4255);
or U5044 (N_5044,N_4281,N_4508);
nand U5045 (N_5045,N_4310,N_4017);
or U5046 (N_5046,N_4927,N_4512);
and U5047 (N_5047,N_4549,N_4104);
nor U5048 (N_5048,N_4171,N_4421);
nor U5049 (N_5049,N_4273,N_4894);
and U5050 (N_5050,N_4192,N_4142);
nand U5051 (N_5051,N_4878,N_4254);
and U5052 (N_5052,N_4673,N_4536);
nand U5053 (N_5053,N_4694,N_4682);
nand U5054 (N_5054,N_4425,N_4111);
nand U5055 (N_5055,N_4260,N_4771);
nor U5056 (N_5056,N_4917,N_4915);
nor U5057 (N_5057,N_4553,N_4451);
or U5058 (N_5058,N_4144,N_4642);
and U5059 (N_5059,N_4856,N_4225);
or U5060 (N_5060,N_4564,N_4297);
and U5061 (N_5061,N_4724,N_4173);
and U5062 (N_5062,N_4853,N_4474);
and U5063 (N_5063,N_4344,N_4195);
and U5064 (N_5064,N_4263,N_4080);
or U5065 (N_5065,N_4960,N_4105);
nand U5066 (N_5066,N_4308,N_4582);
and U5067 (N_5067,N_4064,N_4230);
nor U5068 (N_5068,N_4674,N_4587);
nand U5069 (N_5069,N_4740,N_4730);
or U5070 (N_5070,N_4416,N_4999);
or U5071 (N_5071,N_4665,N_4646);
or U5072 (N_5072,N_4690,N_4184);
nor U5073 (N_5073,N_4815,N_4353);
or U5074 (N_5074,N_4054,N_4211);
or U5075 (N_5075,N_4407,N_4338);
and U5076 (N_5076,N_4361,N_4622);
nor U5077 (N_5077,N_4548,N_4728);
or U5078 (N_5078,N_4057,N_4699);
and U5079 (N_5079,N_4649,N_4656);
nor U5080 (N_5080,N_4129,N_4075);
nand U5081 (N_5081,N_4428,N_4065);
nand U5082 (N_5082,N_4029,N_4368);
xnor U5083 (N_5083,N_4957,N_4882);
and U5084 (N_5084,N_4519,N_4365);
or U5085 (N_5085,N_4830,N_4590);
nor U5086 (N_5086,N_4817,N_4120);
nand U5087 (N_5087,N_4351,N_4007);
and U5088 (N_5088,N_4109,N_4966);
or U5089 (N_5089,N_4496,N_4187);
xnor U5090 (N_5090,N_4355,N_4052);
nor U5091 (N_5091,N_4183,N_4194);
or U5092 (N_5092,N_4130,N_4323);
nor U5093 (N_5093,N_4953,N_4949);
nand U5094 (N_5094,N_4232,N_4342);
and U5095 (N_5095,N_4293,N_4588);
or U5096 (N_5096,N_4875,N_4110);
nand U5097 (N_5097,N_4715,N_4454);
and U5098 (N_5098,N_4555,N_4776);
nor U5099 (N_5099,N_4589,N_4290);
nor U5100 (N_5100,N_4401,N_4480);
nor U5101 (N_5101,N_4529,N_4586);
xnor U5102 (N_5102,N_4288,N_4006);
nor U5103 (N_5103,N_4838,N_4973);
or U5104 (N_5104,N_4855,N_4727);
nor U5105 (N_5105,N_4364,N_4018);
nand U5106 (N_5106,N_4981,N_4637);
nor U5107 (N_5107,N_4544,N_4377);
or U5108 (N_5108,N_4578,N_4667);
nand U5109 (N_5109,N_4576,N_4639);
xnor U5110 (N_5110,N_4531,N_4096);
and U5111 (N_5111,N_4114,N_4038);
nor U5112 (N_5112,N_4085,N_4797);
nor U5113 (N_5113,N_4148,N_4444);
nor U5114 (N_5114,N_4995,N_4443);
or U5115 (N_5115,N_4062,N_4094);
and U5116 (N_5116,N_4487,N_4510);
and U5117 (N_5117,N_4445,N_4827);
nand U5118 (N_5118,N_4807,N_4532);
nor U5119 (N_5119,N_4438,N_4251);
and U5120 (N_5120,N_4891,N_4372);
xor U5121 (N_5121,N_4567,N_4920);
nand U5122 (N_5122,N_4721,N_4880);
nand U5123 (N_5123,N_4936,N_4371);
or U5124 (N_5124,N_4534,N_4153);
nand U5125 (N_5125,N_4628,N_4975);
or U5126 (N_5126,N_4800,N_4491);
xnor U5127 (N_5127,N_4471,N_4528);
xnor U5128 (N_5128,N_4884,N_4557);
and U5129 (N_5129,N_4219,N_4654);
or U5130 (N_5130,N_4046,N_4909);
nor U5131 (N_5131,N_4131,N_4573);
xor U5132 (N_5132,N_4895,N_4424);
or U5133 (N_5133,N_4616,N_4193);
or U5134 (N_5134,N_4942,N_4116);
and U5135 (N_5135,N_4442,N_4751);
and U5136 (N_5136,N_4926,N_4711);
nor U5137 (N_5137,N_4068,N_4241);
nand U5138 (N_5138,N_4707,N_4785);
and U5139 (N_5139,N_4358,N_4516);
and U5140 (N_5140,N_4825,N_4087);
or U5141 (N_5141,N_4581,N_4412);
xnor U5142 (N_5142,N_4620,N_4483);
xnor U5143 (N_5143,N_4359,N_4989);
and U5144 (N_5144,N_4823,N_4295);
nor U5145 (N_5145,N_4208,N_4466);
xnor U5146 (N_5146,N_4473,N_4441);
and U5147 (N_5147,N_4947,N_4747);
and U5148 (N_5148,N_4292,N_4593);
nor U5149 (N_5149,N_4239,N_4027);
or U5150 (N_5150,N_4410,N_4313);
nor U5151 (N_5151,N_4312,N_4765);
and U5152 (N_5152,N_4826,N_4687);
or U5153 (N_5153,N_4294,N_4127);
nand U5154 (N_5154,N_4340,N_4634);
or U5155 (N_5155,N_4954,N_4925);
or U5156 (N_5156,N_4860,N_4228);
xnor U5157 (N_5157,N_4962,N_4077);
or U5158 (N_5158,N_4074,N_4864);
and U5159 (N_5159,N_4339,N_4242);
nand U5160 (N_5160,N_4501,N_4161);
or U5161 (N_5161,N_4788,N_4782);
nand U5162 (N_5162,N_4097,N_4088);
or U5163 (N_5163,N_4202,N_4533);
nor U5164 (N_5164,N_4152,N_4786);
nor U5165 (N_5165,N_4659,N_4139);
nand U5166 (N_5166,N_4155,N_4630);
and U5167 (N_5167,N_4822,N_4906);
xnor U5168 (N_5168,N_4118,N_4922);
nor U5169 (N_5169,N_4803,N_4774);
nor U5170 (N_5170,N_4019,N_4349);
or U5171 (N_5171,N_4931,N_4490);
or U5172 (N_5172,N_4267,N_4331);
xnor U5173 (N_5173,N_4167,N_4221);
nor U5174 (N_5174,N_4705,N_4503);
and U5175 (N_5175,N_4092,N_4988);
nand U5176 (N_5176,N_4051,N_4840);
or U5177 (N_5177,N_4597,N_4769);
xor U5178 (N_5178,N_4413,N_4240);
nand U5179 (N_5179,N_4050,N_4504);
nand U5180 (N_5180,N_4126,N_4967);
and U5181 (N_5181,N_4898,N_4662);
or U5182 (N_5182,N_4712,N_4737);
nor U5183 (N_5183,N_4513,N_4735);
and U5184 (N_5184,N_4778,N_4961);
and U5185 (N_5185,N_4063,N_4089);
and U5186 (N_5186,N_4043,N_4676);
or U5187 (N_5187,N_4579,N_4157);
or U5188 (N_5188,N_4763,N_4964);
and U5189 (N_5189,N_4541,N_4857);
nor U5190 (N_5190,N_4602,N_4390);
nor U5191 (N_5191,N_4831,N_4783);
nor U5192 (N_5192,N_4370,N_4458);
or U5193 (N_5193,N_4469,N_4849);
and U5194 (N_5194,N_4623,N_4436);
and U5195 (N_5195,N_4258,N_4484);
nand U5196 (N_5196,N_4283,N_4492);
or U5197 (N_5197,N_4617,N_4414);
or U5198 (N_5198,N_4790,N_4760);
and U5199 (N_5199,N_4610,N_4816);
and U5200 (N_5200,N_4515,N_4181);
or U5201 (N_5201,N_4409,N_4350);
nand U5202 (N_5202,N_4482,N_4556);
and U5203 (N_5203,N_4393,N_4431);
or U5204 (N_5204,N_4124,N_4383);
nor U5205 (N_5205,N_4276,N_4986);
and U5206 (N_5206,N_4601,N_4369);
nor U5207 (N_5207,N_4095,N_4757);
or U5208 (N_5208,N_4614,N_4214);
nor U5209 (N_5209,N_4893,N_4236);
nor U5210 (N_5210,N_4011,N_4958);
and U5211 (N_5211,N_4714,N_4980);
nor U5212 (N_5212,N_4701,N_4575);
or U5213 (N_5213,N_4668,N_4341);
nor U5214 (N_5214,N_4268,N_4327);
nor U5215 (N_5215,N_4172,N_4044);
nand U5216 (N_5216,N_4117,N_4854);
or U5217 (N_5217,N_4794,N_4269);
nand U5218 (N_5218,N_4346,N_4993);
nor U5219 (N_5219,N_4708,N_4309);
and U5220 (N_5220,N_4012,N_4819);
or U5221 (N_5221,N_4698,N_4220);
or U5222 (N_5222,N_4923,N_4389);
nor U5223 (N_5223,N_4851,N_4262);
nor U5224 (N_5224,N_4625,N_4619);
and U5225 (N_5225,N_4222,N_4385);
or U5226 (N_5226,N_4217,N_4021);
nand U5227 (N_5227,N_4767,N_4937);
or U5228 (N_5228,N_4387,N_4813);
nand U5229 (N_5229,N_4595,N_4569);
and U5230 (N_5230,N_4561,N_4979);
nand U5231 (N_5231,N_4603,N_4653);
nor U5232 (N_5232,N_4231,N_4605);
nor U5233 (N_5233,N_4804,N_4031);
and U5234 (N_5234,N_4672,N_4560);
nor U5235 (N_5235,N_4005,N_4462);
nand U5236 (N_5236,N_4216,N_4078);
nand U5237 (N_5237,N_4990,N_4460);
nand U5238 (N_5238,N_4468,N_4795);
nor U5239 (N_5239,N_4257,N_4761);
and U5240 (N_5240,N_4086,N_4688);
and U5241 (N_5241,N_4867,N_4974);
nor U5242 (N_5242,N_4596,N_4160);
or U5243 (N_5243,N_4305,N_4554);
or U5244 (N_5244,N_4879,N_4233);
and U5245 (N_5245,N_4186,N_4526);
nor U5246 (N_5246,N_4218,N_4150);
nand U5247 (N_5247,N_4861,N_4360);
nand U5248 (N_5248,N_4475,N_4844);
and U5249 (N_5249,N_4343,N_4396);
and U5250 (N_5250,N_4618,N_4417);
or U5251 (N_5251,N_4833,N_4481);
xnor U5252 (N_5252,N_4572,N_4704);
and U5253 (N_5253,N_4380,N_4584);
or U5254 (N_5254,N_4061,N_4518);
or U5255 (N_5255,N_4523,N_4318);
and U5256 (N_5256,N_4729,N_4537);
or U5257 (N_5257,N_4356,N_4180);
nor U5258 (N_5258,N_4169,N_4099);
nor U5259 (N_5259,N_4400,N_4877);
and U5260 (N_5260,N_4448,N_4415);
nor U5261 (N_5261,N_4430,N_4820);
and U5262 (N_5262,N_4014,N_4681);
nand U5263 (N_5263,N_4032,N_4899);
nand U5264 (N_5264,N_4456,N_4502);
or U5265 (N_5265,N_4736,N_4635);
nand U5266 (N_5266,N_4397,N_4550);
and U5267 (N_5267,N_4754,N_4189);
nor U5268 (N_5268,N_4810,N_4780);
nand U5269 (N_5269,N_4395,N_4801);
nand U5270 (N_5270,N_4237,N_4522);
and U5271 (N_5271,N_4284,N_4259);
and U5272 (N_5272,N_4559,N_4386);
xor U5273 (N_5273,N_4873,N_4102);
and U5274 (N_5274,N_4170,N_4796);
nor U5275 (N_5275,N_4624,N_4896);
or U5276 (N_5276,N_4322,N_4100);
nor U5277 (N_5277,N_4082,N_4055);
or U5278 (N_5278,N_4982,N_4889);
nand U5279 (N_5279,N_4022,N_4463);
or U5280 (N_5280,N_4744,N_4373);
nor U5281 (N_5281,N_4378,N_4178);
nor U5282 (N_5282,N_4806,N_4594);
nand U5283 (N_5283,N_4366,N_4651);
or U5284 (N_5284,N_4278,N_4244);
or U5285 (N_5285,N_4081,N_4835);
nor U5286 (N_5286,N_4770,N_4337);
nor U5287 (N_5287,N_4916,N_4107);
or U5288 (N_5288,N_4627,N_4275);
or U5289 (N_5289,N_4374,N_4955);
or U5290 (N_5290,N_4607,N_4566);
nor U5291 (N_5291,N_4158,N_4067);
or U5292 (N_5292,N_4459,N_4048);
or U5293 (N_5293,N_4427,N_4141);
nand U5294 (N_5294,N_4479,N_4629);
nand U5295 (N_5295,N_4328,N_4084);
and U5296 (N_5296,N_4787,N_4314);
nor U5297 (N_5297,N_4570,N_4119);
nor U5298 (N_5298,N_4224,N_4453);
and U5299 (N_5299,N_4745,N_4223);
or U5300 (N_5300,N_4315,N_4606);
and U5301 (N_5301,N_4773,N_4429);
or U5302 (N_5302,N_4154,N_4449);
nand U5303 (N_5303,N_4660,N_4320);
or U5304 (N_5304,N_4886,N_4212);
and U5305 (N_5305,N_4166,N_4702);
nor U5306 (N_5306,N_4836,N_4398);
and U5307 (N_5307,N_4072,N_4904);
nand U5308 (N_5308,N_4406,N_4025);
and U5309 (N_5309,N_4201,N_4739);
nand U5310 (N_5310,N_4903,N_4488);
nor U5311 (N_5311,N_4197,N_4959);
or U5312 (N_5312,N_4034,N_4779);
nor U5313 (N_5313,N_4741,N_4805);
nand U5314 (N_5314,N_4689,N_4028);
or U5315 (N_5315,N_4015,N_4326);
nand U5316 (N_5316,N_4121,N_4000);
nor U5317 (N_5317,N_4821,N_4209);
nor U5318 (N_5318,N_4302,N_4766);
nor U5319 (N_5319,N_4514,N_4041);
nand U5320 (N_5320,N_4272,N_4792);
or U5321 (N_5321,N_4264,N_4932);
and U5322 (N_5322,N_4775,N_4843);
or U5323 (N_5323,N_4935,N_4538);
nor U5324 (N_5324,N_4500,N_4367);
nand U5325 (N_5325,N_4306,N_4168);
and U5326 (N_5326,N_4024,N_4669);
nor U5327 (N_5327,N_4261,N_4571);
and U5328 (N_5328,N_4872,N_4405);
nand U5329 (N_5329,N_4563,N_4650);
or U5330 (N_5330,N_4963,N_4978);
or U5331 (N_5331,N_4693,N_4679);
nand U5332 (N_5332,N_4664,N_4948);
or U5333 (N_5333,N_4432,N_4495);
or U5334 (N_5334,N_4997,N_4307);
nand U5335 (N_5335,N_4887,N_4921);
and U5336 (N_5336,N_4738,N_4485);
nor U5337 (N_5337,N_4725,N_4493);
and U5338 (N_5338,N_4066,N_4182);
nor U5339 (N_5339,N_4098,N_4834);
nor U5340 (N_5340,N_4394,N_4723);
and U5341 (N_5341,N_4545,N_4511);
nor U5342 (N_5342,N_4842,N_4122);
and U5343 (N_5343,N_4143,N_4977);
nand U5344 (N_5344,N_4700,N_4733);
or U5345 (N_5345,N_4848,N_4049);
or U5346 (N_5346,N_4753,N_4863);
and U5347 (N_5347,N_4941,N_4379);
or U5348 (N_5348,N_4506,N_4036);
and U5349 (N_5349,N_4521,N_4001);
and U5350 (N_5350,N_4562,N_4621);
or U5351 (N_5351,N_4108,N_4083);
and U5352 (N_5352,N_4939,N_4115);
and U5353 (N_5353,N_4073,N_4140);
and U5354 (N_5354,N_4151,N_4497);
and U5355 (N_5355,N_4437,N_4717);
or U5356 (N_5356,N_4713,N_4539);
nand U5357 (N_5357,N_4091,N_4802);
and U5358 (N_5358,N_4008,N_4256);
nand U5359 (N_5359,N_4004,N_4552);
nand U5360 (N_5360,N_4663,N_4408);
or U5361 (N_5361,N_4190,N_4914);
nor U5362 (N_5362,N_4638,N_4832);
and U5363 (N_5363,N_4332,N_4695);
xor U5364 (N_5364,N_4238,N_4457);
nand U5365 (N_5365,N_4299,N_4608);
and U5366 (N_5366,N_4229,N_4330);
and U5367 (N_5367,N_4991,N_4363);
nand U5368 (N_5368,N_4862,N_4357);
nand U5369 (N_5369,N_4858,N_4298);
or U5370 (N_5370,N_4781,N_4568);
nor U5371 (N_5371,N_4868,N_4509);
and U5372 (N_5372,N_4009,N_4574);
or U5373 (N_5373,N_4666,N_4023);
nand U5374 (N_5374,N_4136,N_4113);
or U5375 (N_5375,N_4235,N_4994);
or U5376 (N_5376,N_4248,N_4900);
or U5377 (N_5377,N_4969,N_4447);
or U5378 (N_5378,N_4934,N_4888);
nor U5379 (N_5379,N_4507,N_4558);
and U5380 (N_5380,N_4227,N_4112);
and U5381 (N_5381,N_4285,N_4998);
nand U5382 (N_5382,N_4426,N_4722);
nand U5383 (N_5383,N_4686,N_4865);
or U5384 (N_5384,N_4984,N_4253);
nor U5385 (N_5385,N_4706,N_4030);
nor U5386 (N_5386,N_4641,N_4163);
nand U5387 (N_5387,N_4946,N_4246);
xor U5388 (N_5388,N_4035,N_4841);
and U5389 (N_5389,N_4101,N_4042);
nor U5390 (N_5390,N_4632,N_4274);
nor U5391 (N_5391,N_4210,N_4423);
nor U5392 (N_5392,N_4719,N_4837);
nand U5393 (N_5393,N_4477,N_4289);
and U5394 (N_5394,N_4317,N_4697);
nor U5395 (N_5395,N_4726,N_4734);
nor U5396 (N_5396,N_4996,N_4613);
and U5397 (N_5397,N_4658,N_4125);
or U5398 (N_5398,N_4846,N_4912);
nand U5399 (N_5399,N_4759,N_4200);
nand U5400 (N_5400,N_4334,N_4215);
nor U5401 (N_5401,N_4433,N_4933);
xor U5402 (N_5402,N_4972,N_4750);
xnor U5403 (N_5403,N_4583,N_4203);
nor U5404 (N_5404,N_4392,N_4684);
nand U5405 (N_5405,N_4478,N_4828);
and U5406 (N_5406,N_4876,N_4234);
and U5407 (N_5407,N_4615,N_4058);
nor U5408 (N_5408,N_4420,N_4648);
and U5409 (N_5409,N_4418,N_4951);
or U5410 (N_5410,N_4040,N_4388);
nor U5411 (N_5411,N_4090,N_4461);
nor U5412 (N_5412,N_4467,N_4908);
nor U5413 (N_5413,N_4709,N_4808);
nand U5414 (N_5414,N_4304,N_4185);
or U5415 (N_5415,N_4079,N_4499);
or U5416 (N_5416,N_4551,N_4633);
or U5417 (N_5417,N_4985,N_4291);
xnor U5418 (N_5418,N_4631,N_4419);
nand U5419 (N_5419,N_4199,N_4976);
nor U5420 (N_5420,N_4325,N_4696);
nor U5421 (N_5421,N_4455,N_4026);
or U5422 (N_5422,N_4685,N_4020);
nor U5423 (N_5423,N_4732,N_4940);
and U5424 (N_5424,N_4647,N_4530);
nor U5425 (N_5425,N_4045,N_4535);
nor U5426 (N_5426,N_4956,N_4243);
or U5427 (N_5427,N_4965,N_4422);
and U5428 (N_5428,N_4464,N_4316);
and U5429 (N_5429,N_4013,N_4784);
and U5430 (N_5430,N_4191,N_4446);
nand U5431 (N_5431,N_4945,N_4162);
or U5432 (N_5432,N_4159,N_4764);
and U5433 (N_5433,N_4897,N_4652);
nor U5434 (N_5434,N_4156,N_4003);
nand U5435 (N_5435,N_4103,N_4404);
or U5436 (N_5436,N_4179,N_4439);
and U5437 (N_5437,N_4345,N_4311);
nor U5438 (N_5438,N_4010,N_4918);
or U5439 (N_5439,N_4626,N_4205);
nand U5440 (N_5440,N_4196,N_4675);
and U5441 (N_5441,N_4883,N_4106);
or U5442 (N_5442,N_4213,N_4146);
nor U5443 (N_5443,N_4645,N_4016);
and U5444 (N_5444,N_4132,N_4391);
nand U5445 (N_5445,N_4093,N_4402);
or U5446 (N_5446,N_4716,N_4525);
nor U5447 (N_5447,N_4207,N_4677);
and U5448 (N_5448,N_4206,N_4749);
and U5449 (N_5449,N_4746,N_4056);
nand U5450 (N_5450,N_4076,N_4655);
nor U5451 (N_5451,N_4286,N_4282);
and U5452 (N_5452,N_4793,N_4748);
and U5453 (N_5453,N_4577,N_4718);
nor U5454 (N_5454,N_4585,N_4381);
xor U5455 (N_5455,N_4542,N_4300);
and U5456 (N_5456,N_4752,N_4069);
nor U5457 (N_5457,N_4599,N_4060);
nand U5458 (N_5458,N_4640,N_4683);
or U5459 (N_5459,N_4465,N_4609);
nor U5460 (N_5460,N_4850,N_4657);
nand U5461 (N_5461,N_4384,N_4910);
and U5462 (N_5462,N_4943,N_4435);
or U5463 (N_5463,N_4204,N_4517);
nor U5464 (N_5464,N_4452,N_4756);
and U5465 (N_5465,N_4128,N_4280);
and U5466 (N_5466,N_4164,N_4303);
or U5467 (N_5467,N_4799,N_4580);
nor U5468 (N_5468,N_4987,N_4362);
or U5469 (N_5469,N_4524,N_4354);
nand U5470 (N_5470,N_4983,N_4907);
nor U5471 (N_5471,N_4670,N_4138);
nor U5472 (N_5472,N_4919,N_4037);
or U5473 (N_5473,N_4944,N_4486);
xor U5474 (N_5474,N_4059,N_4177);
nor U5475 (N_5475,N_4279,N_4871);
xor U5476 (N_5476,N_4175,N_4399);
and U5477 (N_5477,N_4333,N_4188);
and U5478 (N_5478,N_4071,N_4494);
nor U5479 (N_5479,N_4489,N_4809);
nand U5480 (N_5480,N_4287,N_4968);
nand U5481 (N_5481,N_4905,N_4145);
and U5482 (N_5482,N_4971,N_4604);
or U5483 (N_5483,N_4265,N_4636);
nor U5484 (N_5484,N_4411,N_4811);
nor U5485 (N_5485,N_4952,N_4277);
nand U5486 (N_5486,N_4527,N_4890);
nand U5487 (N_5487,N_4540,N_4176);
or U5488 (N_5488,N_4250,N_4789);
and U5489 (N_5489,N_4592,N_4375);
nor U5490 (N_5490,N_4661,N_4847);
and U5491 (N_5491,N_4818,N_4611);
nor U5492 (N_5492,N_4505,N_4547);
and U5493 (N_5493,N_4870,N_4520);
or U5494 (N_5494,N_4772,N_4123);
nand U5495 (N_5495,N_4376,N_4692);
or U5496 (N_5496,N_4866,N_4777);
and U5497 (N_5497,N_4165,N_4938);
nor U5498 (N_5498,N_4911,N_4929);
or U5499 (N_5499,N_4198,N_4321);
or U5500 (N_5500,N_4449,N_4693);
or U5501 (N_5501,N_4837,N_4570);
or U5502 (N_5502,N_4186,N_4457);
nor U5503 (N_5503,N_4717,N_4132);
or U5504 (N_5504,N_4341,N_4484);
nor U5505 (N_5505,N_4412,N_4728);
nor U5506 (N_5506,N_4839,N_4336);
nor U5507 (N_5507,N_4460,N_4351);
and U5508 (N_5508,N_4697,N_4311);
nand U5509 (N_5509,N_4909,N_4442);
or U5510 (N_5510,N_4152,N_4516);
and U5511 (N_5511,N_4679,N_4191);
and U5512 (N_5512,N_4600,N_4998);
nand U5513 (N_5513,N_4461,N_4901);
or U5514 (N_5514,N_4366,N_4187);
and U5515 (N_5515,N_4331,N_4554);
nor U5516 (N_5516,N_4783,N_4330);
and U5517 (N_5517,N_4321,N_4448);
or U5518 (N_5518,N_4069,N_4239);
nand U5519 (N_5519,N_4946,N_4365);
nor U5520 (N_5520,N_4982,N_4974);
or U5521 (N_5521,N_4873,N_4254);
or U5522 (N_5522,N_4178,N_4960);
and U5523 (N_5523,N_4662,N_4545);
nand U5524 (N_5524,N_4750,N_4236);
or U5525 (N_5525,N_4641,N_4698);
nand U5526 (N_5526,N_4087,N_4158);
nand U5527 (N_5527,N_4096,N_4610);
or U5528 (N_5528,N_4941,N_4084);
or U5529 (N_5529,N_4101,N_4921);
or U5530 (N_5530,N_4182,N_4487);
nand U5531 (N_5531,N_4964,N_4248);
and U5532 (N_5532,N_4318,N_4810);
and U5533 (N_5533,N_4684,N_4969);
nor U5534 (N_5534,N_4847,N_4807);
and U5535 (N_5535,N_4310,N_4270);
nand U5536 (N_5536,N_4928,N_4418);
or U5537 (N_5537,N_4196,N_4411);
nand U5538 (N_5538,N_4737,N_4350);
or U5539 (N_5539,N_4357,N_4753);
and U5540 (N_5540,N_4942,N_4243);
nor U5541 (N_5541,N_4446,N_4805);
nor U5542 (N_5542,N_4421,N_4404);
and U5543 (N_5543,N_4539,N_4353);
nand U5544 (N_5544,N_4687,N_4477);
nor U5545 (N_5545,N_4965,N_4497);
nor U5546 (N_5546,N_4471,N_4561);
nand U5547 (N_5547,N_4223,N_4381);
and U5548 (N_5548,N_4040,N_4346);
nor U5549 (N_5549,N_4366,N_4257);
or U5550 (N_5550,N_4442,N_4193);
or U5551 (N_5551,N_4939,N_4560);
and U5552 (N_5552,N_4887,N_4218);
and U5553 (N_5553,N_4428,N_4549);
nand U5554 (N_5554,N_4549,N_4837);
nand U5555 (N_5555,N_4309,N_4183);
nand U5556 (N_5556,N_4505,N_4604);
nor U5557 (N_5557,N_4032,N_4188);
and U5558 (N_5558,N_4100,N_4081);
and U5559 (N_5559,N_4000,N_4968);
or U5560 (N_5560,N_4498,N_4465);
or U5561 (N_5561,N_4134,N_4448);
and U5562 (N_5562,N_4265,N_4374);
nand U5563 (N_5563,N_4765,N_4515);
nor U5564 (N_5564,N_4887,N_4889);
or U5565 (N_5565,N_4607,N_4741);
nand U5566 (N_5566,N_4986,N_4020);
or U5567 (N_5567,N_4761,N_4535);
and U5568 (N_5568,N_4569,N_4311);
nand U5569 (N_5569,N_4917,N_4772);
or U5570 (N_5570,N_4230,N_4423);
nand U5571 (N_5571,N_4517,N_4963);
or U5572 (N_5572,N_4395,N_4357);
xor U5573 (N_5573,N_4439,N_4199);
nor U5574 (N_5574,N_4421,N_4559);
and U5575 (N_5575,N_4380,N_4349);
nand U5576 (N_5576,N_4035,N_4936);
nand U5577 (N_5577,N_4931,N_4208);
nand U5578 (N_5578,N_4690,N_4944);
or U5579 (N_5579,N_4534,N_4580);
or U5580 (N_5580,N_4823,N_4439);
xnor U5581 (N_5581,N_4011,N_4986);
xor U5582 (N_5582,N_4266,N_4687);
nor U5583 (N_5583,N_4043,N_4875);
or U5584 (N_5584,N_4481,N_4694);
and U5585 (N_5585,N_4930,N_4367);
and U5586 (N_5586,N_4299,N_4216);
or U5587 (N_5587,N_4488,N_4384);
nor U5588 (N_5588,N_4415,N_4723);
and U5589 (N_5589,N_4542,N_4398);
xnor U5590 (N_5590,N_4506,N_4296);
or U5591 (N_5591,N_4507,N_4390);
or U5592 (N_5592,N_4682,N_4758);
nand U5593 (N_5593,N_4669,N_4989);
xor U5594 (N_5594,N_4939,N_4943);
or U5595 (N_5595,N_4861,N_4764);
xor U5596 (N_5596,N_4069,N_4259);
and U5597 (N_5597,N_4014,N_4330);
nor U5598 (N_5598,N_4348,N_4816);
or U5599 (N_5599,N_4278,N_4423);
nand U5600 (N_5600,N_4044,N_4928);
or U5601 (N_5601,N_4998,N_4395);
and U5602 (N_5602,N_4376,N_4662);
and U5603 (N_5603,N_4416,N_4746);
nor U5604 (N_5604,N_4952,N_4737);
nor U5605 (N_5605,N_4925,N_4483);
nand U5606 (N_5606,N_4839,N_4380);
nor U5607 (N_5607,N_4547,N_4852);
and U5608 (N_5608,N_4342,N_4089);
or U5609 (N_5609,N_4706,N_4269);
and U5610 (N_5610,N_4179,N_4469);
nor U5611 (N_5611,N_4359,N_4145);
or U5612 (N_5612,N_4761,N_4996);
or U5613 (N_5613,N_4231,N_4702);
nand U5614 (N_5614,N_4266,N_4468);
nor U5615 (N_5615,N_4735,N_4646);
nand U5616 (N_5616,N_4913,N_4949);
nor U5617 (N_5617,N_4059,N_4746);
nor U5618 (N_5618,N_4536,N_4616);
nand U5619 (N_5619,N_4100,N_4809);
nor U5620 (N_5620,N_4982,N_4112);
or U5621 (N_5621,N_4584,N_4759);
nand U5622 (N_5622,N_4194,N_4785);
and U5623 (N_5623,N_4600,N_4223);
or U5624 (N_5624,N_4495,N_4341);
nand U5625 (N_5625,N_4560,N_4653);
or U5626 (N_5626,N_4326,N_4949);
or U5627 (N_5627,N_4288,N_4414);
and U5628 (N_5628,N_4601,N_4241);
or U5629 (N_5629,N_4589,N_4612);
and U5630 (N_5630,N_4920,N_4464);
nor U5631 (N_5631,N_4143,N_4672);
nand U5632 (N_5632,N_4506,N_4268);
nor U5633 (N_5633,N_4140,N_4632);
or U5634 (N_5634,N_4244,N_4478);
nor U5635 (N_5635,N_4811,N_4375);
nor U5636 (N_5636,N_4665,N_4905);
nor U5637 (N_5637,N_4973,N_4763);
nand U5638 (N_5638,N_4018,N_4422);
nor U5639 (N_5639,N_4297,N_4574);
nand U5640 (N_5640,N_4121,N_4087);
and U5641 (N_5641,N_4926,N_4124);
or U5642 (N_5642,N_4645,N_4724);
nand U5643 (N_5643,N_4048,N_4258);
xor U5644 (N_5644,N_4632,N_4204);
and U5645 (N_5645,N_4871,N_4877);
nor U5646 (N_5646,N_4464,N_4104);
and U5647 (N_5647,N_4640,N_4453);
and U5648 (N_5648,N_4929,N_4723);
nor U5649 (N_5649,N_4658,N_4798);
or U5650 (N_5650,N_4943,N_4577);
or U5651 (N_5651,N_4725,N_4948);
or U5652 (N_5652,N_4402,N_4432);
and U5653 (N_5653,N_4467,N_4374);
xor U5654 (N_5654,N_4479,N_4752);
or U5655 (N_5655,N_4975,N_4281);
and U5656 (N_5656,N_4915,N_4983);
and U5657 (N_5657,N_4088,N_4652);
nand U5658 (N_5658,N_4922,N_4699);
nor U5659 (N_5659,N_4943,N_4428);
nor U5660 (N_5660,N_4509,N_4962);
or U5661 (N_5661,N_4993,N_4082);
and U5662 (N_5662,N_4298,N_4141);
and U5663 (N_5663,N_4805,N_4087);
or U5664 (N_5664,N_4350,N_4160);
nand U5665 (N_5665,N_4272,N_4879);
nand U5666 (N_5666,N_4567,N_4699);
nand U5667 (N_5667,N_4014,N_4165);
nand U5668 (N_5668,N_4395,N_4181);
nand U5669 (N_5669,N_4093,N_4117);
and U5670 (N_5670,N_4071,N_4776);
nand U5671 (N_5671,N_4613,N_4652);
or U5672 (N_5672,N_4386,N_4728);
and U5673 (N_5673,N_4184,N_4063);
nor U5674 (N_5674,N_4041,N_4366);
or U5675 (N_5675,N_4236,N_4850);
or U5676 (N_5676,N_4308,N_4159);
and U5677 (N_5677,N_4129,N_4759);
or U5678 (N_5678,N_4877,N_4130);
or U5679 (N_5679,N_4317,N_4718);
nand U5680 (N_5680,N_4365,N_4832);
and U5681 (N_5681,N_4149,N_4453);
nor U5682 (N_5682,N_4129,N_4212);
or U5683 (N_5683,N_4667,N_4483);
nand U5684 (N_5684,N_4825,N_4269);
and U5685 (N_5685,N_4400,N_4488);
and U5686 (N_5686,N_4836,N_4843);
and U5687 (N_5687,N_4037,N_4390);
and U5688 (N_5688,N_4825,N_4658);
or U5689 (N_5689,N_4918,N_4711);
and U5690 (N_5690,N_4264,N_4722);
and U5691 (N_5691,N_4618,N_4612);
and U5692 (N_5692,N_4923,N_4271);
nand U5693 (N_5693,N_4163,N_4129);
nor U5694 (N_5694,N_4019,N_4340);
nor U5695 (N_5695,N_4742,N_4560);
nand U5696 (N_5696,N_4051,N_4300);
and U5697 (N_5697,N_4254,N_4402);
and U5698 (N_5698,N_4014,N_4589);
or U5699 (N_5699,N_4733,N_4392);
nor U5700 (N_5700,N_4069,N_4263);
nand U5701 (N_5701,N_4437,N_4410);
nor U5702 (N_5702,N_4607,N_4896);
nand U5703 (N_5703,N_4212,N_4551);
nor U5704 (N_5704,N_4988,N_4989);
and U5705 (N_5705,N_4778,N_4232);
or U5706 (N_5706,N_4556,N_4712);
and U5707 (N_5707,N_4691,N_4587);
or U5708 (N_5708,N_4962,N_4948);
and U5709 (N_5709,N_4679,N_4089);
nor U5710 (N_5710,N_4869,N_4085);
nor U5711 (N_5711,N_4947,N_4769);
nor U5712 (N_5712,N_4443,N_4593);
or U5713 (N_5713,N_4023,N_4597);
and U5714 (N_5714,N_4546,N_4121);
or U5715 (N_5715,N_4542,N_4946);
nand U5716 (N_5716,N_4913,N_4653);
and U5717 (N_5717,N_4775,N_4952);
nor U5718 (N_5718,N_4921,N_4803);
and U5719 (N_5719,N_4710,N_4932);
or U5720 (N_5720,N_4422,N_4687);
or U5721 (N_5721,N_4473,N_4630);
and U5722 (N_5722,N_4856,N_4971);
nand U5723 (N_5723,N_4144,N_4771);
xor U5724 (N_5724,N_4193,N_4323);
or U5725 (N_5725,N_4203,N_4033);
nand U5726 (N_5726,N_4508,N_4581);
nand U5727 (N_5727,N_4848,N_4923);
xor U5728 (N_5728,N_4711,N_4259);
and U5729 (N_5729,N_4370,N_4212);
and U5730 (N_5730,N_4243,N_4796);
nor U5731 (N_5731,N_4848,N_4333);
nor U5732 (N_5732,N_4073,N_4401);
xor U5733 (N_5733,N_4771,N_4856);
nand U5734 (N_5734,N_4440,N_4815);
or U5735 (N_5735,N_4240,N_4171);
or U5736 (N_5736,N_4045,N_4185);
nand U5737 (N_5737,N_4004,N_4503);
nand U5738 (N_5738,N_4142,N_4006);
and U5739 (N_5739,N_4070,N_4263);
or U5740 (N_5740,N_4829,N_4408);
nor U5741 (N_5741,N_4799,N_4876);
nand U5742 (N_5742,N_4988,N_4530);
and U5743 (N_5743,N_4486,N_4844);
nand U5744 (N_5744,N_4671,N_4244);
and U5745 (N_5745,N_4189,N_4560);
and U5746 (N_5746,N_4512,N_4407);
or U5747 (N_5747,N_4022,N_4435);
nor U5748 (N_5748,N_4631,N_4730);
nor U5749 (N_5749,N_4275,N_4329);
nor U5750 (N_5750,N_4381,N_4855);
and U5751 (N_5751,N_4642,N_4799);
or U5752 (N_5752,N_4232,N_4498);
nor U5753 (N_5753,N_4373,N_4553);
and U5754 (N_5754,N_4859,N_4865);
nor U5755 (N_5755,N_4762,N_4664);
nor U5756 (N_5756,N_4191,N_4190);
and U5757 (N_5757,N_4588,N_4053);
or U5758 (N_5758,N_4520,N_4697);
or U5759 (N_5759,N_4340,N_4558);
and U5760 (N_5760,N_4928,N_4425);
or U5761 (N_5761,N_4579,N_4648);
nand U5762 (N_5762,N_4449,N_4265);
or U5763 (N_5763,N_4116,N_4057);
nand U5764 (N_5764,N_4517,N_4506);
and U5765 (N_5765,N_4971,N_4921);
or U5766 (N_5766,N_4019,N_4490);
nand U5767 (N_5767,N_4195,N_4550);
nor U5768 (N_5768,N_4857,N_4803);
or U5769 (N_5769,N_4203,N_4043);
nor U5770 (N_5770,N_4064,N_4548);
or U5771 (N_5771,N_4710,N_4430);
and U5772 (N_5772,N_4148,N_4413);
or U5773 (N_5773,N_4258,N_4892);
and U5774 (N_5774,N_4595,N_4238);
or U5775 (N_5775,N_4382,N_4171);
and U5776 (N_5776,N_4711,N_4250);
and U5777 (N_5777,N_4092,N_4393);
nor U5778 (N_5778,N_4323,N_4070);
or U5779 (N_5779,N_4580,N_4400);
nor U5780 (N_5780,N_4245,N_4280);
nand U5781 (N_5781,N_4748,N_4814);
nor U5782 (N_5782,N_4079,N_4868);
and U5783 (N_5783,N_4372,N_4511);
nor U5784 (N_5784,N_4539,N_4130);
nor U5785 (N_5785,N_4378,N_4286);
nand U5786 (N_5786,N_4725,N_4243);
or U5787 (N_5787,N_4173,N_4488);
and U5788 (N_5788,N_4327,N_4847);
nor U5789 (N_5789,N_4351,N_4234);
or U5790 (N_5790,N_4615,N_4492);
and U5791 (N_5791,N_4168,N_4404);
nand U5792 (N_5792,N_4112,N_4909);
or U5793 (N_5793,N_4740,N_4859);
nor U5794 (N_5794,N_4931,N_4873);
and U5795 (N_5795,N_4673,N_4313);
or U5796 (N_5796,N_4303,N_4527);
nand U5797 (N_5797,N_4199,N_4210);
nor U5798 (N_5798,N_4838,N_4331);
or U5799 (N_5799,N_4296,N_4482);
and U5800 (N_5800,N_4720,N_4171);
nand U5801 (N_5801,N_4318,N_4345);
and U5802 (N_5802,N_4880,N_4021);
or U5803 (N_5803,N_4667,N_4889);
nand U5804 (N_5804,N_4381,N_4257);
nor U5805 (N_5805,N_4321,N_4171);
nor U5806 (N_5806,N_4530,N_4768);
nand U5807 (N_5807,N_4724,N_4186);
nand U5808 (N_5808,N_4809,N_4211);
nor U5809 (N_5809,N_4692,N_4911);
or U5810 (N_5810,N_4443,N_4298);
nand U5811 (N_5811,N_4900,N_4436);
or U5812 (N_5812,N_4220,N_4297);
xor U5813 (N_5813,N_4770,N_4603);
nand U5814 (N_5814,N_4927,N_4608);
or U5815 (N_5815,N_4459,N_4452);
or U5816 (N_5816,N_4188,N_4880);
nand U5817 (N_5817,N_4069,N_4420);
or U5818 (N_5818,N_4800,N_4466);
or U5819 (N_5819,N_4506,N_4167);
or U5820 (N_5820,N_4845,N_4775);
and U5821 (N_5821,N_4720,N_4186);
or U5822 (N_5822,N_4379,N_4803);
nor U5823 (N_5823,N_4185,N_4094);
nor U5824 (N_5824,N_4694,N_4250);
or U5825 (N_5825,N_4403,N_4201);
nor U5826 (N_5826,N_4528,N_4556);
nand U5827 (N_5827,N_4634,N_4407);
or U5828 (N_5828,N_4500,N_4160);
or U5829 (N_5829,N_4034,N_4711);
or U5830 (N_5830,N_4888,N_4406);
and U5831 (N_5831,N_4330,N_4420);
nor U5832 (N_5832,N_4641,N_4506);
and U5833 (N_5833,N_4550,N_4686);
nand U5834 (N_5834,N_4323,N_4197);
nor U5835 (N_5835,N_4426,N_4410);
nand U5836 (N_5836,N_4992,N_4171);
nand U5837 (N_5837,N_4086,N_4338);
nor U5838 (N_5838,N_4093,N_4071);
or U5839 (N_5839,N_4607,N_4184);
or U5840 (N_5840,N_4946,N_4485);
nand U5841 (N_5841,N_4840,N_4014);
or U5842 (N_5842,N_4716,N_4158);
xnor U5843 (N_5843,N_4638,N_4090);
nor U5844 (N_5844,N_4203,N_4929);
and U5845 (N_5845,N_4430,N_4180);
or U5846 (N_5846,N_4218,N_4804);
or U5847 (N_5847,N_4610,N_4022);
and U5848 (N_5848,N_4097,N_4249);
and U5849 (N_5849,N_4951,N_4341);
nor U5850 (N_5850,N_4130,N_4804);
nand U5851 (N_5851,N_4082,N_4588);
xnor U5852 (N_5852,N_4510,N_4410);
xnor U5853 (N_5853,N_4240,N_4893);
or U5854 (N_5854,N_4421,N_4901);
nor U5855 (N_5855,N_4827,N_4650);
or U5856 (N_5856,N_4877,N_4566);
or U5857 (N_5857,N_4140,N_4764);
or U5858 (N_5858,N_4336,N_4747);
nand U5859 (N_5859,N_4058,N_4606);
nor U5860 (N_5860,N_4929,N_4704);
or U5861 (N_5861,N_4523,N_4616);
and U5862 (N_5862,N_4249,N_4687);
nand U5863 (N_5863,N_4949,N_4128);
or U5864 (N_5864,N_4879,N_4010);
nand U5865 (N_5865,N_4803,N_4653);
nand U5866 (N_5866,N_4229,N_4915);
and U5867 (N_5867,N_4745,N_4731);
or U5868 (N_5868,N_4576,N_4627);
nor U5869 (N_5869,N_4365,N_4750);
nor U5870 (N_5870,N_4865,N_4737);
and U5871 (N_5871,N_4964,N_4461);
or U5872 (N_5872,N_4375,N_4294);
or U5873 (N_5873,N_4035,N_4047);
nand U5874 (N_5874,N_4497,N_4974);
and U5875 (N_5875,N_4115,N_4980);
nand U5876 (N_5876,N_4139,N_4251);
nor U5877 (N_5877,N_4595,N_4543);
nor U5878 (N_5878,N_4954,N_4226);
or U5879 (N_5879,N_4659,N_4358);
xnor U5880 (N_5880,N_4774,N_4749);
nor U5881 (N_5881,N_4247,N_4528);
nor U5882 (N_5882,N_4114,N_4425);
and U5883 (N_5883,N_4358,N_4484);
or U5884 (N_5884,N_4280,N_4295);
nor U5885 (N_5885,N_4269,N_4830);
nor U5886 (N_5886,N_4334,N_4609);
nand U5887 (N_5887,N_4237,N_4777);
and U5888 (N_5888,N_4648,N_4846);
nor U5889 (N_5889,N_4124,N_4982);
nand U5890 (N_5890,N_4854,N_4466);
nand U5891 (N_5891,N_4339,N_4999);
or U5892 (N_5892,N_4542,N_4438);
or U5893 (N_5893,N_4394,N_4997);
nor U5894 (N_5894,N_4797,N_4507);
and U5895 (N_5895,N_4988,N_4611);
nand U5896 (N_5896,N_4401,N_4092);
nand U5897 (N_5897,N_4605,N_4244);
nor U5898 (N_5898,N_4683,N_4822);
and U5899 (N_5899,N_4287,N_4765);
and U5900 (N_5900,N_4179,N_4619);
or U5901 (N_5901,N_4610,N_4390);
nor U5902 (N_5902,N_4651,N_4551);
or U5903 (N_5903,N_4152,N_4491);
nor U5904 (N_5904,N_4184,N_4029);
and U5905 (N_5905,N_4250,N_4972);
or U5906 (N_5906,N_4917,N_4407);
or U5907 (N_5907,N_4458,N_4049);
and U5908 (N_5908,N_4334,N_4491);
or U5909 (N_5909,N_4143,N_4854);
or U5910 (N_5910,N_4161,N_4222);
or U5911 (N_5911,N_4796,N_4836);
or U5912 (N_5912,N_4462,N_4227);
or U5913 (N_5913,N_4337,N_4892);
or U5914 (N_5914,N_4599,N_4651);
or U5915 (N_5915,N_4278,N_4951);
nor U5916 (N_5916,N_4204,N_4586);
and U5917 (N_5917,N_4901,N_4281);
and U5918 (N_5918,N_4527,N_4741);
and U5919 (N_5919,N_4605,N_4076);
and U5920 (N_5920,N_4915,N_4685);
nor U5921 (N_5921,N_4854,N_4013);
nand U5922 (N_5922,N_4004,N_4901);
or U5923 (N_5923,N_4875,N_4592);
or U5924 (N_5924,N_4590,N_4190);
and U5925 (N_5925,N_4331,N_4306);
and U5926 (N_5926,N_4765,N_4649);
nand U5927 (N_5927,N_4000,N_4507);
nand U5928 (N_5928,N_4225,N_4565);
nand U5929 (N_5929,N_4459,N_4017);
or U5930 (N_5930,N_4282,N_4661);
nand U5931 (N_5931,N_4202,N_4898);
or U5932 (N_5932,N_4685,N_4713);
or U5933 (N_5933,N_4946,N_4065);
nor U5934 (N_5934,N_4550,N_4965);
and U5935 (N_5935,N_4172,N_4066);
and U5936 (N_5936,N_4701,N_4201);
nand U5937 (N_5937,N_4602,N_4676);
or U5938 (N_5938,N_4161,N_4424);
or U5939 (N_5939,N_4414,N_4943);
nand U5940 (N_5940,N_4904,N_4315);
xnor U5941 (N_5941,N_4299,N_4510);
and U5942 (N_5942,N_4567,N_4045);
nand U5943 (N_5943,N_4647,N_4067);
and U5944 (N_5944,N_4899,N_4873);
or U5945 (N_5945,N_4034,N_4391);
and U5946 (N_5946,N_4897,N_4221);
nand U5947 (N_5947,N_4866,N_4184);
or U5948 (N_5948,N_4905,N_4061);
nor U5949 (N_5949,N_4815,N_4044);
or U5950 (N_5950,N_4583,N_4770);
or U5951 (N_5951,N_4893,N_4841);
and U5952 (N_5952,N_4104,N_4482);
or U5953 (N_5953,N_4476,N_4636);
nor U5954 (N_5954,N_4671,N_4031);
or U5955 (N_5955,N_4508,N_4512);
and U5956 (N_5956,N_4702,N_4044);
nor U5957 (N_5957,N_4516,N_4206);
nand U5958 (N_5958,N_4521,N_4855);
or U5959 (N_5959,N_4526,N_4197);
or U5960 (N_5960,N_4247,N_4402);
nor U5961 (N_5961,N_4164,N_4574);
nor U5962 (N_5962,N_4439,N_4393);
and U5963 (N_5963,N_4624,N_4851);
and U5964 (N_5964,N_4207,N_4972);
nand U5965 (N_5965,N_4626,N_4829);
and U5966 (N_5966,N_4637,N_4594);
or U5967 (N_5967,N_4759,N_4411);
nand U5968 (N_5968,N_4776,N_4059);
or U5969 (N_5969,N_4204,N_4877);
nor U5970 (N_5970,N_4221,N_4576);
nor U5971 (N_5971,N_4047,N_4530);
or U5972 (N_5972,N_4008,N_4320);
nand U5973 (N_5973,N_4106,N_4905);
or U5974 (N_5974,N_4828,N_4813);
and U5975 (N_5975,N_4563,N_4719);
nand U5976 (N_5976,N_4490,N_4571);
and U5977 (N_5977,N_4346,N_4226);
nor U5978 (N_5978,N_4394,N_4544);
and U5979 (N_5979,N_4255,N_4241);
nand U5980 (N_5980,N_4804,N_4751);
nor U5981 (N_5981,N_4849,N_4026);
and U5982 (N_5982,N_4159,N_4230);
and U5983 (N_5983,N_4220,N_4004);
and U5984 (N_5984,N_4239,N_4673);
nor U5985 (N_5985,N_4615,N_4486);
nor U5986 (N_5986,N_4808,N_4013);
nor U5987 (N_5987,N_4998,N_4138);
or U5988 (N_5988,N_4669,N_4047);
xor U5989 (N_5989,N_4865,N_4346);
nor U5990 (N_5990,N_4123,N_4368);
nor U5991 (N_5991,N_4209,N_4251);
nand U5992 (N_5992,N_4394,N_4677);
or U5993 (N_5993,N_4807,N_4113);
nor U5994 (N_5994,N_4639,N_4139);
nor U5995 (N_5995,N_4415,N_4165);
and U5996 (N_5996,N_4961,N_4167);
nand U5997 (N_5997,N_4022,N_4492);
and U5998 (N_5998,N_4654,N_4373);
nand U5999 (N_5999,N_4013,N_4294);
or U6000 (N_6000,N_5272,N_5012);
and U6001 (N_6001,N_5350,N_5660);
nor U6002 (N_6002,N_5924,N_5200);
nor U6003 (N_6003,N_5715,N_5850);
nand U6004 (N_6004,N_5489,N_5337);
or U6005 (N_6005,N_5655,N_5956);
or U6006 (N_6006,N_5409,N_5454);
or U6007 (N_6007,N_5895,N_5885);
and U6008 (N_6008,N_5762,N_5898);
and U6009 (N_6009,N_5801,N_5434);
nor U6010 (N_6010,N_5168,N_5731);
nor U6011 (N_6011,N_5056,N_5998);
nor U6012 (N_6012,N_5349,N_5439);
and U6013 (N_6013,N_5588,N_5061);
nand U6014 (N_6014,N_5029,N_5468);
nor U6015 (N_6015,N_5965,N_5093);
nand U6016 (N_6016,N_5204,N_5065);
and U6017 (N_6017,N_5685,N_5818);
nand U6018 (N_6018,N_5481,N_5677);
and U6019 (N_6019,N_5743,N_5985);
or U6020 (N_6020,N_5907,N_5375);
nand U6021 (N_6021,N_5530,N_5886);
nand U6022 (N_6022,N_5329,N_5799);
nand U6023 (N_6023,N_5425,N_5193);
or U6024 (N_6024,N_5797,N_5086);
and U6025 (N_6025,N_5559,N_5458);
and U6026 (N_6026,N_5927,N_5922);
and U6027 (N_6027,N_5037,N_5054);
nor U6028 (N_6028,N_5158,N_5095);
nor U6029 (N_6029,N_5150,N_5900);
and U6030 (N_6030,N_5803,N_5394);
or U6031 (N_6031,N_5014,N_5167);
nor U6032 (N_6032,N_5978,N_5858);
or U6033 (N_6033,N_5546,N_5007);
and U6034 (N_6034,N_5179,N_5804);
or U6035 (N_6035,N_5328,N_5967);
and U6036 (N_6036,N_5631,N_5341);
or U6037 (N_6037,N_5739,N_5210);
xor U6038 (N_6038,N_5391,N_5909);
or U6039 (N_6039,N_5059,N_5115);
and U6040 (N_6040,N_5820,N_5396);
and U6041 (N_6041,N_5825,N_5628);
nand U6042 (N_6042,N_5526,N_5064);
and U6043 (N_6043,N_5157,N_5625);
nor U6044 (N_6044,N_5618,N_5240);
nand U6045 (N_6045,N_5867,N_5979);
and U6046 (N_6046,N_5791,N_5138);
and U6047 (N_6047,N_5494,N_5667);
or U6048 (N_6048,N_5925,N_5194);
nand U6049 (N_6049,N_5798,N_5902);
and U6050 (N_6050,N_5950,N_5321);
and U6051 (N_6051,N_5078,N_5892);
nor U6052 (N_6052,N_5835,N_5219);
nor U6053 (N_6053,N_5683,N_5433);
or U6054 (N_6054,N_5670,N_5103);
and U6055 (N_6055,N_5497,N_5897);
xnor U6056 (N_6056,N_5241,N_5876);
nor U6057 (N_6057,N_5044,N_5399);
nor U6058 (N_6058,N_5267,N_5230);
or U6059 (N_6059,N_5148,N_5424);
and U6060 (N_6060,N_5675,N_5878);
nor U6061 (N_6061,N_5414,N_5382);
and U6062 (N_6062,N_5624,N_5453);
nor U6063 (N_6063,N_5912,N_5383);
nor U6064 (N_6064,N_5969,N_5948);
nor U6065 (N_6065,N_5988,N_5020);
nand U6066 (N_6066,N_5510,N_5034);
nor U6067 (N_6067,N_5750,N_5567);
nor U6068 (N_6068,N_5451,N_5467);
and U6069 (N_6069,N_5543,N_5827);
nor U6070 (N_6070,N_5006,N_5852);
and U6071 (N_6071,N_5268,N_5342);
or U6072 (N_6072,N_5218,N_5916);
or U6073 (N_6073,N_5220,N_5380);
nor U6074 (N_6074,N_5700,N_5811);
nor U6075 (N_6075,N_5822,N_5785);
and U6076 (N_6076,N_5865,N_5203);
nand U6077 (N_6077,N_5903,N_5857);
or U6078 (N_6078,N_5122,N_5493);
nand U6079 (N_6079,N_5788,N_5830);
or U6080 (N_6080,N_5415,N_5197);
nand U6081 (N_6081,N_5163,N_5478);
or U6082 (N_6082,N_5263,N_5066);
nand U6083 (N_6083,N_5420,N_5609);
nor U6084 (N_6084,N_5590,N_5226);
nand U6085 (N_6085,N_5067,N_5513);
or U6086 (N_6086,N_5110,N_5235);
and U6087 (N_6087,N_5643,N_5090);
and U6088 (N_6088,N_5534,N_5834);
nor U6089 (N_6089,N_5854,N_5695);
nand U6090 (N_6090,N_5792,N_5484);
and U6091 (N_6091,N_5701,N_5175);
nand U6092 (N_6092,N_5729,N_5404);
nor U6093 (N_6093,N_5509,N_5351);
or U6094 (N_6094,N_5340,N_5612);
and U6095 (N_6095,N_5836,N_5547);
or U6096 (N_6096,N_5536,N_5072);
nand U6097 (N_6097,N_5352,N_5908);
nor U6098 (N_6098,N_5302,N_5046);
or U6099 (N_6099,N_5395,N_5958);
and U6100 (N_6100,N_5918,N_5787);
and U6101 (N_6101,N_5173,N_5233);
and U6102 (N_6102,N_5053,N_5275);
or U6103 (N_6103,N_5953,N_5725);
nand U6104 (N_6104,N_5539,N_5440);
nor U6105 (N_6105,N_5594,N_5027);
or U6106 (N_6106,N_5309,N_5511);
or U6107 (N_6107,N_5455,N_5605);
and U6108 (N_6108,N_5097,N_5705);
nor U6109 (N_6109,N_5068,N_5370);
nand U6110 (N_6110,N_5627,N_5418);
or U6111 (N_6111,N_5602,N_5744);
nor U6112 (N_6112,N_5401,N_5585);
nand U6113 (N_6113,N_5776,N_5595);
xnor U6114 (N_6114,N_5741,N_5472);
nor U6115 (N_6115,N_5707,N_5149);
and U6116 (N_6116,N_5664,N_5055);
nor U6117 (N_6117,N_5023,N_5751);
or U6118 (N_6118,N_5291,N_5764);
or U6119 (N_6119,N_5265,N_5807);
or U6120 (N_6120,N_5809,N_5782);
or U6121 (N_6121,N_5123,N_5459);
nand U6122 (N_6122,N_5698,N_5819);
xor U6123 (N_6123,N_5155,N_5249);
nand U6124 (N_6124,N_5336,N_5199);
nor U6125 (N_6125,N_5102,N_5773);
or U6126 (N_6126,N_5413,N_5877);
and U6127 (N_6127,N_5222,N_5506);
nand U6128 (N_6128,N_5768,N_5777);
and U6129 (N_6129,N_5558,N_5284);
nor U6130 (N_6130,N_5889,N_5929);
and U6131 (N_6131,N_5737,N_5471);
nand U6132 (N_6132,N_5507,N_5862);
or U6133 (N_6133,N_5607,N_5362);
nand U6134 (N_6134,N_5151,N_5369);
or U6135 (N_6135,N_5180,N_5872);
nand U6136 (N_6136,N_5614,N_5621);
nand U6137 (N_6137,N_5673,N_5243);
nor U6138 (N_6138,N_5174,N_5063);
nand U6139 (N_6139,N_5774,N_5699);
or U6140 (N_6140,N_5575,N_5079);
nor U6141 (N_6141,N_5320,N_5390);
or U6142 (N_6142,N_5091,N_5387);
nor U6143 (N_6143,N_5429,N_5718);
nor U6144 (N_6144,N_5997,N_5719);
or U6145 (N_6145,N_5160,N_5146);
or U6146 (N_6146,N_5659,N_5231);
and U6147 (N_6147,N_5278,N_5738);
nor U6148 (N_6148,N_5264,N_5448);
or U6149 (N_6149,N_5600,N_5665);
and U6150 (N_6150,N_5361,N_5554);
nand U6151 (N_6151,N_5931,N_5951);
nor U6152 (N_6152,N_5080,N_5704);
nand U6153 (N_6153,N_5645,N_5623);
and U6154 (N_6154,N_5247,N_5295);
nand U6155 (N_6155,N_5790,N_5153);
nand U6156 (N_6156,N_5259,N_5388);
or U6157 (N_6157,N_5863,N_5565);
or U6158 (N_6158,N_5270,N_5474);
or U6159 (N_6159,N_5255,N_5552);
nor U6160 (N_6160,N_5649,N_5205);
nand U6161 (N_6161,N_5887,N_5528);
nor U6162 (N_6162,N_5315,N_5195);
nor U6163 (N_6163,N_5873,N_5587);
and U6164 (N_6164,N_5124,N_5300);
and U6165 (N_6165,N_5058,N_5374);
nor U6166 (N_6166,N_5734,N_5540);
nand U6167 (N_6167,N_5282,N_5299);
nor U6168 (N_6168,N_5775,N_5533);
nand U6169 (N_6169,N_5288,N_5217);
and U6170 (N_6170,N_5982,N_5136);
nor U6171 (N_6171,N_5561,N_5723);
or U6172 (N_6172,N_5444,N_5947);
and U6173 (N_6173,N_5470,N_5116);
and U6174 (N_6174,N_5626,N_5426);
or U6175 (N_6175,N_5457,N_5682);
or U6176 (N_6176,N_5258,N_5227);
or U6177 (N_6177,N_5347,N_5129);
and U6178 (N_6178,N_5893,N_5469);
and U6179 (N_6179,N_5112,N_5154);
nor U6180 (N_6180,N_5159,N_5672);
or U6181 (N_6181,N_5488,N_5518);
or U6182 (N_6182,N_5652,N_5579);
nor U6183 (N_6183,N_5962,N_5441);
nand U6184 (N_6184,N_5745,N_5514);
or U6185 (N_6185,N_5896,N_5688);
or U6186 (N_6186,N_5742,N_5573);
or U6187 (N_6187,N_5525,N_5169);
or U6188 (N_6188,N_5304,N_5188);
and U6189 (N_6189,N_5131,N_5772);
nor U6190 (N_6190,N_5324,N_5646);
nand U6191 (N_6191,N_5901,N_5726);
or U6192 (N_6192,N_5991,N_5201);
nor U6193 (N_6193,N_5608,N_5339);
nand U6194 (N_6194,N_5757,N_5187);
and U6195 (N_6195,N_5717,N_5890);
or U6196 (N_6196,N_5164,N_5832);
nand U6197 (N_6197,N_5606,N_5465);
or U6198 (N_6198,N_5040,N_5856);
or U6199 (N_6199,N_5844,N_5244);
or U6200 (N_6200,N_5177,N_5689);
nand U6201 (N_6201,N_5431,N_5557);
or U6202 (N_6202,N_5353,N_5030);
nor U6203 (N_6203,N_5330,N_5373);
nand U6204 (N_6204,N_5538,N_5117);
and U6205 (N_6205,N_5582,N_5276);
nor U6206 (N_6206,N_5555,N_5196);
and U6207 (N_6207,N_5580,N_5930);
and U6208 (N_6208,N_5941,N_5301);
and U6209 (N_6209,N_5333,N_5516);
nand U6210 (N_6210,N_5716,N_5476);
nor U6211 (N_6211,N_5041,N_5008);
or U6212 (N_6212,N_5911,N_5833);
nor U6213 (N_6213,N_5831,N_5126);
and U6214 (N_6214,N_5935,N_5944);
or U6215 (N_6215,N_5297,N_5307);
nand U6216 (N_6216,N_5566,N_5814);
nand U6217 (N_6217,N_5840,N_5118);
nand U6218 (N_6218,N_5989,N_5239);
nand U6219 (N_6219,N_5428,N_5313);
or U6220 (N_6220,N_5636,N_5142);
xor U6221 (N_6221,N_5132,N_5881);
nand U6222 (N_6222,N_5882,N_5372);
nor U6223 (N_6223,N_5823,N_5905);
and U6224 (N_6224,N_5505,N_5245);
nand U6225 (N_6225,N_5871,N_5828);
nor U6226 (N_6226,N_5043,N_5974);
nor U6227 (N_6227,N_5593,N_5613);
xor U6228 (N_6228,N_5868,N_5225);
and U6229 (N_6229,N_5971,N_5326);
and U6230 (N_6230,N_5562,N_5162);
nand U6231 (N_6231,N_5325,N_5855);
and U6232 (N_6232,N_5592,N_5308);
and U6233 (N_6233,N_5354,N_5416);
nand U6234 (N_6234,N_5100,N_5691);
nor U6235 (N_6235,N_5371,N_5793);
nor U6236 (N_6236,N_5815,N_5954);
or U6237 (N_6237,N_5316,N_5121);
or U6238 (N_6238,N_5894,N_5541);
or U6239 (N_6239,N_5487,N_5730);
or U6240 (N_6240,N_5501,N_5763);
nand U6241 (N_6241,N_5161,N_5386);
nand U6242 (N_6242,N_5586,N_5632);
nand U6243 (N_6243,N_5917,N_5109);
or U6244 (N_6244,N_5687,N_5224);
nor U6245 (N_6245,N_5708,N_5026);
or U6246 (N_6246,N_5570,N_5410);
and U6247 (N_6247,N_5702,N_5760);
nand U6248 (N_6248,N_5517,N_5943);
and U6249 (N_6249,N_5223,N_5498);
nand U6250 (N_6250,N_5190,N_5732);
or U6251 (N_6251,N_5666,N_5789);
and U6252 (N_6252,N_5746,N_5955);
nand U6253 (N_6253,N_5111,N_5283);
or U6254 (N_6254,N_5145,N_5527);
nand U6255 (N_6255,N_5523,N_5186);
nor U6256 (N_6256,N_5092,N_5460);
nand U6257 (N_6257,N_5213,N_5492);
and U6258 (N_6258,N_5082,N_5359);
and U6259 (N_6259,N_5904,N_5860);
nand U6260 (N_6260,N_5128,N_5826);
nor U6261 (N_6261,N_5071,N_5601);
nor U6262 (N_6262,N_5697,N_5398);
or U6263 (N_6263,N_5089,N_5211);
nand U6264 (N_6264,N_5994,N_5192);
and U6265 (N_6265,N_5345,N_5537);
nand U6266 (N_6266,N_5479,N_5520);
or U6267 (N_6267,N_5464,N_5269);
and U6268 (N_6268,N_5846,N_5942);
or U6269 (N_6269,N_5678,N_5630);
and U6270 (N_6270,N_5057,N_5266);
nor U6271 (N_6271,N_5843,N_5692);
nand U6272 (N_6272,N_5781,N_5368);
nand U6273 (N_6273,N_5004,N_5417);
or U6274 (N_6274,N_5019,N_5668);
nor U6275 (N_6275,N_5294,N_5170);
or U6276 (N_6276,N_5946,N_5812);
nand U6277 (N_6277,N_5839,N_5183);
and U6278 (N_6278,N_5184,N_5237);
nand U6279 (N_6279,N_5796,N_5456);
xnor U6280 (N_6280,N_5419,N_5710);
and U6281 (N_6281,N_5038,N_5310);
nor U6282 (N_6282,N_5544,N_5611);
nor U6283 (N_6283,N_5133,N_5049);
nor U6284 (N_6284,N_5740,N_5591);
nand U6285 (N_6285,N_5770,N_5752);
or U6286 (N_6286,N_5077,N_5490);
nand U6287 (N_6287,N_5845,N_5654);
or U6288 (N_6288,N_5025,N_5619);
nor U6289 (N_6289,N_5135,N_5713);
or U6290 (N_6290,N_5005,N_5550);
nor U6291 (N_6291,N_5615,N_5436);
and U6292 (N_6292,N_5913,N_5759);
xnor U6293 (N_6293,N_5771,N_5553);
and U6294 (N_6294,N_5721,N_5966);
or U6295 (N_6295,N_5191,N_5393);
and U6296 (N_6296,N_5859,N_5888);
and U6297 (N_6297,N_5273,N_5577);
and U6298 (N_6298,N_5596,N_5604);
or U6299 (N_6299,N_5281,N_5015);
nand U6300 (N_6300,N_5334,N_5599);
nor U6301 (N_6301,N_5661,N_5031);
and U6302 (N_6302,N_5178,N_5018);
or U6303 (N_6303,N_5576,N_5322);
nor U6304 (N_6304,N_5366,N_5084);
nand U6305 (N_6305,N_5870,N_5016);
and U6306 (N_6306,N_5290,N_5296);
or U6307 (N_6307,N_5069,N_5920);
nor U6308 (N_6308,N_5070,N_5853);
or U6309 (N_6309,N_5589,N_5246);
or U6310 (N_6310,N_5216,N_5653);
nor U6311 (N_6311,N_5945,N_5292);
nand U6312 (N_6312,N_5319,N_5363);
and U6313 (N_6313,N_5221,N_5634);
and U6314 (N_6314,N_5332,N_5254);
xnor U6315 (N_6315,N_5480,N_5389);
and U6316 (N_6316,N_5022,N_5551);
nand U6317 (N_6317,N_5185,N_5344);
nand U6318 (N_6318,N_5094,N_5957);
nand U6319 (N_6319,N_5684,N_5849);
nor U6320 (N_6320,N_5817,N_5262);
and U6321 (N_6321,N_5314,N_5009);
nand U6322 (N_6322,N_5141,N_5786);
xor U6323 (N_6323,N_5829,N_5236);
nand U6324 (N_6324,N_5001,N_5838);
nand U6325 (N_6325,N_5081,N_5800);
and U6326 (N_6326,N_5866,N_5143);
nor U6327 (N_6327,N_5584,N_5984);
nor U6328 (N_6328,N_5769,N_5209);
and U6329 (N_6329,N_5364,N_5202);
or U6330 (N_6330,N_5560,N_5610);
nand U6331 (N_6331,N_5156,N_5252);
nor U6332 (N_6332,N_5676,N_5648);
and U6333 (N_6333,N_5357,N_5408);
or U6334 (N_6334,N_5039,N_5317);
nand U6335 (N_6335,N_5542,N_5977);
nand U6336 (N_6336,N_5432,N_5712);
nand U6337 (N_6337,N_5189,N_5635);
and U6338 (N_6338,N_5050,N_5709);
nor U6339 (N_6339,N_5442,N_5842);
or U6340 (N_6340,N_5172,N_5808);
nor U6341 (N_6341,N_5435,N_5411);
or U6342 (N_6342,N_5761,N_5564);
nor U6343 (N_6343,N_5011,N_5312);
or U6344 (N_6344,N_5208,N_5932);
nand U6345 (N_6345,N_5983,N_5139);
and U6346 (N_6346,N_5215,N_5921);
nor U6347 (N_6347,N_5392,N_5075);
or U6348 (N_6348,N_5311,N_5503);
nand U6349 (N_6349,N_5754,N_5597);
nor U6350 (N_6350,N_5271,N_5358);
and U6351 (N_6351,N_5406,N_5622);
xor U6352 (N_6352,N_5412,N_5473);
nor U6353 (N_6353,N_5238,N_5140);
nand U6354 (N_6354,N_5171,N_5884);
and U6355 (N_6355,N_5105,N_5214);
nand U6356 (N_6356,N_5286,N_5937);
or U6357 (N_6357,N_5874,N_5035);
nand U6358 (N_6358,N_5674,N_5348);
or U6359 (N_6359,N_5360,N_5995);
nor U6360 (N_6360,N_5335,N_5466);
or U6361 (N_6361,N_5166,N_5934);
or U6362 (N_6362,N_5926,N_5073);
or U6363 (N_6363,N_5783,N_5650);
nor U6364 (N_6364,N_5234,N_5365);
and U6365 (N_6365,N_5475,N_5367);
nand U6366 (N_6366,N_5959,N_5280);
nor U6367 (N_6367,N_5229,N_5861);
nand U6368 (N_6368,N_5722,N_5658);
nor U6369 (N_6369,N_5747,N_5960);
or U6370 (N_6370,N_5875,N_5879);
nor U6371 (N_6371,N_5690,N_5671);
and U6372 (N_6372,N_5651,N_5108);
or U6373 (N_6373,N_5724,N_5021);
and U6374 (N_6374,N_5938,N_5500);
nor U6375 (N_6375,N_5134,N_5285);
nor U6376 (N_6376,N_5165,N_5933);
and U6377 (N_6377,N_5101,N_5765);
and U6378 (N_6378,N_5794,N_5640);
nand U6379 (N_6379,N_5563,N_5421);
nor U6380 (N_6380,N_5638,N_5795);
nand U6381 (N_6381,N_5633,N_5923);
or U6382 (N_6382,N_5125,N_5293);
and U6383 (N_6383,N_5515,N_5405);
nor U6384 (N_6384,N_5970,N_5806);
and U6385 (N_6385,N_5107,N_5438);
nand U6386 (N_6386,N_5512,N_5574);
nor U6387 (N_6387,N_5940,N_5848);
nor U6388 (N_6388,N_5629,N_5706);
or U6389 (N_6389,N_5376,N_5976);
and U6390 (N_6390,N_5104,N_5728);
nor U6391 (N_6391,N_5961,N_5910);
and U6392 (N_6392,N_5378,N_5987);
and U6393 (N_6393,N_5096,N_5346);
nor U6394 (N_6394,N_5338,N_5711);
nand U6395 (N_6395,N_5990,N_5805);
or U6396 (N_6396,N_5379,N_5549);
and U6397 (N_6397,N_5381,N_5445);
nand U6398 (N_6398,N_5569,N_5568);
nand U6399 (N_6399,N_5522,N_5919);
nand U6400 (N_6400,N_5486,N_5703);
and U6401 (N_6401,N_5578,N_5013);
nor U6402 (N_6402,N_5450,N_5869);
or U6403 (N_6403,N_5972,N_5062);
and U6404 (N_6404,N_5355,N_5696);
nand U6405 (N_6405,N_5289,N_5099);
and U6406 (N_6406,N_5813,N_5051);
or U6407 (N_6407,N_5641,N_5647);
nor U6408 (N_6408,N_5083,N_5686);
and U6409 (N_6409,N_5485,N_5356);
nand U6410 (N_6410,N_5242,N_5727);
xor U6411 (N_6411,N_5531,N_5694);
or U6412 (N_6412,N_5212,N_5810);
nor U6413 (N_6413,N_5274,N_5250);
nand U6414 (N_6414,N_5519,N_5403);
nand U6415 (N_6415,N_5427,N_5137);
nor U6416 (N_6416,N_5087,N_5571);
and U6417 (N_6417,N_5939,N_5644);
xor U6418 (N_6418,N_5060,N_5402);
nand U6419 (N_6419,N_5508,N_5257);
and U6420 (N_6420,N_5261,N_5603);
and U6421 (N_6421,N_5847,N_5993);
and U6422 (N_6422,N_5656,N_5028);
and U6423 (N_6423,N_5986,N_5524);
and U6424 (N_6424,N_5521,N_5074);
and U6425 (N_6425,N_5598,N_5120);
and U6426 (N_6426,N_5113,N_5767);
and U6427 (N_6427,N_5864,N_5779);
nand U6428 (N_6428,N_5837,N_5377);
or U6429 (N_6429,N_5446,N_5277);
nor U6430 (N_6430,N_5980,N_5251);
or U6431 (N_6431,N_5581,N_5130);
nand U6432 (N_6432,N_5891,N_5152);
or U6433 (N_6433,N_5407,N_5327);
xor U6434 (N_6434,N_5663,N_5949);
xor U6435 (N_6435,N_5232,N_5915);
nor U6436 (N_6436,N_5303,N_5981);
and U6437 (N_6437,N_5447,N_5318);
or U6438 (N_6438,N_5642,N_5298);
or U6439 (N_6439,N_5323,N_5748);
or U6440 (N_6440,N_5914,N_5483);
nand U6441 (N_6441,N_5545,N_5975);
and U6442 (N_6442,N_5106,N_5529);
nor U6443 (N_6443,N_5749,N_5936);
nor U6444 (N_6444,N_5182,N_5422);
and U6445 (N_6445,N_5256,N_5906);
and U6446 (N_6446,N_5778,N_5000);
or U6447 (N_6447,N_5952,N_5802);
or U6448 (N_6448,N_5088,N_5693);
nor U6449 (N_6449,N_5010,N_5400);
nor U6450 (N_6450,N_5824,N_5755);
nor U6451 (N_6451,N_5669,N_5502);
or U6452 (N_6452,N_5287,N_5461);
and U6453 (N_6453,N_5033,N_5657);
nor U6454 (N_6454,N_5964,N_5076);
or U6455 (N_6455,N_5114,N_5821);
or U6456 (N_6456,N_5181,N_5639);
nor U6457 (N_6457,N_5883,N_5780);
and U6458 (N_6458,N_5504,N_5766);
nor U6459 (N_6459,N_5532,N_5462);
or U6460 (N_6460,N_5996,N_5968);
and U6461 (N_6461,N_5583,N_5085);
or U6462 (N_6462,N_5127,N_5616);
xnor U6463 (N_6463,N_5198,N_5999);
nor U6464 (N_6464,N_5963,N_5880);
nor U6465 (N_6465,N_5680,N_5003);
nand U6466 (N_6466,N_5207,N_5397);
nand U6467 (N_6467,N_5098,N_5343);
or U6468 (N_6468,N_5305,N_5206);
nand U6469 (N_6469,N_5253,N_5851);
xor U6470 (N_6470,N_5758,N_5248);
nand U6471 (N_6471,N_5681,N_5032);
nor U6472 (N_6472,N_5384,N_5548);
or U6473 (N_6473,N_5714,N_5176);
xor U6474 (N_6474,N_5385,N_5042);
nand U6475 (N_6475,N_5992,N_5620);
or U6476 (N_6476,N_5260,N_5449);
nor U6477 (N_6477,N_5662,N_5899);
or U6478 (N_6478,N_5784,N_5482);
nor U6479 (N_6479,N_5753,N_5228);
nor U6480 (N_6480,N_5017,N_5720);
nor U6481 (N_6481,N_5452,N_5279);
nor U6482 (N_6482,N_5443,N_5556);
or U6483 (N_6483,N_5119,N_5572);
nand U6484 (N_6484,N_5841,N_5437);
or U6485 (N_6485,N_5045,N_5052);
nor U6486 (N_6486,N_5973,N_5816);
and U6487 (N_6487,N_5499,N_5430);
nor U6488 (N_6488,N_5002,N_5736);
and U6489 (N_6489,N_5679,N_5756);
nor U6490 (N_6490,N_5928,N_5144);
or U6491 (N_6491,N_5496,N_5047);
or U6492 (N_6492,N_5463,N_5617);
nand U6493 (N_6493,N_5535,N_5423);
nor U6494 (N_6494,N_5036,N_5331);
nor U6495 (N_6495,N_5048,N_5147);
or U6496 (N_6496,N_5477,N_5495);
and U6497 (N_6497,N_5024,N_5735);
and U6498 (N_6498,N_5306,N_5733);
or U6499 (N_6499,N_5637,N_5491);
nor U6500 (N_6500,N_5002,N_5984);
and U6501 (N_6501,N_5184,N_5518);
and U6502 (N_6502,N_5863,N_5505);
and U6503 (N_6503,N_5048,N_5702);
xor U6504 (N_6504,N_5941,N_5700);
or U6505 (N_6505,N_5030,N_5099);
or U6506 (N_6506,N_5905,N_5387);
nand U6507 (N_6507,N_5018,N_5834);
nor U6508 (N_6508,N_5608,N_5811);
or U6509 (N_6509,N_5988,N_5637);
or U6510 (N_6510,N_5626,N_5888);
or U6511 (N_6511,N_5983,N_5309);
and U6512 (N_6512,N_5962,N_5260);
nor U6513 (N_6513,N_5797,N_5785);
and U6514 (N_6514,N_5790,N_5556);
or U6515 (N_6515,N_5947,N_5984);
nand U6516 (N_6516,N_5522,N_5675);
nand U6517 (N_6517,N_5143,N_5506);
or U6518 (N_6518,N_5971,N_5567);
and U6519 (N_6519,N_5717,N_5954);
nand U6520 (N_6520,N_5589,N_5617);
and U6521 (N_6521,N_5325,N_5349);
nand U6522 (N_6522,N_5889,N_5400);
nand U6523 (N_6523,N_5093,N_5396);
and U6524 (N_6524,N_5268,N_5571);
and U6525 (N_6525,N_5004,N_5891);
xnor U6526 (N_6526,N_5518,N_5988);
and U6527 (N_6527,N_5348,N_5924);
nand U6528 (N_6528,N_5739,N_5379);
nand U6529 (N_6529,N_5260,N_5385);
and U6530 (N_6530,N_5936,N_5280);
nand U6531 (N_6531,N_5121,N_5243);
nor U6532 (N_6532,N_5979,N_5776);
nand U6533 (N_6533,N_5091,N_5123);
nand U6534 (N_6534,N_5235,N_5257);
xnor U6535 (N_6535,N_5365,N_5052);
nand U6536 (N_6536,N_5884,N_5905);
or U6537 (N_6537,N_5049,N_5397);
nor U6538 (N_6538,N_5614,N_5360);
and U6539 (N_6539,N_5322,N_5055);
or U6540 (N_6540,N_5059,N_5958);
or U6541 (N_6541,N_5592,N_5760);
and U6542 (N_6542,N_5229,N_5090);
nor U6543 (N_6543,N_5173,N_5869);
and U6544 (N_6544,N_5584,N_5160);
or U6545 (N_6545,N_5828,N_5309);
and U6546 (N_6546,N_5506,N_5688);
and U6547 (N_6547,N_5122,N_5410);
and U6548 (N_6548,N_5643,N_5590);
or U6549 (N_6549,N_5222,N_5977);
or U6550 (N_6550,N_5528,N_5486);
and U6551 (N_6551,N_5175,N_5583);
and U6552 (N_6552,N_5838,N_5323);
nand U6553 (N_6553,N_5399,N_5418);
nand U6554 (N_6554,N_5501,N_5126);
and U6555 (N_6555,N_5333,N_5903);
nand U6556 (N_6556,N_5110,N_5319);
nand U6557 (N_6557,N_5106,N_5953);
nand U6558 (N_6558,N_5715,N_5354);
nand U6559 (N_6559,N_5448,N_5248);
or U6560 (N_6560,N_5146,N_5727);
nand U6561 (N_6561,N_5651,N_5202);
and U6562 (N_6562,N_5076,N_5311);
and U6563 (N_6563,N_5346,N_5463);
or U6564 (N_6564,N_5145,N_5795);
nand U6565 (N_6565,N_5040,N_5160);
nor U6566 (N_6566,N_5474,N_5508);
and U6567 (N_6567,N_5600,N_5581);
or U6568 (N_6568,N_5235,N_5979);
or U6569 (N_6569,N_5609,N_5610);
and U6570 (N_6570,N_5216,N_5682);
nor U6571 (N_6571,N_5827,N_5103);
nand U6572 (N_6572,N_5426,N_5658);
or U6573 (N_6573,N_5988,N_5422);
and U6574 (N_6574,N_5080,N_5652);
or U6575 (N_6575,N_5156,N_5381);
nor U6576 (N_6576,N_5998,N_5660);
and U6577 (N_6577,N_5339,N_5107);
nand U6578 (N_6578,N_5709,N_5081);
or U6579 (N_6579,N_5882,N_5059);
xnor U6580 (N_6580,N_5893,N_5890);
or U6581 (N_6581,N_5214,N_5253);
nand U6582 (N_6582,N_5933,N_5086);
or U6583 (N_6583,N_5634,N_5403);
nand U6584 (N_6584,N_5178,N_5137);
and U6585 (N_6585,N_5481,N_5893);
or U6586 (N_6586,N_5644,N_5649);
and U6587 (N_6587,N_5100,N_5071);
and U6588 (N_6588,N_5738,N_5067);
or U6589 (N_6589,N_5883,N_5614);
nand U6590 (N_6590,N_5943,N_5539);
and U6591 (N_6591,N_5327,N_5915);
nor U6592 (N_6592,N_5064,N_5732);
and U6593 (N_6593,N_5843,N_5938);
and U6594 (N_6594,N_5938,N_5172);
nand U6595 (N_6595,N_5825,N_5995);
nor U6596 (N_6596,N_5427,N_5858);
and U6597 (N_6597,N_5218,N_5297);
nand U6598 (N_6598,N_5282,N_5668);
nor U6599 (N_6599,N_5229,N_5325);
or U6600 (N_6600,N_5411,N_5334);
or U6601 (N_6601,N_5654,N_5408);
nand U6602 (N_6602,N_5691,N_5034);
and U6603 (N_6603,N_5338,N_5131);
and U6604 (N_6604,N_5229,N_5523);
nand U6605 (N_6605,N_5629,N_5828);
nor U6606 (N_6606,N_5501,N_5076);
and U6607 (N_6607,N_5425,N_5633);
and U6608 (N_6608,N_5727,N_5628);
or U6609 (N_6609,N_5203,N_5860);
or U6610 (N_6610,N_5124,N_5174);
nand U6611 (N_6611,N_5723,N_5462);
and U6612 (N_6612,N_5139,N_5535);
nor U6613 (N_6613,N_5770,N_5008);
or U6614 (N_6614,N_5857,N_5844);
and U6615 (N_6615,N_5000,N_5646);
nand U6616 (N_6616,N_5449,N_5312);
and U6617 (N_6617,N_5591,N_5320);
nor U6618 (N_6618,N_5338,N_5104);
and U6619 (N_6619,N_5252,N_5492);
or U6620 (N_6620,N_5367,N_5278);
xnor U6621 (N_6621,N_5572,N_5880);
and U6622 (N_6622,N_5394,N_5940);
or U6623 (N_6623,N_5638,N_5782);
and U6624 (N_6624,N_5924,N_5486);
nand U6625 (N_6625,N_5640,N_5693);
xnor U6626 (N_6626,N_5773,N_5450);
or U6627 (N_6627,N_5954,N_5089);
and U6628 (N_6628,N_5148,N_5063);
xnor U6629 (N_6629,N_5058,N_5581);
nand U6630 (N_6630,N_5034,N_5841);
or U6631 (N_6631,N_5462,N_5166);
nor U6632 (N_6632,N_5009,N_5933);
or U6633 (N_6633,N_5844,N_5758);
nand U6634 (N_6634,N_5432,N_5858);
and U6635 (N_6635,N_5255,N_5067);
or U6636 (N_6636,N_5511,N_5050);
and U6637 (N_6637,N_5084,N_5417);
and U6638 (N_6638,N_5125,N_5807);
nand U6639 (N_6639,N_5189,N_5748);
and U6640 (N_6640,N_5580,N_5233);
nand U6641 (N_6641,N_5631,N_5387);
nor U6642 (N_6642,N_5773,N_5223);
nor U6643 (N_6643,N_5077,N_5671);
or U6644 (N_6644,N_5905,N_5782);
nand U6645 (N_6645,N_5746,N_5114);
nand U6646 (N_6646,N_5037,N_5612);
or U6647 (N_6647,N_5435,N_5142);
nand U6648 (N_6648,N_5804,N_5111);
and U6649 (N_6649,N_5002,N_5838);
nor U6650 (N_6650,N_5634,N_5877);
or U6651 (N_6651,N_5566,N_5423);
or U6652 (N_6652,N_5259,N_5685);
and U6653 (N_6653,N_5728,N_5249);
or U6654 (N_6654,N_5784,N_5588);
nor U6655 (N_6655,N_5431,N_5795);
and U6656 (N_6656,N_5217,N_5179);
and U6657 (N_6657,N_5918,N_5769);
nand U6658 (N_6658,N_5203,N_5226);
nand U6659 (N_6659,N_5969,N_5699);
and U6660 (N_6660,N_5803,N_5156);
nand U6661 (N_6661,N_5449,N_5646);
nand U6662 (N_6662,N_5331,N_5393);
or U6663 (N_6663,N_5317,N_5952);
and U6664 (N_6664,N_5539,N_5198);
or U6665 (N_6665,N_5475,N_5086);
and U6666 (N_6666,N_5905,N_5488);
and U6667 (N_6667,N_5254,N_5437);
or U6668 (N_6668,N_5532,N_5674);
nand U6669 (N_6669,N_5229,N_5789);
or U6670 (N_6670,N_5686,N_5248);
nand U6671 (N_6671,N_5813,N_5911);
nor U6672 (N_6672,N_5203,N_5173);
nand U6673 (N_6673,N_5013,N_5884);
nor U6674 (N_6674,N_5691,N_5172);
and U6675 (N_6675,N_5980,N_5289);
and U6676 (N_6676,N_5321,N_5657);
nand U6677 (N_6677,N_5248,N_5349);
nor U6678 (N_6678,N_5591,N_5327);
nand U6679 (N_6679,N_5319,N_5492);
or U6680 (N_6680,N_5408,N_5655);
nor U6681 (N_6681,N_5788,N_5170);
nand U6682 (N_6682,N_5087,N_5156);
and U6683 (N_6683,N_5811,N_5399);
and U6684 (N_6684,N_5314,N_5235);
nor U6685 (N_6685,N_5182,N_5826);
nand U6686 (N_6686,N_5673,N_5092);
nor U6687 (N_6687,N_5989,N_5163);
and U6688 (N_6688,N_5290,N_5157);
and U6689 (N_6689,N_5522,N_5893);
and U6690 (N_6690,N_5156,N_5000);
nor U6691 (N_6691,N_5502,N_5036);
or U6692 (N_6692,N_5089,N_5591);
nor U6693 (N_6693,N_5798,N_5598);
nor U6694 (N_6694,N_5901,N_5936);
nand U6695 (N_6695,N_5583,N_5750);
xor U6696 (N_6696,N_5902,N_5474);
nor U6697 (N_6697,N_5573,N_5164);
nand U6698 (N_6698,N_5962,N_5797);
and U6699 (N_6699,N_5033,N_5784);
or U6700 (N_6700,N_5381,N_5264);
nand U6701 (N_6701,N_5625,N_5476);
or U6702 (N_6702,N_5132,N_5367);
nand U6703 (N_6703,N_5418,N_5657);
or U6704 (N_6704,N_5002,N_5147);
and U6705 (N_6705,N_5195,N_5262);
or U6706 (N_6706,N_5685,N_5490);
or U6707 (N_6707,N_5915,N_5364);
nor U6708 (N_6708,N_5628,N_5992);
xnor U6709 (N_6709,N_5231,N_5424);
nor U6710 (N_6710,N_5276,N_5212);
and U6711 (N_6711,N_5300,N_5039);
and U6712 (N_6712,N_5497,N_5037);
and U6713 (N_6713,N_5617,N_5875);
and U6714 (N_6714,N_5749,N_5103);
and U6715 (N_6715,N_5419,N_5717);
nor U6716 (N_6716,N_5364,N_5110);
or U6717 (N_6717,N_5753,N_5316);
nand U6718 (N_6718,N_5292,N_5878);
or U6719 (N_6719,N_5993,N_5831);
nor U6720 (N_6720,N_5608,N_5890);
nor U6721 (N_6721,N_5888,N_5827);
and U6722 (N_6722,N_5222,N_5990);
nor U6723 (N_6723,N_5220,N_5251);
nand U6724 (N_6724,N_5884,N_5253);
and U6725 (N_6725,N_5373,N_5051);
nor U6726 (N_6726,N_5934,N_5642);
nor U6727 (N_6727,N_5329,N_5123);
nand U6728 (N_6728,N_5523,N_5448);
nand U6729 (N_6729,N_5620,N_5248);
or U6730 (N_6730,N_5101,N_5405);
or U6731 (N_6731,N_5571,N_5217);
nand U6732 (N_6732,N_5654,N_5705);
or U6733 (N_6733,N_5889,N_5181);
nand U6734 (N_6734,N_5231,N_5007);
nand U6735 (N_6735,N_5584,N_5995);
xor U6736 (N_6736,N_5803,N_5873);
or U6737 (N_6737,N_5237,N_5406);
and U6738 (N_6738,N_5404,N_5549);
nor U6739 (N_6739,N_5424,N_5999);
nor U6740 (N_6740,N_5648,N_5663);
nor U6741 (N_6741,N_5043,N_5733);
nor U6742 (N_6742,N_5490,N_5686);
nor U6743 (N_6743,N_5847,N_5878);
nand U6744 (N_6744,N_5687,N_5519);
nor U6745 (N_6745,N_5760,N_5810);
xnor U6746 (N_6746,N_5291,N_5031);
and U6747 (N_6747,N_5942,N_5049);
and U6748 (N_6748,N_5740,N_5589);
and U6749 (N_6749,N_5185,N_5288);
or U6750 (N_6750,N_5356,N_5304);
xnor U6751 (N_6751,N_5019,N_5229);
nand U6752 (N_6752,N_5189,N_5461);
nor U6753 (N_6753,N_5363,N_5154);
and U6754 (N_6754,N_5560,N_5581);
or U6755 (N_6755,N_5193,N_5319);
nand U6756 (N_6756,N_5452,N_5182);
nand U6757 (N_6757,N_5807,N_5143);
nand U6758 (N_6758,N_5745,N_5783);
nand U6759 (N_6759,N_5439,N_5401);
and U6760 (N_6760,N_5241,N_5551);
nand U6761 (N_6761,N_5936,N_5036);
or U6762 (N_6762,N_5681,N_5127);
nand U6763 (N_6763,N_5461,N_5935);
and U6764 (N_6764,N_5850,N_5954);
or U6765 (N_6765,N_5828,N_5647);
or U6766 (N_6766,N_5921,N_5607);
nand U6767 (N_6767,N_5634,N_5693);
or U6768 (N_6768,N_5478,N_5277);
or U6769 (N_6769,N_5661,N_5549);
nor U6770 (N_6770,N_5690,N_5674);
nand U6771 (N_6771,N_5718,N_5945);
nor U6772 (N_6772,N_5375,N_5374);
and U6773 (N_6773,N_5446,N_5177);
nand U6774 (N_6774,N_5997,N_5830);
or U6775 (N_6775,N_5607,N_5418);
nor U6776 (N_6776,N_5158,N_5903);
and U6777 (N_6777,N_5785,N_5864);
nand U6778 (N_6778,N_5910,N_5334);
and U6779 (N_6779,N_5926,N_5463);
and U6780 (N_6780,N_5471,N_5429);
and U6781 (N_6781,N_5778,N_5980);
nor U6782 (N_6782,N_5626,N_5756);
or U6783 (N_6783,N_5123,N_5241);
or U6784 (N_6784,N_5393,N_5555);
nor U6785 (N_6785,N_5459,N_5909);
nor U6786 (N_6786,N_5163,N_5232);
nand U6787 (N_6787,N_5314,N_5898);
nand U6788 (N_6788,N_5921,N_5487);
nor U6789 (N_6789,N_5028,N_5046);
nand U6790 (N_6790,N_5335,N_5894);
nand U6791 (N_6791,N_5200,N_5262);
and U6792 (N_6792,N_5381,N_5793);
and U6793 (N_6793,N_5867,N_5920);
or U6794 (N_6794,N_5981,N_5092);
nand U6795 (N_6795,N_5907,N_5171);
and U6796 (N_6796,N_5658,N_5669);
nor U6797 (N_6797,N_5162,N_5072);
xnor U6798 (N_6798,N_5216,N_5324);
nand U6799 (N_6799,N_5051,N_5165);
nor U6800 (N_6800,N_5914,N_5187);
or U6801 (N_6801,N_5763,N_5714);
and U6802 (N_6802,N_5810,N_5605);
nand U6803 (N_6803,N_5753,N_5839);
nor U6804 (N_6804,N_5957,N_5238);
nor U6805 (N_6805,N_5346,N_5840);
and U6806 (N_6806,N_5555,N_5103);
nor U6807 (N_6807,N_5460,N_5853);
nor U6808 (N_6808,N_5067,N_5001);
nor U6809 (N_6809,N_5406,N_5554);
nand U6810 (N_6810,N_5073,N_5250);
nand U6811 (N_6811,N_5152,N_5928);
and U6812 (N_6812,N_5884,N_5417);
and U6813 (N_6813,N_5645,N_5679);
or U6814 (N_6814,N_5345,N_5065);
nor U6815 (N_6815,N_5082,N_5319);
nor U6816 (N_6816,N_5053,N_5420);
or U6817 (N_6817,N_5706,N_5860);
nand U6818 (N_6818,N_5983,N_5247);
nor U6819 (N_6819,N_5694,N_5482);
or U6820 (N_6820,N_5002,N_5690);
nand U6821 (N_6821,N_5343,N_5736);
nand U6822 (N_6822,N_5516,N_5653);
and U6823 (N_6823,N_5577,N_5389);
nand U6824 (N_6824,N_5007,N_5779);
nand U6825 (N_6825,N_5995,N_5274);
nand U6826 (N_6826,N_5289,N_5172);
nor U6827 (N_6827,N_5660,N_5962);
and U6828 (N_6828,N_5195,N_5899);
nand U6829 (N_6829,N_5453,N_5746);
nand U6830 (N_6830,N_5115,N_5923);
or U6831 (N_6831,N_5788,N_5873);
nand U6832 (N_6832,N_5618,N_5275);
nand U6833 (N_6833,N_5111,N_5017);
or U6834 (N_6834,N_5347,N_5941);
or U6835 (N_6835,N_5640,N_5584);
or U6836 (N_6836,N_5057,N_5509);
or U6837 (N_6837,N_5718,N_5244);
and U6838 (N_6838,N_5608,N_5914);
and U6839 (N_6839,N_5491,N_5745);
or U6840 (N_6840,N_5570,N_5318);
nand U6841 (N_6841,N_5908,N_5905);
nor U6842 (N_6842,N_5833,N_5695);
or U6843 (N_6843,N_5703,N_5515);
or U6844 (N_6844,N_5943,N_5933);
or U6845 (N_6845,N_5354,N_5890);
or U6846 (N_6846,N_5121,N_5856);
and U6847 (N_6847,N_5337,N_5659);
or U6848 (N_6848,N_5208,N_5418);
nand U6849 (N_6849,N_5054,N_5283);
and U6850 (N_6850,N_5420,N_5553);
nand U6851 (N_6851,N_5784,N_5404);
xor U6852 (N_6852,N_5308,N_5666);
nor U6853 (N_6853,N_5813,N_5832);
and U6854 (N_6854,N_5816,N_5439);
nand U6855 (N_6855,N_5843,N_5690);
nor U6856 (N_6856,N_5448,N_5814);
nor U6857 (N_6857,N_5294,N_5823);
and U6858 (N_6858,N_5586,N_5182);
nor U6859 (N_6859,N_5288,N_5652);
nor U6860 (N_6860,N_5358,N_5050);
nand U6861 (N_6861,N_5311,N_5425);
or U6862 (N_6862,N_5694,N_5758);
or U6863 (N_6863,N_5189,N_5438);
and U6864 (N_6864,N_5426,N_5101);
nor U6865 (N_6865,N_5808,N_5031);
nand U6866 (N_6866,N_5873,N_5961);
nand U6867 (N_6867,N_5134,N_5350);
and U6868 (N_6868,N_5018,N_5775);
nor U6869 (N_6869,N_5376,N_5984);
nand U6870 (N_6870,N_5889,N_5615);
or U6871 (N_6871,N_5868,N_5436);
nor U6872 (N_6872,N_5884,N_5042);
nor U6873 (N_6873,N_5835,N_5325);
nand U6874 (N_6874,N_5420,N_5684);
and U6875 (N_6875,N_5119,N_5004);
nor U6876 (N_6876,N_5357,N_5625);
nor U6877 (N_6877,N_5195,N_5551);
or U6878 (N_6878,N_5498,N_5493);
and U6879 (N_6879,N_5469,N_5360);
and U6880 (N_6880,N_5400,N_5662);
nor U6881 (N_6881,N_5397,N_5561);
nand U6882 (N_6882,N_5167,N_5008);
nor U6883 (N_6883,N_5457,N_5294);
nand U6884 (N_6884,N_5999,N_5130);
and U6885 (N_6885,N_5470,N_5715);
nand U6886 (N_6886,N_5339,N_5353);
and U6887 (N_6887,N_5029,N_5785);
or U6888 (N_6888,N_5922,N_5912);
or U6889 (N_6889,N_5551,N_5181);
and U6890 (N_6890,N_5911,N_5499);
or U6891 (N_6891,N_5114,N_5819);
nor U6892 (N_6892,N_5243,N_5151);
or U6893 (N_6893,N_5367,N_5075);
or U6894 (N_6894,N_5785,N_5465);
nand U6895 (N_6895,N_5303,N_5573);
nand U6896 (N_6896,N_5544,N_5637);
nor U6897 (N_6897,N_5555,N_5013);
or U6898 (N_6898,N_5688,N_5615);
or U6899 (N_6899,N_5923,N_5386);
nor U6900 (N_6900,N_5208,N_5455);
and U6901 (N_6901,N_5055,N_5625);
and U6902 (N_6902,N_5620,N_5211);
or U6903 (N_6903,N_5193,N_5850);
nor U6904 (N_6904,N_5622,N_5036);
nand U6905 (N_6905,N_5674,N_5702);
nor U6906 (N_6906,N_5012,N_5684);
nor U6907 (N_6907,N_5295,N_5650);
nor U6908 (N_6908,N_5625,N_5761);
nor U6909 (N_6909,N_5235,N_5552);
nand U6910 (N_6910,N_5858,N_5362);
nand U6911 (N_6911,N_5098,N_5065);
nand U6912 (N_6912,N_5020,N_5189);
and U6913 (N_6913,N_5116,N_5854);
nand U6914 (N_6914,N_5777,N_5552);
nand U6915 (N_6915,N_5711,N_5771);
xnor U6916 (N_6916,N_5931,N_5461);
nand U6917 (N_6917,N_5661,N_5082);
nand U6918 (N_6918,N_5692,N_5755);
nand U6919 (N_6919,N_5007,N_5516);
and U6920 (N_6920,N_5032,N_5170);
and U6921 (N_6921,N_5412,N_5526);
or U6922 (N_6922,N_5622,N_5054);
nor U6923 (N_6923,N_5005,N_5573);
nor U6924 (N_6924,N_5582,N_5923);
or U6925 (N_6925,N_5756,N_5366);
nor U6926 (N_6926,N_5078,N_5226);
or U6927 (N_6927,N_5171,N_5375);
and U6928 (N_6928,N_5812,N_5340);
nor U6929 (N_6929,N_5169,N_5299);
and U6930 (N_6930,N_5318,N_5252);
or U6931 (N_6931,N_5726,N_5636);
nor U6932 (N_6932,N_5298,N_5736);
nor U6933 (N_6933,N_5076,N_5778);
nand U6934 (N_6934,N_5344,N_5424);
or U6935 (N_6935,N_5512,N_5024);
nor U6936 (N_6936,N_5503,N_5409);
nor U6937 (N_6937,N_5547,N_5619);
and U6938 (N_6938,N_5536,N_5132);
nand U6939 (N_6939,N_5062,N_5043);
nor U6940 (N_6940,N_5962,N_5674);
nand U6941 (N_6941,N_5543,N_5716);
nand U6942 (N_6942,N_5389,N_5905);
nand U6943 (N_6943,N_5442,N_5385);
and U6944 (N_6944,N_5909,N_5686);
or U6945 (N_6945,N_5440,N_5647);
nand U6946 (N_6946,N_5397,N_5648);
or U6947 (N_6947,N_5028,N_5012);
nor U6948 (N_6948,N_5858,N_5158);
and U6949 (N_6949,N_5993,N_5411);
and U6950 (N_6950,N_5821,N_5540);
nand U6951 (N_6951,N_5500,N_5231);
nand U6952 (N_6952,N_5342,N_5997);
nor U6953 (N_6953,N_5014,N_5260);
nand U6954 (N_6954,N_5401,N_5537);
or U6955 (N_6955,N_5605,N_5898);
nand U6956 (N_6956,N_5324,N_5878);
or U6957 (N_6957,N_5420,N_5355);
nor U6958 (N_6958,N_5062,N_5522);
nand U6959 (N_6959,N_5565,N_5293);
and U6960 (N_6960,N_5500,N_5358);
nand U6961 (N_6961,N_5094,N_5530);
and U6962 (N_6962,N_5189,N_5253);
and U6963 (N_6963,N_5570,N_5167);
or U6964 (N_6964,N_5006,N_5120);
nor U6965 (N_6965,N_5187,N_5047);
or U6966 (N_6966,N_5089,N_5114);
or U6967 (N_6967,N_5535,N_5685);
nor U6968 (N_6968,N_5741,N_5029);
nor U6969 (N_6969,N_5856,N_5781);
nor U6970 (N_6970,N_5124,N_5761);
nand U6971 (N_6971,N_5770,N_5514);
nand U6972 (N_6972,N_5299,N_5888);
xor U6973 (N_6973,N_5476,N_5194);
and U6974 (N_6974,N_5621,N_5983);
nand U6975 (N_6975,N_5131,N_5119);
or U6976 (N_6976,N_5907,N_5683);
and U6977 (N_6977,N_5137,N_5628);
or U6978 (N_6978,N_5445,N_5466);
or U6979 (N_6979,N_5597,N_5755);
and U6980 (N_6980,N_5375,N_5240);
or U6981 (N_6981,N_5187,N_5212);
nand U6982 (N_6982,N_5630,N_5968);
nor U6983 (N_6983,N_5323,N_5412);
nor U6984 (N_6984,N_5588,N_5827);
nor U6985 (N_6985,N_5293,N_5377);
xnor U6986 (N_6986,N_5303,N_5662);
or U6987 (N_6987,N_5979,N_5113);
and U6988 (N_6988,N_5958,N_5273);
and U6989 (N_6989,N_5076,N_5352);
nand U6990 (N_6990,N_5592,N_5940);
nor U6991 (N_6991,N_5261,N_5705);
or U6992 (N_6992,N_5494,N_5088);
nor U6993 (N_6993,N_5741,N_5517);
and U6994 (N_6994,N_5262,N_5088);
and U6995 (N_6995,N_5608,N_5749);
nor U6996 (N_6996,N_5619,N_5887);
nor U6997 (N_6997,N_5383,N_5090);
nor U6998 (N_6998,N_5223,N_5346);
or U6999 (N_6999,N_5039,N_5730);
nor U7000 (N_7000,N_6407,N_6724);
or U7001 (N_7001,N_6196,N_6757);
and U7002 (N_7002,N_6140,N_6643);
nand U7003 (N_7003,N_6533,N_6108);
or U7004 (N_7004,N_6134,N_6043);
nor U7005 (N_7005,N_6094,N_6373);
and U7006 (N_7006,N_6613,N_6631);
and U7007 (N_7007,N_6932,N_6656);
nand U7008 (N_7008,N_6055,N_6572);
nand U7009 (N_7009,N_6560,N_6679);
or U7010 (N_7010,N_6078,N_6951);
and U7011 (N_7011,N_6761,N_6093);
and U7012 (N_7012,N_6375,N_6429);
or U7013 (N_7013,N_6061,N_6592);
nand U7014 (N_7014,N_6880,N_6746);
nor U7015 (N_7015,N_6374,N_6386);
and U7016 (N_7016,N_6050,N_6004);
and U7017 (N_7017,N_6694,N_6851);
and U7018 (N_7018,N_6818,N_6769);
nor U7019 (N_7019,N_6170,N_6228);
and U7020 (N_7020,N_6481,N_6739);
and U7021 (N_7021,N_6683,N_6822);
and U7022 (N_7022,N_6537,N_6837);
or U7023 (N_7023,N_6030,N_6825);
nand U7024 (N_7024,N_6100,N_6911);
nand U7025 (N_7025,N_6603,N_6401);
and U7026 (N_7026,N_6436,N_6570);
and U7027 (N_7027,N_6203,N_6827);
and U7028 (N_7028,N_6852,N_6379);
and U7029 (N_7029,N_6113,N_6075);
nand U7030 (N_7030,N_6678,N_6080);
nand U7031 (N_7031,N_6142,N_6706);
or U7032 (N_7032,N_6342,N_6815);
and U7033 (N_7033,N_6072,N_6276);
nor U7034 (N_7034,N_6277,N_6018);
or U7035 (N_7035,N_6202,N_6855);
or U7036 (N_7036,N_6102,N_6836);
nor U7037 (N_7037,N_6531,N_6669);
nand U7038 (N_7038,N_6804,N_6843);
nor U7039 (N_7039,N_6971,N_6892);
and U7040 (N_7040,N_6728,N_6652);
nand U7041 (N_7041,N_6771,N_6514);
and U7042 (N_7042,N_6947,N_6714);
or U7043 (N_7043,N_6585,N_6478);
nand U7044 (N_7044,N_6943,N_6922);
nor U7045 (N_7045,N_6405,N_6027);
and U7046 (N_7046,N_6748,N_6279);
nand U7047 (N_7047,N_6285,N_6150);
nor U7048 (N_7048,N_6176,N_6680);
nor U7049 (N_7049,N_6430,N_6488);
and U7050 (N_7050,N_6336,N_6053);
nand U7051 (N_7051,N_6487,N_6909);
nor U7052 (N_7052,N_6853,N_6366);
or U7053 (N_7053,N_6816,N_6671);
nand U7054 (N_7054,N_6251,N_6567);
nand U7055 (N_7055,N_6907,N_6049);
nor U7056 (N_7056,N_6525,N_6508);
or U7057 (N_7057,N_6916,N_6608);
nand U7058 (N_7058,N_6109,N_6565);
nor U7059 (N_7059,N_6820,N_6453);
nand U7060 (N_7060,N_6958,N_6335);
nand U7061 (N_7061,N_6247,N_6883);
and U7062 (N_7062,N_6520,N_6280);
nor U7063 (N_7063,N_6225,N_6237);
and U7064 (N_7064,N_6329,N_6629);
nand U7065 (N_7065,N_6535,N_6370);
nand U7066 (N_7066,N_6920,N_6242);
or U7067 (N_7067,N_6675,N_6929);
nor U7068 (N_7068,N_6458,N_6547);
nor U7069 (N_7069,N_6115,N_6505);
xor U7070 (N_7070,N_6474,N_6167);
nand U7071 (N_7071,N_6814,N_6086);
and U7072 (N_7072,N_6116,N_6574);
or U7073 (N_7073,N_6779,N_6701);
and U7074 (N_7074,N_6924,N_6578);
and U7075 (N_7075,N_6212,N_6026);
and U7076 (N_7076,N_6665,N_6979);
and U7077 (N_7077,N_6128,N_6464);
nand U7078 (N_7078,N_6034,N_6637);
nor U7079 (N_7079,N_6135,N_6318);
nor U7080 (N_7080,N_6653,N_6685);
or U7081 (N_7081,N_6391,N_6890);
nor U7082 (N_7082,N_6513,N_6785);
nor U7083 (N_7083,N_6503,N_6839);
nand U7084 (N_7084,N_6058,N_6173);
nor U7085 (N_7085,N_6500,N_6138);
or U7086 (N_7086,N_6421,N_6648);
and U7087 (N_7087,N_6449,N_6586);
nand U7088 (N_7088,N_6324,N_6232);
and U7089 (N_7089,N_6522,N_6862);
xnor U7090 (N_7090,N_6927,N_6642);
nand U7091 (N_7091,N_6337,N_6729);
nor U7092 (N_7092,N_6137,N_6017);
nand U7093 (N_7093,N_6938,N_6333);
and U7094 (N_7094,N_6295,N_6045);
xor U7095 (N_7095,N_6633,N_6409);
or U7096 (N_7096,N_6306,N_6301);
xnor U7097 (N_7097,N_6768,N_6549);
nand U7098 (N_7098,N_6332,N_6492);
or U7099 (N_7099,N_6227,N_6986);
and U7100 (N_7100,N_6817,N_6496);
nor U7101 (N_7101,N_6250,N_6670);
nor U7102 (N_7102,N_6551,N_6649);
nor U7103 (N_7103,N_6796,N_6201);
or U7104 (N_7104,N_6598,N_6107);
or U7105 (N_7105,N_6721,N_6161);
nor U7106 (N_7106,N_6681,N_6912);
nor U7107 (N_7107,N_6023,N_6730);
and U7108 (N_7108,N_6845,N_6975);
or U7109 (N_7109,N_6299,N_6666);
and U7110 (N_7110,N_6172,N_6493);
nor U7111 (N_7111,N_6068,N_6622);
or U7112 (N_7112,N_6392,N_6339);
nand U7113 (N_7113,N_6261,N_6527);
nor U7114 (N_7114,N_6347,N_6861);
and U7115 (N_7115,N_6805,N_6103);
or U7116 (N_7116,N_6127,N_6431);
nor U7117 (N_7117,N_6051,N_6315);
and U7118 (N_7118,N_6088,N_6165);
or U7119 (N_7119,N_6850,N_6899);
xor U7120 (N_7120,N_6001,N_6254);
nor U7121 (N_7121,N_6011,N_6184);
or U7122 (N_7122,N_6399,N_6171);
or U7123 (N_7123,N_6544,N_6282);
nand U7124 (N_7124,N_6875,N_6566);
nand U7125 (N_7125,N_6069,N_6793);
or U7126 (N_7126,N_6052,N_6390);
xnor U7127 (N_7127,N_6812,N_6902);
nand U7128 (N_7128,N_6777,N_6654);
nor U7129 (N_7129,N_6650,N_6949);
nand U7130 (N_7130,N_6129,N_6056);
nand U7131 (N_7131,N_6498,N_6266);
or U7132 (N_7132,N_6763,N_6998);
nand U7133 (N_7133,N_6553,N_6331);
or U7134 (N_7134,N_6040,N_6149);
nor U7135 (N_7135,N_6417,N_6047);
nand U7136 (N_7136,N_6614,N_6195);
or U7137 (N_7137,N_6600,N_6864);
and U7138 (N_7138,N_6780,N_6987);
and U7139 (N_7139,N_6575,N_6356);
and U7140 (N_7140,N_6213,N_6569);
and U7141 (N_7141,N_6036,N_6945);
and U7142 (N_7142,N_6542,N_6214);
or U7143 (N_7143,N_6857,N_6286);
nor U7144 (N_7144,N_6993,N_6450);
or U7145 (N_7145,N_6697,N_6305);
nand U7146 (N_7146,N_6709,N_6676);
nor U7147 (N_7147,N_6424,N_6084);
nor U7148 (N_7148,N_6976,N_6956);
nor U7149 (N_7149,N_6605,N_6192);
and U7150 (N_7150,N_6209,N_6766);
or U7151 (N_7151,N_6713,N_6554);
and U7152 (N_7152,N_6787,N_6988);
nor U7153 (N_7153,N_6841,N_6538);
nand U7154 (N_7154,N_6042,N_6781);
or U7155 (N_7155,N_6141,N_6151);
nor U7156 (N_7156,N_6475,N_6744);
nor U7157 (N_7157,N_6489,N_6636);
nor U7158 (N_7158,N_6658,N_6131);
or U7159 (N_7159,N_6733,N_6340);
nand U7160 (N_7160,N_6821,N_6588);
or U7161 (N_7161,N_6263,N_6868);
nor U7162 (N_7162,N_6863,N_6208);
nor U7163 (N_7163,N_6895,N_6381);
xnor U7164 (N_7164,N_6046,N_6219);
nor U7165 (N_7165,N_6917,N_6166);
or U7166 (N_7166,N_6882,N_6459);
and U7167 (N_7167,N_6104,N_6368);
and U7168 (N_7168,N_6910,N_6517);
and U7169 (N_7169,N_6624,N_6668);
or U7170 (N_7170,N_6071,N_6180);
nand U7171 (N_7171,N_6243,N_6185);
nand U7172 (N_7172,N_6904,N_6826);
or U7173 (N_7173,N_6828,N_6903);
and U7174 (N_7174,N_6400,N_6014);
or U7175 (N_7175,N_6162,N_6074);
or U7176 (N_7176,N_6749,N_6918);
or U7177 (N_7177,N_6359,N_6573);
and U7178 (N_7178,N_6581,N_6627);
and U7179 (N_7179,N_6970,N_6874);
nand U7180 (N_7180,N_6363,N_6204);
and U7181 (N_7181,N_6118,N_6959);
and U7182 (N_7182,N_6846,N_6462);
or U7183 (N_7183,N_6523,N_6978);
nand U7184 (N_7184,N_6740,N_6200);
nor U7185 (N_7185,N_6491,N_6274);
xor U7186 (N_7186,N_6898,N_6327);
nand U7187 (N_7187,N_6693,N_6638);
nand U7188 (N_7188,N_6483,N_6007);
or U7189 (N_7189,N_6252,N_6548);
nand U7190 (N_7190,N_6651,N_6473);
nor U7191 (N_7191,N_6296,N_6177);
and U7192 (N_7192,N_6799,N_6041);
nor U7193 (N_7193,N_6169,N_6532);
nand U7194 (N_7194,N_6298,N_6009);
or U7195 (N_7195,N_6419,N_6928);
nor U7196 (N_7196,N_6025,N_6644);
or U7197 (N_7197,N_6054,N_6541);
or U7198 (N_7198,N_6447,N_6550);
nand U7199 (N_7199,N_6906,N_6452);
and U7200 (N_7200,N_6418,N_6869);
nand U7201 (N_7201,N_6854,N_6188);
and U7202 (N_7202,N_6073,N_6490);
or U7203 (N_7203,N_6438,N_6380);
and U7204 (N_7204,N_6915,N_6512);
and U7205 (N_7205,N_6420,N_6844);
and U7206 (N_7206,N_6105,N_6428);
nand U7207 (N_7207,N_6992,N_6394);
nor U7208 (N_7208,N_6408,N_6509);
and U7209 (N_7209,N_6832,N_6194);
and U7210 (N_7210,N_6322,N_6396);
nand U7211 (N_7211,N_6765,N_6376);
and U7212 (N_7212,N_6702,N_6179);
nand U7213 (N_7213,N_6530,N_6230);
nor U7214 (N_7214,N_6302,N_6155);
or U7215 (N_7215,N_6309,N_6722);
nand U7216 (N_7216,N_6265,N_6884);
nand U7217 (N_7217,N_6686,N_6361);
nand U7218 (N_7218,N_6737,N_6595);
nand U7219 (N_7219,N_6321,N_6389);
and U7220 (N_7220,N_6754,N_6536);
nand U7221 (N_7221,N_6433,N_6121);
nand U7222 (N_7222,N_6434,N_6372);
or U7223 (N_7223,N_6346,N_6645);
nor U7224 (N_7224,N_6270,N_6931);
nor U7225 (N_7225,N_6704,N_6939);
nor U7226 (N_7226,N_6002,N_6705);
and U7227 (N_7227,N_6289,N_6344);
nand U7228 (N_7228,N_6031,N_6308);
nor U7229 (N_7229,N_6300,N_6406);
and U7230 (N_7230,N_6634,N_6222);
xnor U7231 (N_7231,N_6881,N_6039);
nor U7232 (N_7232,N_6557,N_6038);
or U7233 (N_7233,N_6096,N_6894);
nand U7234 (N_7234,N_6293,N_6936);
or U7235 (N_7235,N_6905,N_6745);
or U7236 (N_7236,N_6136,N_6620);
nor U7237 (N_7237,N_6000,N_6231);
nand U7238 (N_7238,N_6707,N_6081);
nor U7239 (N_7239,N_6153,N_6476);
nor U7240 (N_7240,N_6619,N_6290);
nor U7241 (N_7241,N_6067,N_6689);
and U7242 (N_7242,N_6995,N_6596);
nor U7243 (N_7243,N_6753,N_6930);
or U7244 (N_7244,N_6360,N_6354);
nand U7245 (N_7245,N_6019,N_6969);
and U7246 (N_7246,N_6085,N_6893);
and U7247 (N_7247,N_6616,N_6989);
nor U7248 (N_7248,N_6253,N_6819);
nand U7249 (N_7249,N_6024,N_6715);
and U7250 (N_7250,N_6568,N_6143);
nand U7251 (N_7251,N_6425,N_6618);
or U7252 (N_7252,N_6504,N_6256);
or U7253 (N_7253,N_6583,N_6580);
nor U7254 (N_7254,N_6524,N_6539);
nand U7255 (N_7255,N_6145,N_6960);
and U7256 (N_7256,N_6692,N_6404);
nor U7257 (N_7257,N_6482,N_6211);
nand U7258 (N_7258,N_6365,N_6840);
and U7259 (N_7259,N_6510,N_6241);
xor U7260 (N_7260,N_6220,N_6558);
nor U7261 (N_7261,N_6092,N_6997);
or U7262 (N_7262,N_6160,N_6888);
or U7263 (N_7263,N_6602,N_6953);
nor U7264 (N_7264,N_6091,N_6807);
nand U7265 (N_7265,N_6786,N_6860);
nand U7266 (N_7266,N_6106,N_6355);
nor U7267 (N_7267,N_6190,N_6593);
nor U7268 (N_7268,N_6798,N_6515);
and U7269 (N_7269,N_6609,N_6772);
nand U7270 (N_7270,N_6782,N_6454);
and U7271 (N_7271,N_6528,N_6168);
nand U7272 (N_7272,N_6157,N_6008);
and U7273 (N_7273,N_6700,N_6062);
nor U7274 (N_7274,N_6224,N_6472);
nand U7275 (N_7275,N_6579,N_6314);
or U7276 (N_7276,N_6788,N_6334);
nor U7277 (N_7277,N_6878,N_6688);
and U7278 (N_7278,N_6506,N_6994);
or U7279 (N_7279,N_6747,N_6199);
nor U7280 (N_7280,N_6885,N_6385);
or U7281 (N_7281,N_6887,N_6552);
or U7282 (N_7282,N_6889,N_6441);
nor U7283 (N_7283,N_6626,N_6245);
nand U7284 (N_7284,N_6639,N_6126);
or U7285 (N_7285,N_6325,N_6234);
or U7286 (N_7286,N_6082,N_6159);
or U7287 (N_7287,N_6980,N_6154);
nor U7288 (N_7288,N_6789,N_6123);
nand U7289 (N_7289,N_6499,N_6662);
and U7290 (N_7290,N_6858,N_6236);
nand U7291 (N_7291,N_6193,N_6288);
or U7292 (N_7292,N_6469,N_6756);
or U7293 (N_7293,N_6991,N_6809);
nand U7294 (N_7294,N_6210,N_6743);
xor U7295 (N_7295,N_6935,N_6221);
nor U7296 (N_7296,N_6182,N_6316);
nand U7297 (N_7297,N_6249,N_6601);
and U7298 (N_7298,N_6268,N_6621);
or U7299 (N_7299,N_6486,N_6925);
and U7300 (N_7300,N_6451,N_6711);
nand U7301 (N_7301,N_6901,N_6823);
nand U7302 (N_7302,N_6238,N_6272);
xor U7303 (N_7303,N_6087,N_6003);
nor U7304 (N_7304,N_6442,N_6708);
nand U7305 (N_7305,N_6217,N_6511);
and U7306 (N_7306,N_6577,N_6687);
nor U7307 (N_7307,N_6132,N_6526);
nor U7308 (N_7308,N_6770,N_6738);
nor U7309 (N_7309,N_6759,N_6156);
and U7310 (N_7310,N_6967,N_6076);
or U7311 (N_7311,N_6114,N_6571);
nand U7312 (N_7312,N_6383,N_6673);
nor U7313 (N_7313,N_6964,N_6873);
or U7314 (N_7314,N_6016,N_6961);
nand U7315 (N_7315,N_6628,N_6727);
or U7316 (N_7316,N_6849,N_6582);
nor U7317 (N_7317,N_6240,N_6948);
xor U7318 (N_7318,N_6507,N_6742);
or U7319 (N_7319,N_6388,N_6985);
nor U7320 (N_7320,N_6133,N_6940);
nand U7321 (N_7321,N_6158,N_6264);
nand U7322 (N_7322,N_6233,N_6833);
or U7323 (N_7323,N_6735,N_6957);
nor U7324 (N_7324,N_6886,N_6303);
nand U7325 (N_7325,N_6358,N_6556);
nand U7326 (N_7326,N_6124,N_6284);
and U7327 (N_7327,N_6750,N_6501);
and U7328 (N_7328,N_6926,N_6005);
and U7329 (N_7329,N_6612,N_6720);
nor U7330 (N_7330,N_6604,N_6647);
nand U7331 (N_7331,N_6364,N_6831);
nor U7332 (N_7332,N_6033,N_6830);
or U7333 (N_7333,N_6235,N_6856);
nor U7334 (N_7334,N_6690,N_6246);
or U7335 (N_7335,N_6802,N_6206);
or U7336 (N_7336,N_6682,N_6540);
nand U7337 (N_7337,N_6632,N_6741);
nor U7338 (N_7338,N_6187,N_6130);
nand U7339 (N_7339,N_6731,N_6012);
nand U7340 (N_7340,N_6269,N_6181);
and U7341 (N_7341,N_6345,N_6963);
or U7342 (N_7342,N_6066,N_6677);
or U7343 (N_7343,N_6393,N_6921);
and U7344 (N_7344,N_6516,N_6981);
and U7345 (N_7345,N_6990,N_6640);
or U7346 (N_7346,N_6435,N_6463);
nand U7347 (N_7347,N_6941,N_6444);
or U7348 (N_7348,N_6294,N_6371);
or U7349 (N_7349,N_6446,N_6937);
nor U7350 (N_7350,N_6271,N_6021);
nor U7351 (N_7351,N_6800,N_6946);
and U7352 (N_7352,N_6457,N_6343);
and U7353 (N_7353,N_6223,N_6350);
and U7354 (N_7354,N_6432,N_6426);
or U7355 (N_7355,N_6952,N_6411);
and U7356 (N_7356,N_6077,N_6767);
or U7357 (N_7357,N_6838,N_6468);
nand U7358 (N_7358,N_6734,N_6144);
nor U7359 (N_7359,N_6467,N_6186);
nor U7360 (N_7360,N_6518,N_6502);
and U7361 (N_7361,N_6664,N_6378);
nand U7362 (N_7362,N_6283,N_6497);
nor U7363 (N_7363,N_6257,N_6872);
and U7364 (N_7364,N_6035,N_6934);
or U7365 (N_7365,N_6764,N_6696);
nor U7366 (N_7366,N_6175,N_6439);
nand U7367 (N_7367,N_6125,N_6752);
and U7368 (N_7368,N_6348,N_6762);
or U7369 (N_7369,N_6362,N_6944);
nand U7370 (N_7370,N_6555,N_6367);
nor U7371 (N_7371,N_6663,N_6465);
or U7372 (N_7372,N_6607,N_6797);
or U7373 (N_7373,N_6037,N_6543);
nor U7374 (N_7374,N_6328,N_6312);
and U7375 (N_7375,N_6723,N_6848);
or U7376 (N_7376,N_6703,N_6529);
nor U7377 (N_7377,N_6323,N_6095);
and U7378 (N_7378,N_6415,N_6477);
and U7379 (N_7379,N_6755,N_6010);
or U7380 (N_7380,N_6972,N_6589);
nand U7381 (N_7381,N_6877,N_6174);
and U7382 (N_7382,N_6695,N_6657);
xor U7383 (N_7383,N_6495,N_6484);
or U7384 (N_7384,N_6122,N_6044);
nand U7385 (N_7385,N_6732,N_6519);
nor U7386 (N_7386,N_6984,N_6659);
or U7387 (N_7387,N_6590,N_6260);
or U7388 (N_7388,N_6774,N_6866);
nor U7389 (N_7389,N_6778,N_6120);
and U7390 (N_7390,N_6891,N_6835);
xnor U7391 (N_7391,N_6006,N_6455);
nand U7392 (N_7392,N_6377,N_6672);
or U7393 (N_7393,N_6353,N_6471);
or U7394 (N_7394,N_6859,N_6965);
or U7395 (N_7395,N_6824,N_6919);
or U7396 (N_7396,N_6413,N_6661);
nand U7397 (N_7397,N_6726,N_6291);
and U7398 (N_7398,N_6865,N_6278);
or U7399 (N_7399,N_6189,N_6258);
and U7400 (N_7400,N_6273,N_6968);
nand U7401 (N_7401,N_6561,N_6423);
nand U7402 (N_7402,N_6028,N_6775);
nor U7403 (N_7403,N_6625,N_6218);
or U7404 (N_7404,N_6834,N_6896);
nor U7405 (N_7405,N_6773,N_6229);
nor U7406 (N_7406,N_6717,N_6416);
and U7407 (N_7407,N_6576,N_6760);
and U7408 (N_7408,N_6545,N_6244);
or U7409 (N_7409,N_6563,N_6466);
nand U7410 (N_7410,N_6599,N_6148);
nor U7411 (N_7411,N_6810,N_6382);
xor U7412 (N_7412,N_6606,N_6908);
xor U7413 (N_7413,N_6089,N_6758);
or U7414 (N_7414,N_6205,N_6674);
nand U7415 (N_7415,N_6032,N_6725);
or U7416 (N_7416,N_6461,N_6262);
and U7417 (N_7417,N_6097,N_6456);
or U7418 (N_7418,N_6801,N_6973);
nor U7419 (N_7419,N_6790,N_6191);
nand U7420 (N_7420,N_6795,N_6448);
nand U7421 (N_7421,N_6617,N_6384);
or U7422 (N_7422,N_6597,N_6445);
nor U7423 (N_7423,N_6326,N_6351);
or U7424 (N_7424,N_6829,N_6317);
or U7425 (N_7425,N_6164,N_6587);
nand U7426 (N_7426,N_6983,N_6139);
nor U7427 (N_7427,N_6410,N_6808);
or U7428 (N_7428,N_6879,N_6402);
nand U7429 (N_7429,N_6776,N_6015);
nor U7430 (N_7430,N_6914,N_6784);
and U7431 (N_7431,N_6803,N_6090);
nor U7432 (N_7432,N_6111,N_6064);
and U7433 (N_7433,N_6630,N_6422);
nand U7434 (N_7434,N_6099,N_6655);
and U7435 (N_7435,N_6440,N_6320);
or U7436 (N_7436,N_6564,N_6255);
nand U7437 (N_7437,N_6546,N_6292);
nor U7438 (N_7438,N_6146,N_6736);
or U7439 (N_7439,N_6641,N_6057);
nand U7440 (N_7440,N_6806,N_6307);
or U7441 (N_7441,N_6395,N_6083);
or U7442 (N_7442,N_6594,N_6398);
nor U7443 (N_7443,N_6313,N_6020);
and U7444 (N_7444,N_6022,N_6876);
nor U7445 (N_7445,N_6267,N_6684);
or U7446 (N_7446,N_6427,N_6534);
and U7447 (N_7447,N_6867,N_6147);
or U7448 (N_7448,N_6611,N_6699);
nor U7449 (N_7449,N_6197,N_6999);
and U7450 (N_7450,N_6369,N_6215);
and U7451 (N_7451,N_6847,N_6387);
or U7452 (N_7452,N_6751,N_6101);
nand U7453 (N_7453,N_6792,N_6623);
nor U7454 (N_7454,N_6259,N_6982);
or U7455 (N_7455,N_6584,N_6610);
and U7456 (N_7456,N_6412,N_6950);
or U7457 (N_7457,N_6112,N_6485);
or U7458 (N_7458,N_6974,N_6954);
nor U7459 (N_7459,N_6691,N_6719);
nand U7460 (N_7460,N_6660,N_6479);
nor U7461 (N_7461,N_6319,N_6239);
or U7462 (N_7462,N_6330,N_6635);
and U7463 (N_7463,N_6842,N_6521);
and U7464 (N_7464,N_6933,N_6281);
nand U7465 (N_7465,N_6470,N_6207);
or U7466 (N_7466,N_6966,N_6338);
nand U7467 (N_7467,N_6065,N_6646);
or U7468 (N_7468,N_6437,N_6152);
nor U7469 (N_7469,N_6226,N_6048);
or U7470 (N_7470,N_6460,N_6480);
and U7471 (N_7471,N_6897,N_6059);
nor U7472 (N_7472,N_6811,N_6063);
nor U7473 (N_7473,N_6117,N_6079);
and U7474 (N_7474,N_6216,N_6716);
nor U7475 (N_7475,N_6349,N_6357);
nand U7476 (N_7476,N_6060,N_6923);
and U7477 (N_7477,N_6562,N_6871);
and U7478 (N_7478,N_6341,N_6794);
and U7479 (N_7479,N_6559,N_6098);
or U7480 (N_7480,N_6275,N_6591);
and U7481 (N_7481,N_6962,N_6977);
nand U7482 (N_7482,N_6119,N_6900);
and U7483 (N_7483,N_6248,N_6813);
nor U7484 (N_7484,N_6178,N_6443);
nand U7485 (N_7485,N_6183,N_6397);
and U7486 (N_7486,N_6110,N_6710);
and U7487 (N_7487,N_6198,N_6403);
nand U7488 (N_7488,N_6029,N_6013);
nor U7489 (N_7489,N_6913,N_6494);
nor U7490 (N_7490,N_6942,N_6310);
and U7491 (N_7491,N_6718,N_6070);
and U7492 (N_7492,N_6955,N_6870);
nand U7493 (N_7493,N_6712,N_6615);
nor U7494 (N_7494,N_6352,N_6297);
nor U7495 (N_7495,N_6996,N_6783);
nor U7496 (N_7496,N_6163,N_6414);
or U7497 (N_7497,N_6667,N_6698);
nor U7498 (N_7498,N_6311,N_6304);
nand U7499 (N_7499,N_6287,N_6791);
nor U7500 (N_7500,N_6170,N_6447);
or U7501 (N_7501,N_6047,N_6193);
nor U7502 (N_7502,N_6028,N_6525);
and U7503 (N_7503,N_6730,N_6775);
or U7504 (N_7504,N_6317,N_6422);
nor U7505 (N_7505,N_6756,N_6810);
or U7506 (N_7506,N_6522,N_6833);
xor U7507 (N_7507,N_6656,N_6405);
or U7508 (N_7508,N_6019,N_6231);
nor U7509 (N_7509,N_6969,N_6906);
or U7510 (N_7510,N_6439,N_6862);
or U7511 (N_7511,N_6317,N_6476);
or U7512 (N_7512,N_6634,N_6258);
nor U7513 (N_7513,N_6428,N_6783);
nor U7514 (N_7514,N_6756,N_6350);
or U7515 (N_7515,N_6967,N_6846);
or U7516 (N_7516,N_6386,N_6164);
nor U7517 (N_7517,N_6759,N_6622);
and U7518 (N_7518,N_6488,N_6870);
and U7519 (N_7519,N_6888,N_6326);
and U7520 (N_7520,N_6527,N_6621);
and U7521 (N_7521,N_6678,N_6469);
and U7522 (N_7522,N_6695,N_6419);
or U7523 (N_7523,N_6829,N_6327);
nor U7524 (N_7524,N_6399,N_6606);
nor U7525 (N_7525,N_6864,N_6839);
and U7526 (N_7526,N_6456,N_6205);
and U7527 (N_7527,N_6894,N_6084);
nand U7528 (N_7528,N_6685,N_6737);
and U7529 (N_7529,N_6404,N_6892);
nor U7530 (N_7530,N_6906,N_6102);
and U7531 (N_7531,N_6177,N_6082);
or U7532 (N_7532,N_6009,N_6714);
nand U7533 (N_7533,N_6783,N_6505);
or U7534 (N_7534,N_6133,N_6582);
nor U7535 (N_7535,N_6054,N_6208);
and U7536 (N_7536,N_6820,N_6627);
nor U7537 (N_7537,N_6841,N_6567);
or U7538 (N_7538,N_6516,N_6446);
and U7539 (N_7539,N_6296,N_6467);
or U7540 (N_7540,N_6640,N_6694);
nor U7541 (N_7541,N_6370,N_6112);
and U7542 (N_7542,N_6199,N_6201);
nand U7543 (N_7543,N_6884,N_6904);
nor U7544 (N_7544,N_6841,N_6935);
nor U7545 (N_7545,N_6606,N_6669);
or U7546 (N_7546,N_6198,N_6646);
nand U7547 (N_7547,N_6784,N_6084);
xnor U7548 (N_7548,N_6058,N_6644);
nand U7549 (N_7549,N_6005,N_6190);
or U7550 (N_7550,N_6929,N_6298);
nand U7551 (N_7551,N_6202,N_6658);
and U7552 (N_7552,N_6917,N_6450);
nor U7553 (N_7553,N_6655,N_6977);
or U7554 (N_7554,N_6179,N_6646);
and U7555 (N_7555,N_6383,N_6176);
nand U7556 (N_7556,N_6224,N_6387);
nand U7557 (N_7557,N_6982,N_6732);
or U7558 (N_7558,N_6011,N_6178);
and U7559 (N_7559,N_6411,N_6603);
nand U7560 (N_7560,N_6911,N_6061);
nor U7561 (N_7561,N_6332,N_6383);
and U7562 (N_7562,N_6183,N_6236);
and U7563 (N_7563,N_6749,N_6621);
nand U7564 (N_7564,N_6930,N_6520);
and U7565 (N_7565,N_6630,N_6890);
and U7566 (N_7566,N_6173,N_6417);
nand U7567 (N_7567,N_6249,N_6658);
xnor U7568 (N_7568,N_6717,N_6557);
or U7569 (N_7569,N_6254,N_6938);
or U7570 (N_7570,N_6602,N_6559);
and U7571 (N_7571,N_6897,N_6151);
nand U7572 (N_7572,N_6838,N_6574);
and U7573 (N_7573,N_6244,N_6156);
nor U7574 (N_7574,N_6900,N_6150);
or U7575 (N_7575,N_6785,N_6240);
and U7576 (N_7576,N_6957,N_6844);
nor U7577 (N_7577,N_6249,N_6956);
or U7578 (N_7578,N_6235,N_6398);
xnor U7579 (N_7579,N_6239,N_6593);
or U7580 (N_7580,N_6459,N_6284);
and U7581 (N_7581,N_6964,N_6903);
nand U7582 (N_7582,N_6720,N_6261);
nor U7583 (N_7583,N_6309,N_6976);
nor U7584 (N_7584,N_6703,N_6789);
xnor U7585 (N_7585,N_6373,N_6095);
nand U7586 (N_7586,N_6318,N_6061);
nor U7587 (N_7587,N_6943,N_6031);
and U7588 (N_7588,N_6887,N_6513);
and U7589 (N_7589,N_6488,N_6682);
or U7590 (N_7590,N_6901,N_6862);
nand U7591 (N_7591,N_6237,N_6759);
nand U7592 (N_7592,N_6413,N_6400);
and U7593 (N_7593,N_6990,N_6945);
nor U7594 (N_7594,N_6922,N_6160);
or U7595 (N_7595,N_6049,N_6759);
nand U7596 (N_7596,N_6275,N_6889);
nor U7597 (N_7597,N_6007,N_6027);
nand U7598 (N_7598,N_6756,N_6424);
nor U7599 (N_7599,N_6742,N_6558);
and U7600 (N_7600,N_6905,N_6415);
or U7601 (N_7601,N_6969,N_6467);
nand U7602 (N_7602,N_6284,N_6736);
or U7603 (N_7603,N_6447,N_6937);
nand U7604 (N_7604,N_6387,N_6852);
xnor U7605 (N_7605,N_6015,N_6848);
or U7606 (N_7606,N_6894,N_6127);
nand U7607 (N_7607,N_6395,N_6217);
or U7608 (N_7608,N_6052,N_6622);
and U7609 (N_7609,N_6416,N_6209);
and U7610 (N_7610,N_6621,N_6189);
nor U7611 (N_7611,N_6477,N_6387);
nor U7612 (N_7612,N_6842,N_6810);
nand U7613 (N_7613,N_6857,N_6519);
and U7614 (N_7614,N_6197,N_6029);
nor U7615 (N_7615,N_6222,N_6477);
nor U7616 (N_7616,N_6502,N_6240);
nand U7617 (N_7617,N_6433,N_6629);
nand U7618 (N_7618,N_6449,N_6257);
or U7619 (N_7619,N_6259,N_6064);
nand U7620 (N_7620,N_6130,N_6624);
nand U7621 (N_7621,N_6321,N_6257);
nor U7622 (N_7622,N_6261,N_6213);
and U7623 (N_7623,N_6999,N_6902);
nand U7624 (N_7624,N_6180,N_6962);
and U7625 (N_7625,N_6733,N_6434);
nor U7626 (N_7626,N_6036,N_6046);
and U7627 (N_7627,N_6971,N_6666);
and U7628 (N_7628,N_6242,N_6548);
or U7629 (N_7629,N_6207,N_6859);
or U7630 (N_7630,N_6322,N_6053);
or U7631 (N_7631,N_6813,N_6545);
xor U7632 (N_7632,N_6325,N_6481);
and U7633 (N_7633,N_6774,N_6587);
nand U7634 (N_7634,N_6505,N_6400);
nor U7635 (N_7635,N_6542,N_6778);
or U7636 (N_7636,N_6475,N_6431);
nor U7637 (N_7637,N_6836,N_6294);
or U7638 (N_7638,N_6501,N_6996);
or U7639 (N_7639,N_6928,N_6284);
or U7640 (N_7640,N_6530,N_6113);
and U7641 (N_7641,N_6635,N_6698);
nand U7642 (N_7642,N_6477,N_6780);
nor U7643 (N_7643,N_6724,N_6074);
xnor U7644 (N_7644,N_6886,N_6451);
and U7645 (N_7645,N_6827,N_6802);
nor U7646 (N_7646,N_6126,N_6395);
nor U7647 (N_7647,N_6110,N_6252);
nand U7648 (N_7648,N_6206,N_6678);
or U7649 (N_7649,N_6645,N_6588);
or U7650 (N_7650,N_6078,N_6706);
or U7651 (N_7651,N_6143,N_6485);
or U7652 (N_7652,N_6351,N_6118);
nor U7653 (N_7653,N_6239,N_6695);
nand U7654 (N_7654,N_6591,N_6457);
nand U7655 (N_7655,N_6943,N_6011);
or U7656 (N_7656,N_6033,N_6938);
and U7657 (N_7657,N_6579,N_6155);
xnor U7658 (N_7658,N_6308,N_6543);
or U7659 (N_7659,N_6924,N_6222);
and U7660 (N_7660,N_6808,N_6722);
and U7661 (N_7661,N_6834,N_6181);
and U7662 (N_7662,N_6616,N_6569);
or U7663 (N_7663,N_6012,N_6926);
or U7664 (N_7664,N_6417,N_6342);
and U7665 (N_7665,N_6716,N_6587);
and U7666 (N_7666,N_6293,N_6372);
or U7667 (N_7667,N_6034,N_6601);
nor U7668 (N_7668,N_6731,N_6802);
nor U7669 (N_7669,N_6851,N_6015);
nor U7670 (N_7670,N_6208,N_6510);
and U7671 (N_7671,N_6075,N_6499);
nand U7672 (N_7672,N_6011,N_6669);
and U7673 (N_7673,N_6113,N_6177);
or U7674 (N_7674,N_6276,N_6850);
nand U7675 (N_7675,N_6240,N_6706);
or U7676 (N_7676,N_6005,N_6179);
or U7677 (N_7677,N_6595,N_6888);
and U7678 (N_7678,N_6873,N_6693);
nor U7679 (N_7679,N_6933,N_6882);
and U7680 (N_7680,N_6097,N_6257);
or U7681 (N_7681,N_6357,N_6738);
and U7682 (N_7682,N_6541,N_6842);
nand U7683 (N_7683,N_6887,N_6748);
nand U7684 (N_7684,N_6630,N_6418);
nor U7685 (N_7685,N_6950,N_6318);
nand U7686 (N_7686,N_6729,N_6021);
nor U7687 (N_7687,N_6201,N_6093);
and U7688 (N_7688,N_6062,N_6146);
or U7689 (N_7689,N_6901,N_6133);
nand U7690 (N_7690,N_6618,N_6749);
nor U7691 (N_7691,N_6435,N_6708);
or U7692 (N_7692,N_6992,N_6871);
or U7693 (N_7693,N_6536,N_6843);
nand U7694 (N_7694,N_6103,N_6569);
nand U7695 (N_7695,N_6693,N_6824);
nor U7696 (N_7696,N_6022,N_6677);
nand U7697 (N_7697,N_6677,N_6643);
xnor U7698 (N_7698,N_6358,N_6605);
nor U7699 (N_7699,N_6282,N_6320);
nand U7700 (N_7700,N_6365,N_6858);
and U7701 (N_7701,N_6296,N_6914);
nand U7702 (N_7702,N_6312,N_6981);
and U7703 (N_7703,N_6545,N_6282);
or U7704 (N_7704,N_6672,N_6318);
nand U7705 (N_7705,N_6643,N_6971);
nand U7706 (N_7706,N_6836,N_6899);
nand U7707 (N_7707,N_6884,N_6620);
or U7708 (N_7708,N_6409,N_6622);
or U7709 (N_7709,N_6125,N_6867);
and U7710 (N_7710,N_6970,N_6403);
and U7711 (N_7711,N_6137,N_6705);
and U7712 (N_7712,N_6421,N_6062);
nor U7713 (N_7713,N_6744,N_6941);
nor U7714 (N_7714,N_6381,N_6732);
nand U7715 (N_7715,N_6706,N_6144);
or U7716 (N_7716,N_6167,N_6555);
nor U7717 (N_7717,N_6133,N_6964);
nand U7718 (N_7718,N_6249,N_6617);
and U7719 (N_7719,N_6841,N_6610);
nor U7720 (N_7720,N_6166,N_6353);
nor U7721 (N_7721,N_6423,N_6633);
and U7722 (N_7722,N_6315,N_6319);
xnor U7723 (N_7723,N_6246,N_6452);
nand U7724 (N_7724,N_6230,N_6758);
nand U7725 (N_7725,N_6509,N_6081);
or U7726 (N_7726,N_6115,N_6045);
nor U7727 (N_7727,N_6043,N_6151);
nor U7728 (N_7728,N_6572,N_6419);
and U7729 (N_7729,N_6743,N_6168);
nand U7730 (N_7730,N_6782,N_6857);
nor U7731 (N_7731,N_6609,N_6855);
nand U7732 (N_7732,N_6293,N_6863);
or U7733 (N_7733,N_6811,N_6196);
nor U7734 (N_7734,N_6681,N_6378);
nor U7735 (N_7735,N_6045,N_6183);
nor U7736 (N_7736,N_6721,N_6222);
or U7737 (N_7737,N_6613,N_6411);
nor U7738 (N_7738,N_6779,N_6042);
and U7739 (N_7739,N_6051,N_6673);
nor U7740 (N_7740,N_6512,N_6173);
and U7741 (N_7741,N_6027,N_6084);
or U7742 (N_7742,N_6745,N_6220);
nand U7743 (N_7743,N_6542,N_6588);
nand U7744 (N_7744,N_6092,N_6404);
and U7745 (N_7745,N_6173,N_6070);
nand U7746 (N_7746,N_6542,N_6835);
nor U7747 (N_7747,N_6019,N_6790);
nand U7748 (N_7748,N_6018,N_6780);
nor U7749 (N_7749,N_6735,N_6114);
nand U7750 (N_7750,N_6319,N_6089);
or U7751 (N_7751,N_6144,N_6007);
nor U7752 (N_7752,N_6519,N_6297);
and U7753 (N_7753,N_6061,N_6519);
and U7754 (N_7754,N_6010,N_6035);
nand U7755 (N_7755,N_6343,N_6868);
or U7756 (N_7756,N_6199,N_6047);
or U7757 (N_7757,N_6942,N_6597);
nor U7758 (N_7758,N_6062,N_6708);
nand U7759 (N_7759,N_6381,N_6837);
and U7760 (N_7760,N_6963,N_6189);
nor U7761 (N_7761,N_6088,N_6074);
nand U7762 (N_7762,N_6763,N_6503);
nand U7763 (N_7763,N_6741,N_6064);
nand U7764 (N_7764,N_6661,N_6594);
and U7765 (N_7765,N_6421,N_6201);
and U7766 (N_7766,N_6955,N_6106);
nand U7767 (N_7767,N_6259,N_6830);
nor U7768 (N_7768,N_6672,N_6555);
nor U7769 (N_7769,N_6371,N_6865);
nand U7770 (N_7770,N_6231,N_6095);
nand U7771 (N_7771,N_6479,N_6606);
or U7772 (N_7772,N_6370,N_6859);
nand U7773 (N_7773,N_6553,N_6060);
and U7774 (N_7774,N_6707,N_6770);
nor U7775 (N_7775,N_6745,N_6052);
and U7776 (N_7776,N_6957,N_6281);
or U7777 (N_7777,N_6949,N_6883);
and U7778 (N_7778,N_6539,N_6779);
nand U7779 (N_7779,N_6430,N_6893);
and U7780 (N_7780,N_6609,N_6540);
and U7781 (N_7781,N_6042,N_6795);
nor U7782 (N_7782,N_6398,N_6144);
and U7783 (N_7783,N_6855,N_6267);
and U7784 (N_7784,N_6105,N_6745);
or U7785 (N_7785,N_6443,N_6004);
nand U7786 (N_7786,N_6304,N_6983);
nand U7787 (N_7787,N_6451,N_6613);
and U7788 (N_7788,N_6945,N_6400);
nand U7789 (N_7789,N_6735,N_6871);
nand U7790 (N_7790,N_6706,N_6683);
and U7791 (N_7791,N_6053,N_6965);
nor U7792 (N_7792,N_6750,N_6982);
nor U7793 (N_7793,N_6728,N_6340);
nand U7794 (N_7794,N_6629,N_6971);
nand U7795 (N_7795,N_6489,N_6184);
and U7796 (N_7796,N_6429,N_6990);
nor U7797 (N_7797,N_6896,N_6193);
nand U7798 (N_7798,N_6288,N_6944);
nor U7799 (N_7799,N_6686,N_6785);
nor U7800 (N_7800,N_6034,N_6113);
or U7801 (N_7801,N_6113,N_6397);
nand U7802 (N_7802,N_6435,N_6215);
or U7803 (N_7803,N_6277,N_6789);
or U7804 (N_7804,N_6138,N_6312);
nand U7805 (N_7805,N_6263,N_6108);
and U7806 (N_7806,N_6889,N_6478);
nand U7807 (N_7807,N_6975,N_6052);
nand U7808 (N_7808,N_6059,N_6896);
or U7809 (N_7809,N_6736,N_6632);
and U7810 (N_7810,N_6626,N_6893);
and U7811 (N_7811,N_6265,N_6474);
nand U7812 (N_7812,N_6517,N_6104);
or U7813 (N_7813,N_6814,N_6033);
nor U7814 (N_7814,N_6991,N_6835);
or U7815 (N_7815,N_6683,N_6461);
nand U7816 (N_7816,N_6361,N_6384);
nor U7817 (N_7817,N_6372,N_6274);
nor U7818 (N_7818,N_6117,N_6491);
nand U7819 (N_7819,N_6247,N_6533);
or U7820 (N_7820,N_6134,N_6318);
and U7821 (N_7821,N_6502,N_6102);
nand U7822 (N_7822,N_6043,N_6720);
nor U7823 (N_7823,N_6638,N_6504);
and U7824 (N_7824,N_6469,N_6827);
or U7825 (N_7825,N_6957,N_6252);
nor U7826 (N_7826,N_6780,N_6981);
and U7827 (N_7827,N_6321,N_6620);
nor U7828 (N_7828,N_6849,N_6455);
or U7829 (N_7829,N_6141,N_6671);
nand U7830 (N_7830,N_6464,N_6104);
nor U7831 (N_7831,N_6673,N_6167);
nor U7832 (N_7832,N_6892,N_6981);
xor U7833 (N_7833,N_6701,N_6918);
or U7834 (N_7834,N_6454,N_6994);
and U7835 (N_7835,N_6207,N_6633);
and U7836 (N_7836,N_6012,N_6386);
nand U7837 (N_7837,N_6147,N_6776);
nand U7838 (N_7838,N_6232,N_6425);
nand U7839 (N_7839,N_6945,N_6658);
nand U7840 (N_7840,N_6003,N_6020);
and U7841 (N_7841,N_6786,N_6410);
nor U7842 (N_7842,N_6733,N_6838);
or U7843 (N_7843,N_6073,N_6072);
and U7844 (N_7844,N_6973,N_6345);
nor U7845 (N_7845,N_6282,N_6021);
nor U7846 (N_7846,N_6165,N_6022);
xor U7847 (N_7847,N_6694,N_6372);
nor U7848 (N_7848,N_6465,N_6219);
or U7849 (N_7849,N_6813,N_6071);
nand U7850 (N_7850,N_6346,N_6988);
nor U7851 (N_7851,N_6298,N_6838);
and U7852 (N_7852,N_6944,N_6514);
nand U7853 (N_7853,N_6529,N_6669);
nand U7854 (N_7854,N_6730,N_6940);
and U7855 (N_7855,N_6612,N_6774);
and U7856 (N_7856,N_6640,N_6057);
or U7857 (N_7857,N_6744,N_6170);
nand U7858 (N_7858,N_6656,N_6835);
nand U7859 (N_7859,N_6653,N_6676);
nor U7860 (N_7860,N_6602,N_6066);
nor U7861 (N_7861,N_6911,N_6426);
and U7862 (N_7862,N_6562,N_6575);
nor U7863 (N_7863,N_6836,N_6276);
or U7864 (N_7864,N_6480,N_6737);
nor U7865 (N_7865,N_6120,N_6565);
nand U7866 (N_7866,N_6255,N_6284);
or U7867 (N_7867,N_6675,N_6785);
nand U7868 (N_7868,N_6599,N_6992);
nand U7869 (N_7869,N_6843,N_6427);
or U7870 (N_7870,N_6559,N_6633);
nand U7871 (N_7871,N_6337,N_6905);
nand U7872 (N_7872,N_6894,N_6324);
xor U7873 (N_7873,N_6256,N_6261);
nor U7874 (N_7874,N_6354,N_6653);
nand U7875 (N_7875,N_6807,N_6189);
and U7876 (N_7876,N_6148,N_6556);
or U7877 (N_7877,N_6564,N_6795);
or U7878 (N_7878,N_6651,N_6892);
nand U7879 (N_7879,N_6401,N_6567);
nand U7880 (N_7880,N_6525,N_6547);
or U7881 (N_7881,N_6510,N_6534);
nor U7882 (N_7882,N_6099,N_6891);
nor U7883 (N_7883,N_6911,N_6188);
nor U7884 (N_7884,N_6154,N_6457);
and U7885 (N_7885,N_6374,N_6476);
and U7886 (N_7886,N_6818,N_6764);
nor U7887 (N_7887,N_6720,N_6330);
or U7888 (N_7888,N_6778,N_6861);
or U7889 (N_7889,N_6938,N_6697);
or U7890 (N_7890,N_6763,N_6769);
nor U7891 (N_7891,N_6136,N_6202);
or U7892 (N_7892,N_6849,N_6833);
and U7893 (N_7893,N_6559,N_6483);
or U7894 (N_7894,N_6109,N_6202);
nand U7895 (N_7895,N_6089,N_6995);
nor U7896 (N_7896,N_6020,N_6436);
or U7897 (N_7897,N_6635,N_6976);
and U7898 (N_7898,N_6350,N_6481);
nor U7899 (N_7899,N_6300,N_6521);
nand U7900 (N_7900,N_6173,N_6251);
nand U7901 (N_7901,N_6675,N_6584);
and U7902 (N_7902,N_6125,N_6815);
nand U7903 (N_7903,N_6889,N_6304);
nand U7904 (N_7904,N_6714,N_6330);
or U7905 (N_7905,N_6475,N_6630);
or U7906 (N_7906,N_6153,N_6718);
nand U7907 (N_7907,N_6281,N_6093);
nor U7908 (N_7908,N_6561,N_6880);
or U7909 (N_7909,N_6776,N_6619);
or U7910 (N_7910,N_6934,N_6383);
nor U7911 (N_7911,N_6200,N_6785);
nor U7912 (N_7912,N_6084,N_6376);
or U7913 (N_7913,N_6769,N_6268);
nand U7914 (N_7914,N_6447,N_6661);
and U7915 (N_7915,N_6055,N_6312);
and U7916 (N_7916,N_6420,N_6881);
xnor U7917 (N_7917,N_6342,N_6591);
nor U7918 (N_7918,N_6660,N_6489);
or U7919 (N_7919,N_6237,N_6339);
and U7920 (N_7920,N_6262,N_6103);
nand U7921 (N_7921,N_6721,N_6567);
and U7922 (N_7922,N_6578,N_6745);
nand U7923 (N_7923,N_6517,N_6250);
nor U7924 (N_7924,N_6943,N_6003);
nand U7925 (N_7925,N_6485,N_6528);
nor U7926 (N_7926,N_6832,N_6186);
nand U7927 (N_7927,N_6947,N_6817);
and U7928 (N_7928,N_6614,N_6353);
nand U7929 (N_7929,N_6062,N_6952);
nor U7930 (N_7930,N_6817,N_6948);
nor U7931 (N_7931,N_6423,N_6217);
nand U7932 (N_7932,N_6286,N_6621);
nand U7933 (N_7933,N_6577,N_6724);
nand U7934 (N_7934,N_6378,N_6529);
and U7935 (N_7935,N_6259,N_6102);
or U7936 (N_7936,N_6681,N_6452);
xor U7937 (N_7937,N_6643,N_6943);
nor U7938 (N_7938,N_6026,N_6354);
nor U7939 (N_7939,N_6959,N_6558);
nand U7940 (N_7940,N_6685,N_6933);
or U7941 (N_7941,N_6057,N_6895);
nor U7942 (N_7942,N_6460,N_6082);
and U7943 (N_7943,N_6451,N_6620);
and U7944 (N_7944,N_6660,N_6757);
and U7945 (N_7945,N_6505,N_6532);
nand U7946 (N_7946,N_6131,N_6195);
and U7947 (N_7947,N_6674,N_6665);
nand U7948 (N_7948,N_6895,N_6562);
and U7949 (N_7949,N_6252,N_6498);
nand U7950 (N_7950,N_6530,N_6572);
or U7951 (N_7951,N_6326,N_6777);
and U7952 (N_7952,N_6641,N_6888);
or U7953 (N_7953,N_6952,N_6001);
nand U7954 (N_7954,N_6358,N_6096);
or U7955 (N_7955,N_6036,N_6753);
or U7956 (N_7956,N_6891,N_6538);
and U7957 (N_7957,N_6426,N_6628);
or U7958 (N_7958,N_6609,N_6476);
nand U7959 (N_7959,N_6622,N_6626);
nand U7960 (N_7960,N_6372,N_6538);
and U7961 (N_7961,N_6266,N_6922);
or U7962 (N_7962,N_6509,N_6647);
nand U7963 (N_7963,N_6488,N_6856);
nor U7964 (N_7964,N_6934,N_6150);
and U7965 (N_7965,N_6482,N_6056);
nand U7966 (N_7966,N_6202,N_6702);
and U7967 (N_7967,N_6533,N_6825);
or U7968 (N_7968,N_6079,N_6862);
and U7969 (N_7969,N_6667,N_6502);
nor U7970 (N_7970,N_6048,N_6640);
nand U7971 (N_7971,N_6847,N_6562);
or U7972 (N_7972,N_6398,N_6443);
nor U7973 (N_7973,N_6656,N_6636);
nand U7974 (N_7974,N_6370,N_6898);
nor U7975 (N_7975,N_6829,N_6584);
nand U7976 (N_7976,N_6758,N_6159);
and U7977 (N_7977,N_6955,N_6866);
nand U7978 (N_7978,N_6919,N_6502);
nand U7979 (N_7979,N_6315,N_6698);
nand U7980 (N_7980,N_6951,N_6851);
and U7981 (N_7981,N_6582,N_6202);
nand U7982 (N_7982,N_6230,N_6335);
and U7983 (N_7983,N_6894,N_6177);
nor U7984 (N_7984,N_6711,N_6460);
nand U7985 (N_7985,N_6027,N_6500);
and U7986 (N_7986,N_6247,N_6495);
or U7987 (N_7987,N_6404,N_6826);
nor U7988 (N_7988,N_6053,N_6704);
nor U7989 (N_7989,N_6694,N_6656);
nand U7990 (N_7990,N_6949,N_6249);
or U7991 (N_7991,N_6052,N_6751);
nand U7992 (N_7992,N_6029,N_6649);
nand U7993 (N_7993,N_6595,N_6956);
or U7994 (N_7994,N_6479,N_6931);
xor U7995 (N_7995,N_6097,N_6998);
nor U7996 (N_7996,N_6456,N_6701);
xnor U7997 (N_7997,N_6522,N_6194);
or U7998 (N_7998,N_6023,N_6755);
nor U7999 (N_7999,N_6304,N_6430);
or U8000 (N_8000,N_7877,N_7281);
nand U8001 (N_8001,N_7033,N_7099);
nor U8002 (N_8002,N_7773,N_7226);
xnor U8003 (N_8003,N_7752,N_7842);
nand U8004 (N_8004,N_7639,N_7674);
nor U8005 (N_8005,N_7107,N_7321);
or U8006 (N_8006,N_7136,N_7519);
and U8007 (N_8007,N_7860,N_7817);
nor U8008 (N_8008,N_7621,N_7022);
or U8009 (N_8009,N_7488,N_7935);
xnor U8010 (N_8010,N_7793,N_7010);
nor U8011 (N_8011,N_7125,N_7075);
xnor U8012 (N_8012,N_7482,N_7581);
and U8013 (N_8013,N_7004,N_7579);
nor U8014 (N_8014,N_7492,N_7953);
or U8015 (N_8015,N_7193,N_7098);
xor U8016 (N_8016,N_7027,N_7588);
and U8017 (N_8017,N_7006,N_7048);
or U8018 (N_8018,N_7376,N_7791);
nor U8019 (N_8019,N_7690,N_7316);
and U8020 (N_8020,N_7122,N_7065);
or U8021 (N_8021,N_7443,N_7744);
and U8022 (N_8022,N_7259,N_7218);
or U8023 (N_8023,N_7634,N_7982);
nand U8024 (N_8024,N_7625,N_7166);
or U8025 (N_8025,N_7780,N_7897);
nor U8026 (N_8026,N_7504,N_7445);
nor U8027 (N_8027,N_7540,N_7499);
or U8028 (N_8028,N_7464,N_7669);
nand U8029 (N_8029,N_7641,N_7180);
and U8030 (N_8030,N_7865,N_7238);
xor U8031 (N_8031,N_7542,N_7798);
and U8032 (N_8032,N_7350,N_7505);
or U8033 (N_8033,N_7570,N_7105);
and U8034 (N_8034,N_7264,N_7101);
nand U8035 (N_8035,N_7926,N_7260);
and U8036 (N_8036,N_7086,N_7450);
nor U8037 (N_8037,N_7196,N_7333);
nor U8038 (N_8038,N_7245,N_7383);
nor U8039 (N_8039,N_7841,N_7007);
nand U8040 (N_8040,N_7473,N_7361);
nor U8041 (N_8041,N_7267,N_7711);
nor U8042 (N_8042,N_7129,N_7262);
nor U8043 (N_8043,N_7019,N_7153);
nand U8044 (N_8044,N_7025,N_7544);
and U8045 (N_8045,N_7756,N_7591);
and U8046 (N_8046,N_7480,N_7633);
nor U8047 (N_8047,N_7269,N_7949);
and U8048 (N_8048,N_7572,N_7317);
nor U8049 (N_8049,N_7044,N_7991);
nand U8050 (N_8050,N_7379,N_7745);
or U8051 (N_8051,N_7067,N_7353);
xor U8052 (N_8052,N_7565,N_7697);
nor U8053 (N_8053,N_7425,N_7160);
or U8054 (N_8054,N_7394,N_7364);
nand U8055 (N_8055,N_7393,N_7093);
or U8056 (N_8056,N_7047,N_7617);
and U8057 (N_8057,N_7430,N_7973);
nor U8058 (N_8058,N_7543,N_7412);
nor U8059 (N_8059,N_7481,N_7679);
and U8060 (N_8060,N_7527,N_7681);
or U8061 (N_8061,N_7762,N_7085);
or U8062 (N_8062,N_7670,N_7867);
and U8063 (N_8063,N_7145,N_7718);
and U8064 (N_8064,N_7653,N_7904);
and U8065 (N_8065,N_7981,N_7700);
or U8066 (N_8066,N_7092,N_7408);
or U8067 (N_8067,N_7380,N_7323);
nand U8068 (N_8068,N_7233,N_7134);
or U8069 (N_8069,N_7255,N_7373);
nor U8070 (N_8070,N_7902,N_7395);
and U8071 (N_8071,N_7298,N_7120);
nor U8072 (N_8072,N_7785,N_7058);
nor U8073 (N_8073,N_7609,N_7080);
nor U8074 (N_8074,N_7636,N_7358);
and U8075 (N_8075,N_7137,N_7938);
xor U8076 (N_8076,N_7293,N_7546);
nand U8077 (N_8077,N_7606,N_7941);
nor U8078 (N_8078,N_7892,N_7231);
nor U8079 (N_8079,N_7875,N_7392);
nor U8080 (N_8080,N_7879,N_7371);
xnor U8081 (N_8081,N_7857,N_7154);
and U8082 (N_8082,N_7734,N_7534);
and U8083 (N_8083,N_7183,N_7169);
nor U8084 (N_8084,N_7549,N_7312);
nand U8085 (N_8085,N_7442,N_7776);
nor U8086 (N_8086,N_7195,N_7498);
or U8087 (N_8087,N_7348,N_7507);
nor U8088 (N_8088,N_7789,N_7405);
or U8089 (N_8089,N_7413,N_7403);
xor U8090 (N_8090,N_7934,N_7295);
nand U8091 (N_8091,N_7850,N_7557);
or U8092 (N_8092,N_7016,N_7208);
and U8093 (N_8093,N_7512,N_7763);
and U8094 (N_8094,N_7645,N_7626);
or U8095 (N_8095,N_7971,N_7320);
or U8096 (N_8096,N_7864,N_7937);
or U8097 (N_8097,N_7400,N_7620);
nor U8098 (N_8098,N_7191,N_7057);
nand U8099 (N_8099,N_7889,N_7123);
nor U8100 (N_8100,N_7873,N_7550);
or U8101 (N_8101,N_7747,N_7244);
nand U8102 (N_8102,N_7113,N_7571);
nor U8103 (N_8103,N_7034,N_7622);
or U8104 (N_8104,N_7087,N_7614);
and U8105 (N_8105,N_7787,N_7375);
and U8106 (N_8106,N_7777,N_7753);
and U8107 (N_8107,N_7040,N_7724);
nor U8108 (N_8108,N_7922,N_7294);
nor U8109 (N_8109,N_7829,N_7503);
nor U8110 (N_8110,N_7150,N_7899);
or U8111 (N_8111,N_7187,N_7852);
or U8112 (N_8112,N_7182,N_7732);
nand U8113 (N_8113,N_7174,N_7657);
nor U8114 (N_8114,N_7382,N_7849);
nor U8115 (N_8115,N_7627,N_7108);
nor U8116 (N_8116,N_7784,N_7460);
or U8117 (N_8117,N_7433,N_7906);
or U8118 (N_8118,N_7330,N_7802);
nor U8119 (N_8119,N_7055,N_7717);
and U8120 (N_8120,N_7215,N_7646);
nand U8121 (N_8121,N_7435,N_7476);
nand U8122 (N_8122,N_7801,N_7072);
nand U8123 (N_8123,N_7313,N_7429);
and U8124 (N_8124,N_7186,N_7288);
and U8125 (N_8125,N_7270,N_7794);
nand U8126 (N_8126,N_7073,N_7268);
nand U8127 (N_8127,N_7750,N_7306);
xor U8128 (N_8128,N_7835,N_7079);
nor U8129 (N_8129,N_7671,N_7173);
nand U8130 (N_8130,N_7969,N_7436);
and U8131 (N_8131,N_7035,N_7642);
xor U8132 (N_8132,N_7112,N_7453);
and U8133 (N_8133,N_7638,N_7538);
nand U8134 (N_8134,N_7685,N_7869);
and U8135 (N_8135,N_7924,N_7804);
nand U8136 (N_8136,N_7957,N_7109);
nand U8137 (N_8137,N_7962,N_7853);
and U8138 (N_8138,N_7847,N_7511);
and U8139 (N_8139,N_7910,N_7159);
and U8140 (N_8140,N_7952,N_7110);
nand U8141 (N_8141,N_7135,N_7983);
or U8142 (N_8142,N_7014,N_7738);
or U8143 (N_8143,N_7629,N_7607);
or U8144 (N_8144,N_7415,N_7918);
and U8145 (N_8145,N_7770,N_7165);
nor U8146 (N_8146,N_7372,N_7782);
or U8147 (N_8147,N_7644,N_7917);
nand U8148 (N_8148,N_7297,N_7664);
nand U8149 (N_8149,N_7525,N_7615);
and U8150 (N_8150,N_7018,N_7583);
nand U8151 (N_8151,N_7448,N_7603);
nor U8152 (N_8152,N_7526,N_7815);
nor U8153 (N_8153,N_7749,N_7198);
nand U8154 (N_8154,N_7469,N_7594);
nand U8155 (N_8155,N_7168,N_7999);
nand U8156 (N_8156,N_7494,N_7704);
nand U8157 (N_8157,N_7531,N_7903);
nor U8158 (N_8158,N_7733,N_7141);
and U8159 (N_8159,N_7530,N_7287);
or U8160 (N_8160,N_7363,N_7928);
nor U8161 (N_8161,N_7725,N_7199);
and U8162 (N_8162,N_7662,N_7828);
nand U8163 (N_8163,N_7727,N_7533);
nand U8164 (N_8164,N_7576,N_7339);
or U8165 (N_8165,N_7740,N_7343);
nand U8166 (N_8166,N_7529,N_7933);
nor U8167 (N_8167,N_7352,N_7030);
nor U8168 (N_8168,N_7508,N_7501);
and U8169 (N_8169,N_7387,N_7000);
nand U8170 (N_8170,N_7523,N_7901);
xor U8171 (N_8171,N_7291,N_7513);
or U8172 (N_8172,N_7795,N_7097);
nand U8173 (N_8173,N_7431,N_7568);
and U8174 (N_8174,N_7856,N_7487);
nor U8175 (N_8175,N_7552,N_7569);
and U8176 (N_8176,N_7694,N_7566);
nor U8177 (N_8177,N_7545,N_7822);
or U8178 (N_8178,N_7252,N_7739);
nand U8179 (N_8179,N_7623,N_7280);
nor U8180 (N_8180,N_7053,N_7536);
or U8181 (N_8181,N_7300,N_7219);
nand U8182 (N_8182,N_7471,N_7968);
nor U8183 (N_8183,N_7500,N_7032);
and U8184 (N_8184,N_7440,N_7462);
nor U8185 (N_8185,N_7585,N_7771);
or U8186 (N_8186,N_7673,N_7987);
and U8187 (N_8187,N_7106,N_7528);
nand U8188 (N_8188,N_7863,N_7289);
nand U8189 (N_8189,N_7781,N_7945);
or U8190 (N_8190,N_7986,N_7359);
nand U8191 (N_8191,N_7146,N_7386);
or U8192 (N_8192,N_7490,N_7021);
nor U8193 (N_8193,N_7551,N_7611);
and U8194 (N_8194,N_7043,N_7103);
nor U8195 (N_8195,N_7036,N_7455);
nand U8196 (N_8196,N_7950,N_7946);
xor U8197 (N_8197,N_7311,N_7742);
and U8198 (N_8198,N_7114,N_7334);
or U8199 (N_8199,N_7959,N_7161);
nand U8200 (N_8200,N_7329,N_7936);
and U8201 (N_8201,N_7305,N_7884);
nand U8202 (N_8202,N_7322,N_7369);
or U8203 (N_8203,N_7883,N_7063);
and U8204 (N_8204,N_7792,N_7223);
and U8205 (N_8205,N_7855,N_7825);
or U8206 (N_8206,N_7046,N_7827);
or U8207 (N_8207,N_7411,N_7596);
nor U8208 (N_8208,N_7558,N_7556);
nand U8209 (N_8209,N_7837,N_7144);
or U8210 (N_8210,N_7871,N_7374);
or U8211 (N_8211,N_7172,N_7489);
nor U8212 (N_8212,N_7211,N_7820);
and U8213 (N_8213,N_7824,N_7819);
xnor U8214 (N_8214,N_7894,N_7438);
nand U8215 (N_8215,N_7327,N_7002);
nor U8216 (N_8216,N_7302,N_7271);
and U8217 (N_8217,N_7060,N_7786);
nand U8218 (N_8218,N_7735,N_7351);
or U8219 (N_8219,N_7406,N_7630);
nand U8220 (N_8220,N_7520,N_7419);
nor U8221 (N_8221,N_7675,N_7265);
or U8222 (N_8222,N_7151,N_7595);
and U8223 (N_8223,N_7832,N_7273);
or U8224 (N_8224,N_7772,N_7128);
or U8225 (N_8225,N_7263,N_7020);
or U8226 (N_8226,N_7584,N_7992);
nand U8227 (N_8227,N_7722,N_7967);
and U8228 (N_8228,N_7993,N_7796);
nor U8229 (N_8229,N_7397,N_7456);
nor U8230 (N_8230,N_7524,N_7800);
or U8231 (N_8231,N_7672,N_7610);
nor U8232 (N_8232,N_7423,N_7390);
and U8233 (N_8233,N_7643,N_7064);
or U8234 (N_8234,N_7966,N_7315);
and U8235 (N_8235,N_7147,N_7447);
nor U8236 (N_8236,N_7619,N_7398);
and U8237 (N_8237,N_7241,N_7258);
nand U8238 (N_8238,N_7580,N_7831);
or U8239 (N_8239,N_7563,N_7844);
nor U8240 (N_8240,N_7342,N_7005);
nand U8241 (N_8241,N_7331,N_7723);
or U8242 (N_8242,N_7054,N_7424);
or U8243 (N_8243,N_7407,N_7517);
and U8244 (N_8244,N_7995,N_7931);
nand U8245 (N_8245,N_7203,N_7340);
and U8246 (N_8246,N_7078,N_7224);
or U8247 (N_8247,N_7111,N_7988);
and U8248 (N_8248,N_7806,N_7236);
or U8249 (N_8249,N_7495,N_7651);
and U8250 (N_8250,N_7071,N_7755);
or U8251 (N_8251,N_7923,N_7748);
or U8252 (N_8252,N_7421,N_7337);
and U8253 (N_8253,N_7309,N_7874);
and U8254 (N_8254,N_7332,N_7210);
or U8255 (N_8255,N_7731,N_7444);
and U8256 (N_8256,N_7721,N_7013);
and U8257 (N_8257,N_7197,N_7213);
xor U8258 (N_8258,N_7942,N_7391);
and U8259 (N_8259,N_7956,N_7285);
nand U8260 (N_8260,N_7848,N_7190);
and U8261 (N_8261,N_7497,N_7121);
or U8262 (N_8262,N_7384,N_7677);
or U8263 (N_8263,N_7457,N_7017);
or U8264 (N_8264,N_7207,N_7547);
and U8265 (N_8265,N_7009,N_7178);
xor U8266 (N_8266,N_7292,N_7091);
or U8267 (N_8267,N_7515,N_7710);
nor U8268 (N_8268,N_7929,N_7237);
or U8269 (N_8269,N_7314,N_7164);
or U8270 (N_8270,N_7227,N_7859);
nor U8271 (N_8271,N_7240,N_7761);
and U8272 (N_8272,N_7496,N_7921);
nor U8273 (N_8273,N_7729,N_7388);
and U8274 (N_8274,N_7077,N_7996);
nor U8275 (N_8275,N_7628,N_7247);
nor U8276 (N_8276,N_7417,N_7872);
or U8277 (N_8277,N_7024,N_7661);
nand U8278 (N_8278,N_7274,N_7676);
or U8279 (N_8279,N_7157,N_7362);
nor U8280 (N_8280,N_7713,N_7925);
or U8281 (N_8281,N_7360,N_7491);
nand U8282 (N_8282,N_7346,N_7900);
nor U8283 (N_8283,N_7728,N_7094);
or U8284 (N_8284,N_7913,N_7797);
and U8285 (N_8285,N_7881,N_7587);
xor U8286 (N_8286,N_7701,N_7712);
and U8287 (N_8287,N_7206,N_7814);
or U8288 (N_8288,N_7624,N_7858);
and U8289 (N_8289,N_7254,N_7600);
nor U8290 (N_8290,N_7344,N_7070);
or U8291 (N_8291,N_7175,N_7031);
xor U8292 (N_8292,N_7640,N_7148);
or U8293 (N_8293,N_7919,N_7308);
nand U8294 (N_8294,N_7011,N_7514);
nor U8295 (N_8295,N_7502,N_7582);
or U8296 (N_8296,N_7068,N_7809);
and U8297 (N_8297,N_7354,N_7483);
nand U8298 (N_8298,N_7970,N_7124);
or U8299 (N_8299,N_7188,N_7759);
xor U8300 (N_8300,N_7001,N_7783);
nor U8301 (N_8301,N_7652,N_7357);
and U8302 (N_8302,N_7414,N_7422);
nand U8303 (N_8303,N_7493,N_7458);
nor U8304 (N_8304,N_7960,N_7803);
nor U8305 (N_8305,N_7768,N_7083);
and U8306 (N_8306,N_7266,N_7807);
and U8307 (N_8307,N_7056,N_7702);
or U8308 (N_8308,N_7707,N_7714);
nand U8309 (N_8309,N_7909,N_7356);
or U8310 (N_8310,N_7696,N_7139);
nor U8311 (N_8311,N_7084,N_7911);
nor U8312 (N_8312,N_7866,N_7667);
and U8313 (N_8313,N_7632,N_7896);
and U8314 (N_8314,N_7251,N_7143);
or U8315 (N_8315,N_7746,N_7573);
and U8316 (N_8316,N_7862,N_7812);
and U8317 (N_8317,N_7541,N_7691);
nor U8318 (N_8318,N_7162,N_7730);
nor U8319 (N_8319,N_7979,N_7474);
nor U8320 (N_8320,N_7559,N_7846);
nor U8321 (N_8321,N_7076,N_7220);
or U8322 (N_8322,N_7066,N_7826);
and U8323 (N_8323,N_7402,N_7420);
and U8324 (N_8324,N_7840,N_7980);
and U8325 (N_8325,N_7916,N_7439);
nor U8326 (N_8326,N_7586,N_7604);
or U8327 (N_8327,N_7484,N_7680);
nor U8328 (N_8328,N_7659,N_7882);
or U8329 (N_8329,N_7049,N_7836);
nor U8330 (N_8330,N_7365,N_7574);
nor U8331 (N_8331,N_7564,N_7616);
nand U8332 (N_8332,N_7518,N_7194);
or U8333 (N_8333,N_7984,N_7880);
and U8334 (N_8334,N_7891,N_7324);
or U8335 (N_8335,N_7612,N_7449);
nand U8336 (N_8336,N_7296,N_7256);
nand U8337 (N_8337,N_7130,N_7041);
nand U8338 (N_8338,N_7964,N_7204);
and U8339 (N_8339,N_7061,N_7378);
nor U8340 (N_8340,N_7336,N_7234);
nand U8341 (N_8341,N_7318,N_7658);
nand U8342 (N_8342,N_7944,N_7286);
nor U8343 (N_8343,N_7301,N_7766);
or U8344 (N_8344,N_7039,N_7509);
nand U8345 (N_8345,N_7716,N_7663);
and U8346 (N_8346,N_7886,N_7149);
nand U8347 (N_8347,N_7965,N_7562);
and U8348 (N_8348,N_7216,N_7069);
nor U8349 (N_8349,N_7854,N_7242);
nand U8350 (N_8350,N_7142,N_7232);
or U8351 (N_8351,N_7341,N_7743);
nor U8352 (N_8352,N_7555,N_7834);
nor U8353 (N_8353,N_7184,N_7026);
nor U8354 (N_8354,N_7823,N_7920);
xor U8355 (N_8355,N_7279,N_7475);
or U8356 (N_8356,N_7290,N_7170);
nor U8357 (N_8357,N_7715,N_7805);
nand U8358 (N_8358,N_7905,N_7985);
and U8359 (N_8359,N_7765,N_7409);
and U8360 (N_8360,N_7126,N_7764);
nand U8361 (N_8361,N_7283,N_7467);
or U8362 (N_8362,N_7119,N_7654);
or U8363 (N_8363,N_7222,N_7775);
nand U8364 (N_8364,N_7441,N_7248);
or U8365 (N_8365,N_7736,N_7851);
nand U8366 (N_8366,N_7666,N_7808);
nand U8367 (N_8367,N_7635,N_7452);
nor U8368 (N_8368,N_7253,N_7947);
or U8369 (N_8369,N_7088,N_7319);
nand U8370 (N_8370,N_7045,N_7532);
nand U8371 (N_8371,N_7769,N_7235);
nand U8372 (N_8372,N_7389,N_7751);
or U8373 (N_8373,N_7876,N_7468);
nor U8374 (N_8374,N_7432,N_7131);
or U8375 (N_8375,N_7757,N_7593);
or U8376 (N_8376,N_7304,N_7209);
nand U8377 (N_8377,N_7156,N_7778);
nand U8378 (N_8378,N_7276,N_7217);
nand U8379 (N_8379,N_7939,N_7328);
and U8380 (N_8380,N_7972,N_7015);
or U8381 (N_8381,N_7096,N_7366);
and U8382 (N_8382,N_7486,N_7649);
and U8383 (N_8383,N_7192,N_7117);
nor U8384 (N_8384,N_7567,N_7102);
or U8385 (N_8385,N_7349,N_7385);
and U8386 (N_8386,N_7127,N_7012);
nand U8387 (N_8387,N_7246,N_7451);
nand U8388 (N_8388,N_7284,N_7930);
and U8389 (N_8389,N_7239,N_7185);
nor U8390 (N_8390,N_7401,N_7466);
nand U8391 (N_8391,N_7335,N_7212);
or U8392 (N_8392,N_7767,N_7741);
or U8393 (N_8393,N_7539,N_7278);
or U8394 (N_8394,N_7427,N_7648);
xnor U8395 (N_8395,N_7948,N_7228);
nand U8396 (N_8396,N_7709,N_7608);
nand U8397 (N_8397,N_7994,N_7958);
and U8398 (N_8398,N_7977,N_7310);
or U8399 (N_8399,N_7434,N_7325);
nand U8400 (N_8400,N_7152,N_7708);
and U8401 (N_8401,N_7760,N_7081);
nand U8402 (N_8402,N_7510,N_7838);
nor U8403 (N_8403,N_7578,N_7613);
and U8404 (N_8404,N_7221,N_7303);
and U8405 (N_8405,N_7693,N_7478);
or U8406 (N_8406,N_7818,N_7975);
or U8407 (N_8407,N_7368,N_7307);
nand U8408 (N_8408,N_7961,N_7575);
nor U8409 (N_8409,N_7100,N_7553);
and U8410 (N_8410,N_7779,N_7463);
or U8411 (N_8411,N_7446,N_7189);
nor U8412 (N_8412,N_7688,N_7684);
and U8413 (N_8413,N_7472,N_7963);
nor U8414 (N_8414,N_7868,N_7506);
and U8415 (N_8415,N_7163,N_7155);
nor U8416 (N_8416,N_7601,N_7116);
nor U8417 (N_8417,N_7890,N_7355);
and U8418 (N_8418,N_7465,N_7719);
and U8419 (N_8419,N_7907,N_7754);
or U8420 (N_8420,N_7454,N_7051);
and U8421 (N_8421,N_7181,N_7811);
nand U8422 (N_8422,N_7275,N_7590);
nor U8423 (N_8423,N_7915,N_7202);
and U8424 (N_8424,N_7370,N_7683);
or U8425 (N_8425,N_7133,N_7138);
and U8426 (N_8426,N_7179,N_7347);
and U8427 (N_8427,N_7790,N_7257);
or U8428 (N_8428,N_7416,N_7647);
or U8429 (N_8429,N_7665,N_7230);
nand U8430 (N_8430,N_7470,N_7655);
and U8431 (N_8431,N_7870,N_7229);
nor U8432 (N_8432,N_7706,N_7932);
nor U8433 (N_8433,N_7698,N_7059);
or U8434 (N_8434,N_7705,N_7176);
or U8435 (N_8435,N_7167,N_7261);
nor U8436 (N_8436,N_7656,N_7437);
or U8437 (N_8437,N_7023,N_7404);
nand U8438 (N_8438,N_7095,N_7893);
xor U8439 (N_8439,N_7477,N_7082);
nand U8440 (N_8440,N_7605,N_7479);
nand U8441 (N_8441,N_7177,N_7535);
nand U8442 (N_8442,N_7758,N_7214);
or U8443 (N_8443,N_7598,N_7720);
or U8444 (N_8444,N_7171,N_7861);
nand U8445 (N_8445,N_7887,N_7399);
nand U8446 (N_8446,N_7943,N_7272);
xor U8447 (N_8447,N_7816,N_7678);
nand U8448 (N_8448,N_7689,N_7998);
nor U8449 (N_8449,N_7833,N_7774);
nand U8450 (N_8450,N_7548,N_7074);
and U8451 (N_8451,N_7821,N_7885);
nor U8452 (N_8452,N_7845,N_7381);
nor U8453 (N_8453,N_7703,N_7990);
or U8454 (N_8454,N_7042,N_7345);
or U8455 (N_8455,N_7912,N_7997);
nor U8456 (N_8456,N_7660,N_7788);
nor U8457 (N_8457,N_7914,N_7249);
nor U8458 (N_8458,N_7602,N_7839);
and U8459 (N_8459,N_7459,N_7118);
nor U8460 (N_8460,N_7485,N_7560);
nand U8461 (N_8461,N_7686,N_7396);
or U8462 (N_8462,N_7277,N_7516);
or U8463 (N_8463,N_7682,N_7028);
and U8464 (N_8464,N_7989,N_7978);
nor U8465 (N_8465,N_7650,N_7089);
nor U8466 (N_8466,N_7940,N_7428);
nor U8467 (N_8467,N_7692,N_7726);
or U8468 (N_8468,N_7737,N_7599);
or U8469 (N_8469,N_7201,N_7461);
nor U8470 (N_8470,N_7050,N_7521);
nor U8471 (N_8471,N_7810,N_7299);
nor U8472 (N_8472,N_7687,N_7062);
and U8473 (N_8473,N_7813,N_7951);
or U8474 (N_8474,N_7898,N_7631);
nand U8475 (N_8475,N_7377,N_7104);
or U8476 (N_8476,N_7037,N_7200);
or U8477 (N_8477,N_7367,N_7843);
or U8478 (N_8478,N_7927,N_7637);
nor U8479 (N_8479,N_7250,N_7955);
and U8480 (N_8480,N_7132,N_7561);
and U8481 (N_8481,N_7976,N_7618);
and U8482 (N_8482,N_7954,N_7140);
nor U8483 (N_8483,N_7577,N_7537);
or U8484 (N_8484,N_7029,N_7830);
or U8485 (N_8485,N_7974,N_7418);
nand U8486 (N_8486,N_7426,N_7052);
xor U8487 (N_8487,N_7410,N_7888);
nor U8488 (N_8488,N_7158,N_7908);
nor U8489 (N_8489,N_7878,N_7592);
and U8490 (N_8490,N_7338,N_7225);
or U8491 (N_8491,N_7205,N_7003);
and U8492 (N_8492,N_7668,N_7115);
or U8493 (N_8493,N_7597,N_7243);
nor U8494 (N_8494,N_7326,N_7695);
nand U8495 (N_8495,N_7282,N_7799);
or U8496 (N_8496,N_7699,N_7589);
nor U8497 (N_8497,N_7038,N_7895);
and U8498 (N_8498,N_7008,N_7554);
nand U8499 (N_8499,N_7522,N_7090);
and U8500 (N_8500,N_7243,N_7324);
nor U8501 (N_8501,N_7607,N_7697);
nand U8502 (N_8502,N_7879,N_7049);
or U8503 (N_8503,N_7208,N_7379);
nand U8504 (N_8504,N_7597,N_7617);
and U8505 (N_8505,N_7690,N_7094);
nor U8506 (N_8506,N_7934,N_7595);
nor U8507 (N_8507,N_7738,N_7387);
nor U8508 (N_8508,N_7608,N_7100);
and U8509 (N_8509,N_7702,N_7803);
xor U8510 (N_8510,N_7859,N_7320);
nor U8511 (N_8511,N_7079,N_7392);
or U8512 (N_8512,N_7924,N_7942);
nand U8513 (N_8513,N_7245,N_7753);
and U8514 (N_8514,N_7379,N_7133);
nand U8515 (N_8515,N_7745,N_7905);
and U8516 (N_8516,N_7788,N_7747);
nand U8517 (N_8517,N_7298,N_7729);
or U8518 (N_8518,N_7438,N_7194);
or U8519 (N_8519,N_7026,N_7653);
nand U8520 (N_8520,N_7975,N_7948);
nor U8521 (N_8521,N_7552,N_7697);
and U8522 (N_8522,N_7641,N_7744);
and U8523 (N_8523,N_7172,N_7843);
nor U8524 (N_8524,N_7039,N_7672);
nor U8525 (N_8525,N_7474,N_7541);
nor U8526 (N_8526,N_7568,N_7920);
or U8527 (N_8527,N_7151,N_7301);
and U8528 (N_8528,N_7161,N_7159);
nor U8529 (N_8529,N_7667,N_7981);
nor U8530 (N_8530,N_7655,N_7029);
nor U8531 (N_8531,N_7932,N_7335);
nand U8532 (N_8532,N_7914,N_7941);
or U8533 (N_8533,N_7405,N_7392);
and U8534 (N_8534,N_7468,N_7776);
nand U8535 (N_8535,N_7578,N_7942);
or U8536 (N_8536,N_7369,N_7751);
nor U8537 (N_8537,N_7696,N_7156);
nor U8538 (N_8538,N_7131,N_7256);
and U8539 (N_8539,N_7561,N_7197);
nor U8540 (N_8540,N_7172,N_7102);
nor U8541 (N_8541,N_7543,N_7305);
nand U8542 (N_8542,N_7396,N_7622);
and U8543 (N_8543,N_7649,N_7091);
and U8544 (N_8544,N_7932,N_7785);
nand U8545 (N_8545,N_7315,N_7559);
nor U8546 (N_8546,N_7851,N_7240);
and U8547 (N_8547,N_7016,N_7422);
nor U8548 (N_8548,N_7181,N_7516);
xnor U8549 (N_8549,N_7052,N_7090);
and U8550 (N_8550,N_7640,N_7458);
and U8551 (N_8551,N_7924,N_7847);
nor U8552 (N_8552,N_7667,N_7799);
or U8553 (N_8553,N_7906,N_7589);
or U8554 (N_8554,N_7213,N_7122);
and U8555 (N_8555,N_7177,N_7028);
nor U8556 (N_8556,N_7616,N_7126);
and U8557 (N_8557,N_7261,N_7841);
nand U8558 (N_8558,N_7671,N_7006);
nand U8559 (N_8559,N_7201,N_7073);
nor U8560 (N_8560,N_7062,N_7116);
nand U8561 (N_8561,N_7764,N_7454);
nor U8562 (N_8562,N_7961,N_7826);
and U8563 (N_8563,N_7695,N_7342);
and U8564 (N_8564,N_7846,N_7084);
and U8565 (N_8565,N_7194,N_7945);
and U8566 (N_8566,N_7977,N_7215);
nor U8567 (N_8567,N_7902,N_7884);
nand U8568 (N_8568,N_7689,N_7604);
or U8569 (N_8569,N_7040,N_7011);
nand U8570 (N_8570,N_7919,N_7808);
nor U8571 (N_8571,N_7288,N_7683);
nand U8572 (N_8572,N_7057,N_7707);
nand U8573 (N_8573,N_7110,N_7043);
nand U8574 (N_8574,N_7105,N_7723);
or U8575 (N_8575,N_7457,N_7396);
nand U8576 (N_8576,N_7811,N_7420);
or U8577 (N_8577,N_7881,N_7351);
nand U8578 (N_8578,N_7609,N_7308);
nand U8579 (N_8579,N_7096,N_7160);
and U8580 (N_8580,N_7700,N_7176);
nor U8581 (N_8581,N_7721,N_7353);
nor U8582 (N_8582,N_7172,N_7319);
and U8583 (N_8583,N_7983,N_7524);
or U8584 (N_8584,N_7265,N_7695);
or U8585 (N_8585,N_7798,N_7447);
nor U8586 (N_8586,N_7763,N_7117);
nor U8587 (N_8587,N_7847,N_7512);
and U8588 (N_8588,N_7977,N_7699);
nor U8589 (N_8589,N_7805,N_7435);
and U8590 (N_8590,N_7780,N_7457);
or U8591 (N_8591,N_7304,N_7553);
nor U8592 (N_8592,N_7443,N_7845);
and U8593 (N_8593,N_7616,N_7257);
xnor U8594 (N_8594,N_7932,N_7280);
nor U8595 (N_8595,N_7565,N_7078);
or U8596 (N_8596,N_7046,N_7768);
nor U8597 (N_8597,N_7422,N_7819);
nor U8598 (N_8598,N_7658,N_7807);
nor U8599 (N_8599,N_7682,N_7892);
nor U8600 (N_8600,N_7882,N_7789);
xor U8601 (N_8601,N_7892,N_7165);
nand U8602 (N_8602,N_7675,N_7142);
and U8603 (N_8603,N_7022,N_7941);
nor U8604 (N_8604,N_7693,N_7200);
or U8605 (N_8605,N_7445,N_7227);
nor U8606 (N_8606,N_7310,N_7492);
or U8607 (N_8607,N_7241,N_7770);
and U8608 (N_8608,N_7270,N_7998);
nand U8609 (N_8609,N_7068,N_7444);
or U8610 (N_8610,N_7383,N_7881);
and U8611 (N_8611,N_7133,N_7911);
or U8612 (N_8612,N_7472,N_7254);
xor U8613 (N_8613,N_7186,N_7278);
or U8614 (N_8614,N_7275,N_7236);
and U8615 (N_8615,N_7459,N_7004);
nor U8616 (N_8616,N_7424,N_7777);
nand U8617 (N_8617,N_7883,N_7937);
nor U8618 (N_8618,N_7577,N_7506);
nand U8619 (N_8619,N_7889,N_7842);
and U8620 (N_8620,N_7760,N_7383);
or U8621 (N_8621,N_7169,N_7418);
or U8622 (N_8622,N_7681,N_7768);
and U8623 (N_8623,N_7523,N_7351);
nor U8624 (N_8624,N_7467,N_7457);
nand U8625 (N_8625,N_7156,N_7460);
nor U8626 (N_8626,N_7547,N_7952);
or U8627 (N_8627,N_7923,N_7112);
nor U8628 (N_8628,N_7852,N_7129);
nor U8629 (N_8629,N_7357,N_7077);
nand U8630 (N_8630,N_7024,N_7498);
or U8631 (N_8631,N_7185,N_7707);
and U8632 (N_8632,N_7260,N_7393);
nand U8633 (N_8633,N_7490,N_7022);
nor U8634 (N_8634,N_7120,N_7779);
nand U8635 (N_8635,N_7869,N_7739);
nor U8636 (N_8636,N_7151,N_7638);
and U8637 (N_8637,N_7374,N_7068);
nor U8638 (N_8638,N_7137,N_7259);
nor U8639 (N_8639,N_7656,N_7521);
and U8640 (N_8640,N_7348,N_7119);
nand U8641 (N_8641,N_7543,N_7858);
nor U8642 (N_8642,N_7523,N_7149);
nor U8643 (N_8643,N_7862,N_7524);
nor U8644 (N_8644,N_7816,N_7955);
nand U8645 (N_8645,N_7742,N_7171);
and U8646 (N_8646,N_7092,N_7720);
and U8647 (N_8647,N_7085,N_7611);
nand U8648 (N_8648,N_7630,N_7531);
nand U8649 (N_8649,N_7850,N_7885);
and U8650 (N_8650,N_7003,N_7544);
nor U8651 (N_8651,N_7850,N_7316);
nand U8652 (N_8652,N_7497,N_7527);
nor U8653 (N_8653,N_7367,N_7552);
nor U8654 (N_8654,N_7859,N_7949);
nand U8655 (N_8655,N_7820,N_7595);
nand U8656 (N_8656,N_7162,N_7247);
or U8657 (N_8657,N_7465,N_7765);
and U8658 (N_8658,N_7352,N_7314);
nor U8659 (N_8659,N_7499,N_7769);
and U8660 (N_8660,N_7294,N_7575);
xor U8661 (N_8661,N_7898,N_7696);
nor U8662 (N_8662,N_7159,N_7227);
or U8663 (N_8663,N_7191,N_7856);
nor U8664 (N_8664,N_7605,N_7210);
nand U8665 (N_8665,N_7696,N_7205);
nor U8666 (N_8666,N_7112,N_7313);
and U8667 (N_8667,N_7901,N_7254);
and U8668 (N_8668,N_7504,N_7215);
or U8669 (N_8669,N_7945,N_7101);
or U8670 (N_8670,N_7959,N_7440);
or U8671 (N_8671,N_7228,N_7549);
nor U8672 (N_8672,N_7582,N_7324);
and U8673 (N_8673,N_7610,N_7575);
and U8674 (N_8674,N_7496,N_7896);
nand U8675 (N_8675,N_7522,N_7152);
and U8676 (N_8676,N_7896,N_7095);
nor U8677 (N_8677,N_7183,N_7596);
nor U8678 (N_8678,N_7799,N_7570);
nand U8679 (N_8679,N_7058,N_7244);
and U8680 (N_8680,N_7764,N_7275);
nor U8681 (N_8681,N_7843,N_7116);
or U8682 (N_8682,N_7587,N_7905);
nand U8683 (N_8683,N_7444,N_7225);
or U8684 (N_8684,N_7905,N_7139);
nand U8685 (N_8685,N_7225,N_7323);
or U8686 (N_8686,N_7809,N_7949);
and U8687 (N_8687,N_7373,N_7729);
nand U8688 (N_8688,N_7355,N_7403);
or U8689 (N_8689,N_7800,N_7867);
nor U8690 (N_8690,N_7181,N_7603);
xnor U8691 (N_8691,N_7695,N_7509);
nor U8692 (N_8692,N_7061,N_7878);
and U8693 (N_8693,N_7240,N_7677);
nand U8694 (N_8694,N_7997,N_7171);
nand U8695 (N_8695,N_7600,N_7715);
and U8696 (N_8696,N_7701,N_7628);
and U8697 (N_8697,N_7512,N_7502);
and U8698 (N_8698,N_7102,N_7840);
and U8699 (N_8699,N_7018,N_7287);
nor U8700 (N_8700,N_7788,N_7306);
nand U8701 (N_8701,N_7704,N_7172);
and U8702 (N_8702,N_7718,N_7960);
nand U8703 (N_8703,N_7742,N_7766);
nand U8704 (N_8704,N_7309,N_7842);
nor U8705 (N_8705,N_7276,N_7779);
or U8706 (N_8706,N_7949,N_7883);
or U8707 (N_8707,N_7095,N_7664);
and U8708 (N_8708,N_7892,N_7418);
or U8709 (N_8709,N_7079,N_7732);
nor U8710 (N_8710,N_7502,N_7829);
nand U8711 (N_8711,N_7989,N_7287);
nor U8712 (N_8712,N_7068,N_7303);
or U8713 (N_8713,N_7210,N_7763);
and U8714 (N_8714,N_7494,N_7272);
nand U8715 (N_8715,N_7031,N_7088);
nor U8716 (N_8716,N_7741,N_7875);
or U8717 (N_8717,N_7948,N_7281);
and U8718 (N_8718,N_7863,N_7644);
nor U8719 (N_8719,N_7954,N_7810);
nor U8720 (N_8720,N_7849,N_7562);
nor U8721 (N_8721,N_7408,N_7163);
and U8722 (N_8722,N_7052,N_7482);
and U8723 (N_8723,N_7424,N_7477);
nor U8724 (N_8724,N_7244,N_7374);
nor U8725 (N_8725,N_7633,N_7572);
nand U8726 (N_8726,N_7233,N_7426);
nand U8727 (N_8727,N_7901,N_7128);
or U8728 (N_8728,N_7235,N_7915);
nor U8729 (N_8729,N_7083,N_7890);
nor U8730 (N_8730,N_7256,N_7412);
xnor U8731 (N_8731,N_7251,N_7148);
and U8732 (N_8732,N_7779,N_7713);
nand U8733 (N_8733,N_7136,N_7112);
xor U8734 (N_8734,N_7922,N_7526);
nand U8735 (N_8735,N_7966,N_7479);
nand U8736 (N_8736,N_7803,N_7646);
and U8737 (N_8737,N_7587,N_7559);
or U8738 (N_8738,N_7243,N_7974);
and U8739 (N_8739,N_7308,N_7043);
or U8740 (N_8740,N_7133,N_7264);
or U8741 (N_8741,N_7679,N_7323);
nor U8742 (N_8742,N_7769,N_7244);
or U8743 (N_8743,N_7173,N_7263);
nor U8744 (N_8744,N_7517,N_7189);
nand U8745 (N_8745,N_7191,N_7631);
or U8746 (N_8746,N_7152,N_7452);
or U8747 (N_8747,N_7120,N_7500);
or U8748 (N_8748,N_7354,N_7344);
nor U8749 (N_8749,N_7623,N_7727);
nor U8750 (N_8750,N_7407,N_7604);
nand U8751 (N_8751,N_7100,N_7947);
nand U8752 (N_8752,N_7798,N_7938);
nand U8753 (N_8753,N_7818,N_7104);
nor U8754 (N_8754,N_7458,N_7555);
or U8755 (N_8755,N_7814,N_7999);
or U8756 (N_8756,N_7853,N_7972);
xor U8757 (N_8757,N_7037,N_7903);
or U8758 (N_8758,N_7934,N_7769);
nor U8759 (N_8759,N_7679,N_7040);
or U8760 (N_8760,N_7525,N_7724);
or U8761 (N_8761,N_7373,N_7793);
nand U8762 (N_8762,N_7941,N_7281);
xnor U8763 (N_8763,N_7019,N_7846);
nor U8764 (N_8764,N_7473,N_7140);
and U8765 (N_8765,N_7505,N_7190);
nand U8766 (N_8766,N_7382,N_7710);
nor U8767 (N_8767,N_7597,N_7103);
or U8768 (N_8768,N_7853,N_7437);
and U8769 (N_8769,N_7092,N_7550);
or U8770 (N_8770,N_7652,N_7094);
nand U8771 (N_8771,N_7647,N_7893);
and U8772 (N_8772,N_7900,N_7674);
nand U8773 (N_8773,N_7431,N_7548);
nor U8774 (N_8774,N_7187,N_7658);
and U8775 (N_8775,N_7485,N_7111);
nand U8776 (N_8776,N_7154,N_7739);
xnor U8777 (N_8777,N_7659,N_7037);
nor U8778 (N_8778,N_7246,N_7017);
or U8779 (N_8779,N_7542,N_7941);
nor U8780 (N_8780,N_7701,N_7533);
nand U8781 (N_8781,N_7770,N_7069);
or U8782 (N_8782,N_7327,N_7484);
or U8783 (N_8783,N_7700,N_7556);
nor U8784 (N_8784,N_7732,N_7265);
and U8785 (N_8785,N_7467,N_7078);
nor U8786 (N_8786,N_7669,N_7783);
nand U8787 (N_8787,N_7756,N_7315);
and U8788 (N_8788,N_7579,N_7048);
nor U8789 (N_8789,N_7707,N_7020);
and U8790 (N_8790,N_7238,N_7202);
or U8791 (N_8791,N_7172,N_7765);
or U8792 (N_8792,N_7653,N_7356);
nand U8793 (N_8793,N_7889,N_7128);
or U8794 (N_8794,N_7542,N_7233);
nand U8795 (N_8795,N_7371,N_7768);
nor U8796 (N_8796,N_7451,N_7353);
or U8797 (N_8797,N_7758,N_7887);
nor U8798 (N_8798,N_7555,N_7690);
nor U8799 (N_8799,N_7692,N_7024);
or U8800 (N_8800,N_7792,N_7148);
and U8801 (N_8801,N_7488,N_7195);
nor U8802 (N_8802,N_7990,N_7878);
or U8803 (N_8803,N_7055,N_7757);
nand U8804 (N_8804,N_7014,N_7318);
nor U8805 (N_8805,N_7202,N_7303);
or U8806 (N_8806,N_7265,N_7982);
nand U8807 (N_8807,N_7354,N_7759);
and U8808 (N_8808,N_7074,N_7848);
or U8809 (N_8809,N_7394,N_7544);
nand U8810 (N_8810,N_7618,N_7726);
or U8811 (N_8811,N_7406,N_7084);
and U8812 (N_8812,N_7099,N_7388);
nand U8813 (N_8813,N_7045,N_7572);
and U8814 (N_8814,N_7868,N_7676);
nand U8815 (N_8815,N_7497,N_7735);
and U8816 (N_8816,N_7121,N_7124);
or U8817 (N_8817,N_7810,N_7212);
nand U8818 (N_8818,N_7209,N_7569);
nor U8819 (N_8819,N_7363,N_7811);
and U8820 (N_8820,N_7257,N_7031);
or U8821 (N_8821,N_7780,N_7852);
and U8822 (N_8822,N_7567,N_7847);
nor U8823 (N_8823,N_7779,N_7179);
and U8824 (N_8824,N_7018,N_7715);
or U8825 (N_8825,N_7264,N_7655);
or U8826 (N_8826,N_7361,N_7642);
xor U8827 (N_8827,N_7379,N_7897);
nand U8828 (N_8828,N_7296,N_7362);
nor U8829 (N_8829,N_7368,N_7038);
xor U8830 (N_8830,N_7462,N_7288);
and U8831 (N_8831,N_7830,N_7498);
nand U8832 (N_8832,N_7978,N_7065);
nand U8833 (N_8833,N_7510,N_7864);
xor U8834 (N_8834,N_7930,N_7135);
or U8835 (N_8835,N_7715,N_7733);
and U8836 (N_8836,N_7044,N_7182);
nand U8837 (N_8837,N_7097,N_7121);
and U8838 (N_8838,N_7591,N_7174);
nand U8839 (N_8839,N_7295,N_7365);
nor U8840 (N_8840,N_7504,N_7701);
nand U8841 (N_8841,N_7842,N_7284);
and U8842 (N_8842,N_7632,N_7149);
or U8843 (N_8843,N_7166,N_7713);
and U8844 (N_8844,N_7424,N_7746);
and U8845 (N_8845,N_7061,N_7697);
and U8846 (N_8846,N_7986,N_7858);
or U8847 (N_8847,N_7167,N_7807);
and U8848 (N_8848,N_7718,N_7162);
nand U8849 (N_8849,N_7842,N_7293);
nor U8850 (N_8850,N_7814,N_7764);
nand U8851 (N_8851,N_7974,N_7053);
nand U8852 (N_8852,N_7111,N_7920);
or U8853 (N_8853,N_7741,N_7706);
nor U8854 (N_8854,N_7354,N_7234);
nand U8855 (N_8855,N_7944,N_7737);
nand U8856 (N_8856,N_7641,N_7202);
and U8857 (N_8857,N_7858,N_7753);
or U8858 (N_8858,N_7653,N_7661);
nor U8859 (N_8859,N_7784,N_7213);
and U8860 (N_8860,N_7524,N_7385);
or U8861 (N_8861,N_7310,N_7937);
and U8862 (N_8862,N_7197,N_7953);
nand U8863 (N_8863,N_7692,N_7199);
and U8864 (N_8864,N_7548,N_7100);
or U8865 (N_8865,N_7685,N_7082);
and U8866 (N_8866,N_7211,N_7317);
or U8867 (N_8867,N_7831,N_7157);
and U8868 (N_8868,N_7133,N_7504);
and U8869 (N_8869,N_7050,N_7861);
or U8870 (N_8870,N_7265,N_7134);
nand U8871 (N_8871,N_7125,N_7570);
nor U8872 (N_8872,N_7609,N_7058);
nand U8873 (N_8873,N_7708,N_7359);
and U8874 (N_8874,N_7245,N_7345);
and U8875 (N_8875,N_7957,N_7836);
or U8876 (N_8876,N_7352,N_7794);
or U8877 (N_8877,N_7402,N_7964);
nand U8878 (N_8878,N_7898,N_7987);
nand U8879 (N_8879,N_7368,N_7245);
and U8880 (N_8880,N_7329,N_7668);
nor U8881 (N_8881,N_7945,N_7815);
nor U8882 (N_8882,N_7532,N_7484);
nand U8883 (N_8883,N_7557,N_7401);
xor U8884 (N_8884,N_7427,N_7957);
or U8885 (N_8885,N_7811,N_7789);
nand U8886 (N_8886,N_7339,N_7942);
nor U8887 (N_8887,N_7208,N_7204);
or U8888 (N_8888,N_7583,N_7122);
and U8889 (N_8889,N_7642,N_7910);
nor U8890 (N_8890,N_7216,N_7140);
or U8891 (N_8891,N_7647,N_7780);
nor U8892 (N_8892,N_7605,N_7511);
nor U8893 (N_8893,N_7462,N_7182);
nand U8894 (N_8894,N_7825,N_7443);
or U8895 (N_8895,N_7898,N_7421);
nor U8896 (N_8896,N_7794,N_7492);
nor U8897 (N_8897,N_7988,N_7311);
or U8898 (N_8898,N_7983,N_7477);
nor U8899 (N_8899,N_7045,N_7504);
or U8900 (N_8900,N_7771,N_7867);
nor U8901 (N_8901,N_7261,N_7471);
or U8902 (N_8902,N_7147,N_7334);
or U8903 (N_8903,N_7450,N_7626);
nand U8904 (N_8904,N_7853,N_7978);
nand U8905 (N_8905,N_7655,N_7543);
nor U8906 (N_8906,N_7225,N_7240);
or U8907 (N_8907,N_7374,N_7898);
nand U8908 (N_8908,N_7070,N_7180);
and U8909 (N_8909,N_7569,N_7912);
or U8910 (N_8910,N_7306,N_7079);
nor U8911 (N_8911,N_7090,N_7020);
and U8912 (N_8912,N_7931,N_7867);
nand U8913 (N_8913,N_7025,N_7545);
nand U8914 (N_8914,N_7913,N_7796);
and U8915 (N_8915,N_7065,N_7776);
nand U8916 (N_8916,N_7099,N_7249);
xor U8917 (N_8917,N_7486,N_7381);
nand U8918 (N_8918,N_7520,N_7912);
nand U8919 (N_8919,N_7697,N_7783);
or U8920 (N_8920,N_7177,N_7998);
nand U8921 (N_8921,N_7369,N_7414);
and U8922 (N_8922,N_7492,N_7520);
and U8923 (N_8923,N_7094,N_7471);
or U8924 (N_8924,N_7967,N_7554);
or U8925 (N_8925,N_7633,N_7715);
nand U8926 (N_8926,N_7783,N_7142);
nand U8927 (N_8927,N_7495,N_7659);
xor U8928 (N_8928,N_7453,N_7524);
or U8929 (N_8929,N_7994,N_7189);
nand U8930 (N_8930,N_7424,N_7268);
or U8931 (N_8931,N_7749,N_7465);
nor U8932 (N_8932,N_7300,N_7329);
nand U8933 (N_8933,N_7879,N_7490);
or U8934 (N_8934,N_7612,N_7630);
or U8935 (N_8935,N_7907,N_7675);
xnor U8936 (N_8936,N_7138,N_7375);
nand U8937 (N_8937,N_7524,N_7070);
nor U8938 (N_8938,N_7482,N_7528);
xor U8939 (N_8939,N_7186,N_7549);
nor U8940 (N_8940,N_7647,N_7592);
or U8941 (N_8941,N_7574,N_7842);
xor U8942 (N_8942,N_7113,N_7134);
xor U8943 (N_8943,N_7248,N_7389);
nand U8944 (N_8944,N_7573,N_7422);
xnor U8945 (N_8945,N_7800,N_7200);
nor U8946 (N_8946,N_7704,N_7260);
or U8947 (N_8947,N_7786,N_7770);
and U8948 (N_8948,N_7059,N_7404);
and U8949 (N_8949,N_7942,N_7770);
and U8950 (N_8950,N_7035,N_7232);
nor U8951 (N_8951,N_7220,N_7731);
nand U8952 (N_8952,N_7160,N_7284);
nand U8953 (N_8953,N_7802,N_7616);
nand U8954 (N_8954,N_7313,N_7670);
nor U8955 (N_8955,N_7369,N_7355);
and U8956 (N_8956,N_7827,N_7085);
nand U8957 (N_8957,N_7071,N_7555);
nand U8958 (N_8958,N_7503,N_7454);
or U8959 (N_8959,N_7633,N_7199);
nor U8960 (N_8960,N_7066,N_7963);
nor U8961 (N_8961,N_7848,N_7761);
or U8962 (N_8962,N_7072,N_7820);
nor U8963 (N_8963,N_7521,N_7923);
nor U8964 (N_8964,N_7046,N_7754);
nand U8965 (N_8965,N_7764,N_7944);
or U8966 (N_8966,N_7301,N_7804);
nand U8967 (N_8967,N_7623,N_7957);
or U8968 (N_8968,N_7534,N_7748);
nand U8969 (N_8969,N_7515,N_7967);
and U8970 (N_8970,N_7235,N_7048);
and U8971 (N_8971,N_7880,N_7330);
xor U8972 (N_8972,N_7199,N_7622);
nor U8973 (N_8973,N_7451,N_7817);
nand U8974 (N_8974,N_7255,N_7288);
nor U8975 (N_8975,N_7584,N_7344);
and U8976 (N_8976,N_7234,N_7509);
and U8977 (N_8977,N_7136,N_7834);
or U8978 (N_8978,N_7203,N_7011);
or U8979 (N_8979,N_7909,N_7170);
nand U8980 (N_8980,N_7224,N_7980);
nor U8981 (N_8981,N_7044,N_7642);
and U8982 (N_8982,N_7111,N_7671);
nand U8983 (N_8983,N_7708,N_7361);
nand U8984 (N_8984,N_7298,N_7475);
nand U8985 (N_8985,N_7313,N_7850);
xnor U8986 (N_8986,N_7959,N_7094);
nand U8987 (N_8987,N_7809,N_7891);
nor U8988 (N_8988,N_7937,N_7188);
and U8989 (N_8989,N_7606,N_7197);
nor U8990 (N_8990,N_7060,N_7425);
nor U8991 (N_8991,N_7386,N_7553);
and U8992 (N_8992,N_7082,N_7802);
and U8993 (N_8993,N_7621,N_7414);
and U8994 (N_8994,N_7249,N_7820);
and U8995 (N_8995,N_7196,N_7060);
or U8996 (N_8996,N_7513,N_7721);
and U8997 (N_8997,N_7039,N_7164);
nor U8998 (N_8998,N_7090,N_7515);
nand U8999 (N_8999,N_7233,N_7397);
nor U9000 (N_9000,N_8427,N_8769);
nand U9001 (N_9001,N_8091,N_8974);
and U9002 (N_9002,N_8824,N_8631);
nand U9003 (N_9003,N_8981,N_8584);
nand U9004 (N_9004,N_8661,N_8809);
nand U9005 (N_9005,N_8508,N_8927);
nand U9006 (N_9006,N_8172,N_8314);
nor U9007 (N_9007,N_8789,N_8212);
nor U9008 (N_9008,N_8840,N_8902);
nor U9009 (N_9009,N_8870,N_8005);
nor U9010 (N_9010,N_8796,N_8050);
nand U9011 (N_9011,N_8200,N_8422);
nor U9012 (N_9012,N_8669,N_8586);
and U9013 (N_9013,N_8764,N_8335);
and U9014 (N_9014,N_8272,N_8514);
nor U9015 (N_9015,N_8786,N_8419);
nand U9016 (N_9016,N_8821,N_8950);
and U9017 (N_9017,N_8806,N_8255);
nor U9018 (N_9018,N_8699,N_8955);
nor U9019 (N_9019,N_8531,N_8970);
or U9020 (N_9020,N_8663,N_8136);
nor U9021 (N_9021,N_8658,N_8767);
or U9022 (N_9022,N_8420,N_8532);
nand U9023 (N_9023,N_8834,N_8180);
or U9024 (N_9024,N_8073,N_8209);
or U9025 (N_9025,N_8889,N_8365);
and U9026 (N_9026,N_8791,N_8907);
nor U9027 (N_9027,N_8971,N_8553);
and U9028 (N_9028,N_8284,N_8718);
nand U9029 (N_9029,N_8910,N_8896);
nor U9030 (N_9030,N_8759,N_8009);
nor U9031 (N_9031,N_8224,N_8317);
and U9032 (N_9032,N_8129,N_8856);
or U9033 (N_9033,N_8758,N_8742);
or U9034 (N_9034,N_8497,N_8325);
or U9035 (N_9035,N_8347,N_8776);
nand U9036 (N_9036,N_8736,N_8096);
or U9037 (N_9037,N_8415,N_8277);
and U9038 (N_9038,N_8945,N_8318);
nand U9039 (N_9039,N_8559,N_8107);
or U9040 (N_9040,N_8310,N_8996);
nand U9041 (N_9041,N_8316,N_8703);
nor U9042 (N_9042,N_8743,N_8930);
nand U9043 (N_9043,N_8363,N_8299);
and U9044 (N_9044,N_8025,N_8720);
xnor U9045 (N_9045,N_8721,N_8991);
and U9046 (N_9046,N_8113,N_8590);
and U9047 (N_9047,N_8875,N_8218);
and U9048 (N_9048,N_8210,N_8751);
or U9049 (N_9049,N_8285,N_8067);
or U9050 (N_9050,N_8071,N_8510);
nand U9051 (N_9051,N_8587,N_8293);
or U9052 (N_9052,N_8802,N_8311);
or U9053 (N_9053,N_8903,N_8487);
or U9054 (N_9054,N_8561,N_8333);
or U9055 (N_9055,N_8213,N_8370);
nand U9056 (N_9056,N_8263,N_8203);
and U9057 (N_9057,N_8612,N_8810);
and U9058 (N_9058,N_8378,N_8577);
or U9059 (N_9059,N_8346,N_8269);
nor U9060 (N_9060,N_8504,N_8899);
and U9061 (N_9061,N_8600,N_8617);
or U9062 (N_9062,N_8949,N_8575);
and U9063 (N_9063,N_8079,N_8001);
and U9064 (N_9064,N_8126,N_8726);
xnor U9065 (N_9065,N_8215,N_8282);
or U9066 (N_9066,N_8053,N_8062);
and U9067 (N_9067,N_8946,N_8233);
nor U9068 (N_9068,N_8155,N_8622);
and U9069 (N_9069,N_8376,N_8765);
or U9070 (N_9070,N_8998,N_8529);
nor U9071 (N_9071,N_8602,N_8513);
nor U9072 (N_9072,N_8994,N_8092);
nand U9073 (N_9073,N_8020,N_8744);
and U9074 (N_9074,N_8516,N_8238);
nand U9075 (N_9075,N_8688,N_8740);
or U9076 (N_9076,N_8247,N_8175);
xnor U9077 (N_9077,N_8109,N_8165);
and U9078 (N_9078,N_8656,N_8579);
nor U9079 (N_9079,N_8519,N_8771);
and U9080 (N_9080,N_8623,N_8204);
nor U9081 (N_9081,N_8002,N_8094);
nand U9082 (N_9082,N_8029,N_8607);
nor U9083 (N_9083,N_8232,N_8156);
nor U9084 (N_9084,N_8312,N_8961);
nand U9085 (N_9085,N_8474,N_8413);
nor U9086 (N_9086,N_8326,N_8278);
or U9087 (N_9087,N_8800,N_8698);
nand U9088 (N_9088,N_8064,N_8489);
and U9089 (N_9089,N_8545,N_8716);
nand U9090 (N_9090,N_8676,N_8948);
nand U9091 (N_9091,N_8841,N_8815);
or U9092 (N_9092,N_8932,N_8491);
or U9093 (N_9093,N_8366,N_8249);
nand U9094 (N_9094,N_8801,N_8262);
nor U9095 (N_9095,N_8027,N_8259);
or U9096 (N_9096,N_8635,N_8547);
nor U9097 (N_9097,N_8443,N_8469);
nand U9098 (N_9098,N_8082,N_8056);
nand U9099 (N_9099,N_8343,N_8000);
nand U9100 (N_9100,N_8075,N_8616);
and U9101 (N_9101,N_8331,N_8681);
or U9102 (N_9102,N_8007,N_8844);
nor U9103 (N_9103,N_8294,N_8476);
or U9104 (N_9104,N_8756,N_8957);
xnor U9105 (N_9105,N_8832,N_8191);
and U9106 (N_9106,N_8395,N_8424);
and U9107 (N_9107,N_8624,N_8780);
or U9108 (N_9108,N_8076,N_8280);
nand U9109 (N_9109,N_8080,N_8013);
nor U9110 (N_9110,N_8749,N_8386);
nand U9111 (N_9111,N_8146,N_8015);
or U9112 (N_9112,N_8568,N_8403);
or U9113 (N_9113,N_8977,N_8863);
nand U9114 (N_9114,N_8201,N_8216);
nand U9115 (N_9115,N_8103,N_8120);
or U9116 (N_9116,N_8667,N_8308);
nand U9117 (N_9117,N_8918,N_8196);
nor U9118 (N_9118,N_8460,N_8535);
or U9119 (N_9119,N_8537,N_8660);
nor U9120 (N_9120,N_8900,N_8356);
or U9121 (N_9121,N_8055,N_8735);
xnor U9122 (N_9122,N_8410,N_8098);
nor U9123 (N_9123,N_8574,N_8913);
nand U9124 (N_9124,N_8620,N_8149);
nor U9125 (N_9125,N_8941,N_8708);
or U9126 (N_9126,N_8515,N_8412);
or U9127 (N_9127,N_8142,N_8604);
nor U9128 (N_9128,N_8954,N_8967);
or U9129 (N_9129,N_8929,N_8125);
nand U9130 (N_9130,N_8524,N_8633);
nor U9131 (N_9131,N_8659,N_8592);
and U9132 (N_9132,N_8234,N_8985);
nand U9133 (N_9133,N_8684,N_8045);
and U9134 (N_9134,N_8770,N_8421);
nor U9135 (N_9135,N_8122,N_8706);
and U9136 (N_9136,N_8244,N_8162);
nor U9137 (N_9137,N_8766,N_8391);
xnor U9138 (N_9138,N_8909,N_8017);
or U9139 (N_9139,N_8106,N_8795);
nor U9140 (N_9140,N_8322,N_8978);
nand U9141 (N_9141,N_8141,N_8748);
nand U9142 (N_9142,N_8127,N_8330);
nand U9143 (N_9143,N_8179,N_8812);
nand U9144 (N_9144,N_8836,N_8662);
nor U9145 (N_9145,N_8372,N_8338);
nand U9146 (N_9146,N_8042,N_8931);
and U9147 (N_9147,N_8072,N_8777);
and U9148 (N_9148,N_8199,N_8986);
nand U9149 (N_9149,N_8467,N_8148);
and U9150 (N_9150,N_8835,N_8747);
or U9151 (N_9151,N_8675,N_8406);
nand U9152 (N_9152,N_8598,N_8921);
xor U9153 (N_9153,N_8454,N_8774);
nor U9154 (N_9154,N_8176,N_8779);
or U9155 (N_9155,N_8193,N_8496);
and U9156 (N_9156,N_8580,N_8606);
nand U9157 (N_9157,N_8479,N_8341);
and U9158 (N_9158,N_8451,N_8868);
nor U9159 (N_9159,N_8446,N_8784);
nand U9160 (N_9160,N_8626,N_8034);
and U9161 (N_9161,N_8026,N_8628);
xor U9162 (N_9162,N_8845,N_8518);
nor U9163 (N_9163,N_8254,N_8827);
nor U9164 (N_9164,N_8066,N_8104);
nor U9165 (N_9165,N_8520,N_8543);
nand U9166 (N_9166,N_8150,N_8877);
nor U9167 (N_9167,N_8551,N_8936);
and U9168 (N_9168,N_8089,N_8274);
nor U9169 (N_9169,N_8905,N_8564);
and U9170 (N_9170,N_8151,N_8083);
or U9171 (N_9171,N_8345,N_8440);
nor U9172 (N_9172,N_8601,N_8118);
nor U9173 (N_9173,N_8677,N_8281);
or U9174 (N_9174,N_8997,N_8337);
or U9175 (N_9175,N_8359,N_8485);
and U9176 (N_9176,N_8980,N_8717);
nor U9177 (N_9177,N_8400,N_8320);
nor U9178 (N_9178,N_8283,N_8984);
or U9179 (N_9179,N_8471,N_8178);
and U9180 (N_9180,N_8527,N_8288);
or U9181 (N_9181,N_8396,N_8043);
or U9182 (N_9182,N_8492,N_8723);
and U9183 (N_9183,N_8682,N_8030);
nor U9184 (N_9184,N_8309,N_8384);
nand U9185 (N_9185,N_8292,N_8174);
or U9186 (N_9186,N_8890,N_8444);
or U9187 (N_9187,N_8933,N_8882);
or U9188 (N_9188,N_8379,N_8979);
or U9189 (N_9189,N_8214,N_8241);
or U9190 (N_9190,N_8762,N_8560);
nand U9191 (N_9191,N_8730,N_8227);
and U9192 (N_9192,N_8100,N_8021);
and U9193 (N_9193,N_8947,N_8158);
xnor U9194 (N_9194,N_8057,N_8582);
and U9195 (N_9195,N_8297,N_8298);
and U9196 (N_9196,N_8265,N_8854);
nor U9197 (N_9197,N_8867,N_8817);
nand U9198 (N_9198,N_8301,N_8495);
or U9199 (N_9199,N_8144,N_8138);
or U9200 (N_9200,N_8303,N_8431);
nor U9201 (N_9201,N_8194,N_8589);
xor U9202 (N_9202,N_8879,N_8585);
nand U9203 (N_9203,N_8432,N_8369);
nor U9204 (N_9204,N_8666,N_8975);
or U9205 (N_9205,N_8611,N_8028);
and U9206 (N_9206,N_8074,N_8869);
nand U9207 (N_9207,N_8047,N_8752);
and U9208 (N_9208,N_8862,N_8168);
nand U9209 (N_9209,N_8920,N_8457);
nor U9210 (N_9210,N_8459,N_8893);
nor U9211 (N_9211,N_8939,N_8135);
nand U9212 (N_9212,N_8099,N_8782);
or U9213 (N_9213,N_8368,N_8266);
or U9214 (N_9214,N_8501,N_8058);
and U9215 (N_9215,N_8694,N_8276);
and U9216 (N_9216,N_8576,N_8052);
nand U9217 (N_9217,N_8897,N_8943);
nand U9218 (N_9218,N_8273,N_8319);
or U9219 (N_9219,N_8493,N_8983);
and U9220 (N_9220,N_8594,N_8336);
nand U9221 (N_9221,N_8010,N_8011);
nor U9222 (N_9222,N_8636,N_8221);
nand U9223 (N_9223,N_8046,N_8797);
nor U9224 (N_9224,N_8304,N_8198);
and U9225 (N_9225,N_8637,N_8544);
or U9226 (N_9226,N_8760,N_8826);
nor U9227 (N_9227,N_8951,N_8012);
nor U9228 (N_9228,N_8701,N_8793);
nand U9229 (N_9229,N_8610,N_8989);
nor U9230 (N_9230,N_8517,N_8039);
nand U9231 (N_9231,N_8383,N_8556);
nand U9232 (N_9232,N_8541,N_8409);
or U9233 (N_9233,N_8220,N_8362);
nand U9234 (N_9234,N_8257,N_8737);
and U9235 (N_9235,N_8966,N_8411);
nand U9236 (N_9236,N_8004,N_8455);
or U9237 (N_9237,N_8145,N_8653);
or U9238 (N_9238,N_8085,N_8202);
nor U9239 (N_9239,N_8300,N_8894);
or U9240 (N_9240,N_8630,N_8239);
or U9241 (N_9241,N_8315,N_8483);
and U9242 (N_9242,N_8917,N_8839);
or U9243 (N_9243,N_8558,N_8063);
nand U9244 (N_9244,N_8621,N_8275);
nand U9245 (N_9245,N_8222,N_8225);
nand U9246 (N_9246,N_8549,N_8402);
and U9247 (N_9247,N_8321,N_8702);
nor U9248 (N_9248,N_8811,N_8952);
nor U9249 (N_9249,N_8704,N_8901);
nor U9250 (N_9250,N_8855,N_8591);
nand U9251 (N_9251,N_8248,N_8696);
nand U9252 (N_9252,N_8242,N_8570);
and U9253 (N_9253,N_8117,N_8334);
and U9254 (N_9254,N_8494,N_8137);
nand U9255 (N_9255,N_8557,N_8710);
xor U9256 (N_9256,N_8525,N_8850);
or U9257 (N_9257,N_8465,N_8552);
nor U9258 (N_9258,N_8246,N_8197);
and U9259 (N_9259,N_8134,N_8357);
or U9260 (N_9260,N_8296,N_8530);
and U9261 (N_9261,N_8783,N_8993);
or U9262 (N_9262,N_8690,N_8187);
nand U9263 (N_9263,N_8538,N_8733);
nand U9264 (N_9264,N_8295,N_8581);
nand U9265 (N_9265,N_8876,N_8511);
and U9266 (N_9266,N_8022,N_8753);
and U9267 (N_9267,N_8323,N_8613);
or U9268 (N_9268,N_8813,N_8567);
and U9269 (N_9269,N_8886,N_8371);
and U9270 (N_9270,N_8472,N_8507);
or U9271 (N_9271,N_8434,N_8734);
nor U9272 (N_9272,N_8049,N_8566);
nand U9273 (N_9273,N_8649,N_8648);
nand U9274 (N_9274,N_8976,N_8482);
nor U9275 (N_9275,N_8087,N_8968);
nand U9276 (N_9276,N_8339,N_8475);
or U9277 (N_9277,N_8037,N_8578);
xnor U9278 (N_9278,N_8188,N_8595);
nand U9279 (N_9279,N_8219,N_8463);
and U9280 (N_9280,N_8763,N_8231);
and U9281 (N_9281,N_8757,N_8289);
nand U9282 (N_9282,N_8674,N_8115);
and U9283 (N_9283,N_8018,N_8668);
or U9284 (N_9284,N_8445,N_8848);
or U9285 (N_9285,N_8924,N_8670);
or U9286 (N_9286,N_8102,N_8822);
and U9287 (N_9287,N_8982,N_8588);
nand U9288 (N_9288,N_8641,N_8707);
and U9289 (N_9289,N_8105,N_8044);
nor U9290 (N_9290,N_8965,N_8429);
nand U9291 (N_9291,N_8192,N_8163);
nand U9292 (N_9292,N_8051,N_8437);
nand U9293 (N_9293,N_8852,N_8036);
or U9294 (N_9294,N_8353,N_8571);
nand U9295 (N_9295,N_8778,N_8938);
nand U9296 (N_9296,N_8640,N_8727);
and U9297 (N_9297,N_8664,N_8256);
nand U9298 (N_9298,N_8700,N_8164);
or U9299 (N_9299,N_8928,N_8060);
and U9300 (N_9300,N_8528,N_8794);
or U9301 (N_9301,N_8804,N_8108);
nor U9302 (N_9302,N_8861,N_8157);
and U9303 (N_9303,N_8332,N_8798);
nand U9304 (N_9304,N_8430,N_8962);
nor U9305 (N_9305,N_8614,N_8678);
or U9306 (N_9306,N_8652,N_8229);
nor U9307 (N_9307,N_8258,N_8781);
or U9308 (N_9308,N_8750,N_8279);
nand U9309 (N_9309,N_8159,N_8773);
nor U9310 (N_9310,N_8672,N_8714);
or U9311 (N_9311,N_8040,N_8599);
or U9312 (N_9312,N_8490,N_8885);
and U9313 (N_9313,N_8837,N_8041);
nor U9314 (N_9314,N_8864,N_8466);
nor U9315 (N_9315,N_8892,N_8593);
and U9316 (N_9316,N_8226,N_8825);
and U9317 (N_9317,N_8884,N_8205);
nand U9318 (N_9318,N_8243,N_8381);
nor U9319 (N_9319,N_8019,N_8123);
nor U9320 (N_9320,N_8114,N_8992);
nor U9321 (N_9321,N_8746,N_8329);
or U9322 (N_9322,N_8912,N_8185);
or U9323 (N_9323,N_8732,N_8898);
or U9324 (N_9324,N_8140,N_8873);
or U9325 (N_9325,N_8435,N_8452);
and U9326 (N_9326,N_8712,N_8268);
and U9327 (N_9327,N_8891,N_8305);
nor U9328 (N_9328,N_8251,N_8691);
nand U9329 (N_9329,N_8872,N_8464);
nand U9330 (N_9330,N_8629,N_8130);
nor U9331 (N_9331,N_8206,N_8388);
nand U9332 (N_9332,N_8679,N_8500);
and U9333 (N_9333,N_8651,N_8697);
or U9334 (N_9334,N_8632,N_8741);
nand U9335 (N_9335,N_8713,N_8240);
nand U9336 (N_9336,N_8853,N_8352);
nand U9337 (N_9337,N_8364,N_8831);
and U9338 (N_9338,N_8680,N_8442);
nand U9339 (N_9339,N_8887,N_8382);
nor U9340 (N_9340,N_8906,N_8934);
xor U9341 (N_9341,N_8542,N_8874);
nor U9342 (N_9342,N_8523,N_8390);
nand U9343 (N_9343,N_8973,N_8245);
nand U9344 (N_9344,N_8503,N_8143);
nor U9345 (N_9345,N_8462,N_8953);
or U9346 (N_9346,N_8625,N_8112);
or U9347 (N_9347,N_8881,N_8167);
or U9348 (N_9348,N_8550,N_8408);
nand U9349 (N_9349,N_8270,N_8646);
or U9350 (N_9350,N_8618,N_8375);
and U9351 (N_9351,N_8423,N_8502);
nor U9352 (N_9352,N_8380,N_8116);
nor U9353 (N_9353,N_8828,N_8392);
nand U9354 (N_9354,N_8858,N_8911);
nand U9355 (N_9355,N_8418,N_8478);
or U9356 (N_9356,N_8878,N_8729);
nor U9357 (N_9357,N_8302,N_8271);
nor U9358 (N_9358,N_8250,N_8189);
nor U9359 (N_9359,N_8035,N_8988);
nand U9360 (N_9360,N_8775,N_8555);
and U9361 (N_9361,N_8919,N_8195);
nor U9362 (N_9362,N_8438,N_8572);
nor U9363 (N_9363,N_8908,N_8054);
or U9364 (N_9364,N_8237,N_8236);
nor U9365 (N_9365,N_8405,N_8807);
or U9366 (N_9366,N_8693,N_8643);
or U9367 (N_9367,N_8436,N_8842);
nor U9368 (N_9368,N_8914,N_8711);
nand U9369 (N_9369,N_8367,N_8433);
and U9370 (N_9370,N_8565,N_8526);
nand U9371 (N_9371,N_8344,N_8692);
and U9372 (N_9372,N_8480,N_8761);
or U9373 (N_9373,N_8521,N_8916);
xnor U9374 (N_9374,N_8642,N_8453);
nand U9375 (N_9375,N_8792,N_8086);
nor U9376 (N_9376,N_8260,N_8389);
or U9377 (N_9377,N_8788,N_8253);
nor U9378 (N_9378,N_8799,N_8447);
and U9379 (N_9379,N_8829,N_8481);
and U9380 (N_9380,N_8871,N_8348);
nand U9381 (N_9381,N_8959,N_8065);
xnor U9382 (N_9382,N_8154,N_8573);
nor U9383 (N_9383,N_8634,N_8385);
nand U9384 (N_9384,N_8654,N_8133);
and U9385 (N_9385,N_8394,N_8851);
xor U9386 (N_9386,N_8399,N_8488);
nand U9387 (N_9387,N_8605,N_8456);
or U9388 (N_9388,N_8166,N_8095);
nand U9389 (N_9389,N_8925,N_8754);
and U9390 (N_9390,N_8173,N_8944);
nand U9391 (N_9391,N_8926,N_8061);
nand U9392 (N_9392,N_8534,N_8358);
nand U9393 (N_9393,N_8417,N_8512);
nor U9394 (N_9394,N_8119,N_8290);
nand U9395 (N_9395,N_8328,N_8006);
or U9396 (N_9396,N_8101,N_8177);
and U9397 (N_9397,N_8728,N_8374);
and U9398 (N_9398,N_8963,N_8361);
or U9399 (N_9399,N_8814,N_8935);
nor U9400 (N_9400,N_8171,N_8498);
and U9401 (N_9401,N_8787,N_8306);
nor U9402 (N_9402,N_8883,N_8078);
nor U9403 (N_9403,N_8428,N_8539);
nor U9404 (N_9404,N_8509,N_8937);
or U9405 (N_9405,N_8003,N_8032);
nor U9406 (N_9406,N_8131,N_8823);
and U9407 (N_9407,N_8808,N_8208);
and U9408 (N_9408,N_8128,N_8499);
or U9409 (N_9409,N_8583,N_8597);
or U9410 (N_9410,N_8738,N_8819);
nor U9411 (N_9411,N_8147,N_8536);
and U9412 (N_9412,N_8596,N_8608);
nand U9413 (N_9413,N_8942,N_8110);
and U9414 (N_9414,N_8818,N_8169);
nand U9415 (N_9415,N_8719,N_8888);
and U9416 (N_9416,N_8709,N_8739);
or U9417 (N_9417,N_8327,N_8077);
nand U9418 (N_9418,N_8686,N_8895);
and U9419 (N_9419,N_8785,N_8458);
nand U9420 (N_9420,N_8695,N_8830);
nand U9421 (N_9421,N_8922,N_8790);
or U9422 (N_9422,N_8070,N_8160);
and U9423 (N_9423,N_8745,N_8068);
nand U9424 (N_9424,N_8722,N_8181);
nand U9425 (N_9425,N_8999,N_8506);
or U9426 (N_9426,N_8803,N_8252);
and U9427 (N_9427,N_8638,N_8705);
nand U9428 (N_9428,N_8161,N_8184);
and U9429 (N_9429,N_8031,N_8286);
xnor U9430 (N_9430,N_8235,N_8228);
and U9431 (N_9431,N_8207,N_8223);
or U9432 (N_9432,N_8153,N_8230);
and U9433 (N_9433,N_8024,N_8373);
xnor U9434 (N_9434,N_8416,N_8414);
nor U9435 (N_9435,N_8647,N_8407);
and U9436 (N_9436,N_8964,N_8340);
or U9437 (N_9437,N_8008,N_8540);
and U9438 (N_9438,N_8639,N_8349);
nor U9439 (N_9439,N_8687,N_8866);
and U9440 (N_9440,N_8190,N_8461);
nor U9441 (N_9441,N_8843,N_8468);
and U9442 (N_9442,N_8211,N_8023);
and U9443 (N_9443,N_8563,N_8090);
or U9444 (N_9444,N_8398,N_8121);
and U9445 (N_9445,N_8940,N_8846);
and U9446 (N_9446,N_8657,N_8152);
nand U9447 (N_9447,N_8644,N_8915);
and U9448 (N_9448,N_8645,N_8533);
and U9449 (N_9449,N_8324,N_8857);
or U9450 (N_9450,N_8673,N_8404);
nor U9451 (N_9451,N_8685,N_8448);
or U9452 (N_9452,N_8397,N_8969);
and U9453 (N_9453,N_8860,N_8111);
or U9454 (N_9454,N_8569,N_8609);
nor U9455 (N_9455,N_8377,N_8849);
or U9456 (N_9456,N_8425,N_8816);
and U9457 (N_9457,N_8615,N_8960);
nor U9458 (N_9458,N_8217,N_8351);
or U9459 (N_9459,N_8833,N_8805);
or U9460 (N_9460,N_8441,N_8562);
and U9461 (N_9461,N_8820,N_8360);
or U9462 (N_9462,N_8342,N_8847);
and U9463 (N_9463,N_8859,N_8655);
nor U9464 (N_9464,N_8261,N_8838);
or U9465 (N_9465,N_8387,N_8904);
nor U9466 (N_9466,N_8183,N_8264);
or U9467 (N_9467,N_8725,N_8470);
nor U9468 (N_9468,N_8139,N_8439);
or U9469 (N_9469,N_8449,N_8132);
or U9470 (N_9470,N_8477,N_8093);
and U9471 (N_9471,N_8548,N_8724);
nor U9472 (N_9472,N_8048,N_8619);
nand U9473 (N_9473,N_8033,N_8473);
nor U9474 (N_9474,N_8522,N_8755);
nor U9475 (N_9475,N_8554,N_8956);
or U9476 (N_9476,N_8990,N_8038);
nand U9477 (N_9477,N_8393,N_8355);
nand U9478 (N_9478,N_8731,N_8097);
nor U9479 (N_9479,N_8267,N_8958);
or U9480 (N_9480,N_8081,N_8865);
or U9481 (N_9481,N_8505,N_8665);
xnor U9482 (N_9482,N_8880,N_8923);
nand U9483 (N_9483,N_8084,N_8689);
nor U9484 (N_9484,N_8627,N_8124);
or U9485 (N_9485,N_8772,N_8307);
nor U9486 (N_9486,N_8354,N_8186);
or U9487 (N_9487,N_8016,N_8972);
and U9488 (N_9488,N_8450,N_8350);
nand U9489 (N_9489,N_8401,N_8088);
and U9490 (N_9490,N_8426,N_8650);
nor U9491 (N_9491,N_8486,N_8546);
or U9492 (N_9492,N_8671,N_8170);
or U9493 (N_9493,N_8059,N_8182);
and U9494 (N_9494,N_8715,N_8987);
nand U9495 (N_9495,N_8768,N_8069);
and U9496 (N_9496,N_8683,N_8484);
nand U9497 (N_9497,N_8995,N_8291);
or U9498 (N_9498,N_8287,N_8603);
and U9499 (N_9499,N_8313,N_8014);
or U9500 (N_9500,N_8491,N_8390);
nor U9501 (N_9501,N_8666,N_8172);
or U9502 (N_9502,N_8984,N_8294);
nand U9503 (N_9503,N_8899,N_8516);
nor U9504 (N_9504,N_8517,N_8556);
or U9505 (N_9505,N_8299,N_8467);
nor U9506 (N_9506,N_8216,N_8214);
or U9507 (N_9507,N_8042,N_8554);
nor U9508 (N_9508,N_8525,N_8513);
or U9509 (N_9509,N_8108,N_8042);
nor U9510 (N_9510,N_8289,N_8764);
and U9511 (N_9511,N_8263,N_8715);
nor U9512 (N_9512,N_8793,N_8607);
or U9513 (N_9513,N_8295,N_8480);
nand U9514 (N_9514,N_8531,N_8213);
nor U9515 (N_9515,N_8536,N_8806);
and U9516 (N_9516,N_8621,N_8510);
xnor U9517 (N_9517,N_8404,N_8629);
nand U9518 (N_9518,N_8078,N_8340);
nor U9519 (N_9519,N_8689,N_8377);
and U9520 (N_9520,N_8126,N_8911);
or U9521 (N_9521,N_8906,N_8859);
and U9522 (N_9522,N_8248,N_8311);
and U9523 (N_9523,N_8346,N_8641);
or U9524 (N_9524,N_8553,N_8231);
and U9525 (N_9525,N_8408,N_8489);
or U9526 (N_9526,N_8421,N_8971);
or U9527 (N_9527,N_8456,N_8369);
and U9528 (N_9528,N_8865,N_8896);
or U9529 (N_9529,N_8898,N_8344);
nor U9530 (N_9530,N_8635,N_8562);
nand U9531 (N_9531,N_8392,N_8490);
nand U9532 (N_9532,N_8811,N_8998);
or U9533 (N_9533,N_8631,N_8385);
and U9534 (N_9534,N_8598,N_8654);
and U9535 (N_9535,N_8338,N_8250);
or U9536 (N_9536,N_8327,N_8046);
and U9537 (N_9537,N_8240,N_8743);
nor U9538 (N_9538,N_8526,N_8825);
xnor U9539 (N_9539,N_8833,N_8494);
and U9540 (N_9540,N_8578,N_8339);
and U9541 (N_9541,N_8578,N_8770);
or U9542 (N_9542,N_8646,N_8714);
or U9543 (N_9543,N_8428,N_8888);
nand U9544 (N_9544,N_8086,N_8005);
and U9545 (N_9545,N_8697,N_8926);
nor U9546 (N_9546,N_8882,N_8709);
nor U9547 (N_9547,N_8803,N_8048);
nand U9548 (N_9548,N_8913,N_8444);
nor U9549 (N_9549,N_8473,N_8713);
nor U9550 (N_9550,N_8752,N_8566);
or U9551 (N_9551,N_8477,N_8677);
nand U9552 (N_9552,N_8035,N_8768);
nand U9553 (N_9553,N_8154,N_8593);
nor U9554 (N_9554,N_8065,N_8994);
nand U9555 (N_9555,N_8341,N_8973);
nand U9556 (N_9556,N_8785,N_8339);
nor U9557 (N_9557,N_8427,N_8131);
and U9558 (N_9558,N_8876,N_8100);
and U9559 (N_9559,N_8972,N_8362);
or U9560 (N_9560,N_8839,N_8265);
nand U9561 (N_9561,N_8567,N_8182);
and U9562 (N_9562,N_8545,N_8654);
or U9563 (N_9563,N_8489,N_8277);
and U9564 (N_9564,N_8998,N_8253);
nand U9565 (N_9565,N_8729,N_8988);
nor U9566 (N_9566,N_8819,N_8995);
or U9567 (N_9567,N_8465,N_8252);
nor U9568 (N_9568,N_8849,N_8511);
or U9569 (N_9569,N_8337,N_8575);
or U9570 (N_9570,N_8596,N_8778);
nor U9571 (N_9571,N_8736,N_8459);
xnor U9572 (N_9572,N_8268,N_8481);
or U9573 (N_9573,N_8159,N_8550);
nand U9574 (N_9574,N_8252,N_8060);
nand U9575 (N_9575,N_8570,N_8013);
nor U9576 (N_9576,N_8929,N_8884);
nand U9577 (N_9577,N_8714,N_8871);
nand U9578 (N_9578,N_8675,N_8071);
nand U9579 (N_9579,N_8881,N_8939);
nor U9580 (N_9580,N_8446,N_8524);
nand U9581 (N_9581,N_8118,N_8390);
nand U9582 (N_9582,N_8539,N_8691);
and U9583 (N_9583,N_8401,N_8775);
nor U9584 (N_9584,N_8147,N_8445);
or U9585 (N_9585,N_8095,N_8860);
or U9586 (N_9586,N_8018,N_8354);
nor U9587 (N_9587,N_8737,N_8371);
nand U9588 (N_9588,N_8095,N_8460);
nand U9589 (N_9589,N_8367,N_8679);
xor U9590 (N_9590,N_8449,N_8481);
or U9591 (N_9591,N_8411,N_8315);
nand U9592 (N_9592,N_8871,N_8058);
or U9593 (N_9593,N_8021,N_8976);
nand U9594 (N_9594,N_8653,N_8593);
or U9595 (N_9595,N_8425,N_8983);
and U9596 (N_9596,N_8628,N_8422);
and U9597 (N_9597,N_8515,N_8055);
nor U9598 (N_9598,N_8015,N_8072);
nor U9599 (N_9599,N_8680,N_8609);
or U9600 (N_9600,N_8982,N_8399);
nand U9601 (N_9601,N_8601,N_8253);
or U9602 (N_9602,N_8788,N_8249);
or U9603 (N_9603,N_8989,N_8392);
and U9604 (N_9604,N_8960,N_8675);
nand U9605 (N_9605,N_8310,N_8379);
nand U9606 (N_9606,N_8280,N_8817);
nor U9607 (N_9607,N_8380,N_8514);
and U9608 (N_9608,N_8682,N_8243);
nor U9609 (N_9609,N_8285,N_8084);
and U9610 (N_9610,N_8752,N_8386);
nor U9611 (N_9611,N_8734,N_8627);
and U9612 (N_9612,N_8084,N_8258);
or U9613 (N_9613,N_8976,N_8454);
or U9614 (N_9614,N_8663,N_8311);
nand U9615 (N_9615,N_8957,N_8313);
or U9616 (N_9616,N_8201,N_8080);
and U9617 (N_9617,N_8063,N_8746);
nor U9618 (N_9618,N_8341,N_8750);
and U9619 (N_9619,N_8383,N_8618);
nor U9620 (N_9620,N_8682,N_8490);
nand U9621 (N_9621,N_8184,N_8206);
xnor U9622 (N_9622,N_8735,N_8987);
nand U9623 (N_9623,N_8477,N_8733);
nor U9624 (N_9624,N_8289,N_8160);
xnor U9625 (N_9625,N_8015,N_8166);
and U9626 (N_9626,N_8140,N_8095);
or U9627 (N_9627,N_8079,N_8211);
nor U9628 (N_9628,N_8044,N_8797);
or U9629 (N_9629,N_8847,N_8605);
nand U9630 (N_9630,N_8653,N_8014);
or U9631 (N_9631,N_8453,N_8746);
nand U9632 (N_9632,N_8087,N_8181);
nor U9633 (N_9633,N_8281,N_8413);
nor U9634 (N_9634,N_8147,N_8175);
nor U9635 (N_9635,N_8326,N_8433);
or U9636 (N_9636,N_8556,N_8829);
or U9637 (N_9637,N_8440,N_8304);
and U9638 (N_9638,N_8361,N_8505);
nor U9639 (N_9639,N_8406,N_8760);
or U9640 (N_9640,N_8573,N_8394);
and U9641 (N_9641,N_8278,N_8468);
and U9642 (N_9642,N_8450,N_8224);
nor U9643 (N_9643,N_8993,N_8297);
and U9644 (N_9644,N_8701,N_8794);
or U9645 (N_9645,N_8061,N_8811);
or U9646 (N_9646,N_8839,N_8901);
nand U9647 (N_9647,N_8502,N_8951);
nand U9648 (N_9648,N_8538,N_8800);
nand U9649 (N_9649,N_8646,N_8349);
or U9650 (N_9650,N_8180,N_8321);
nor U9651 (N_9651,N_8349,N_8144);
nand U9652 (N_9652,N_8519,N_8957);
nand U9653 (N_9653,N_8215,N_8500);
or U9654 (N_9654,N_8321,N_8219);
nand U9655 (N_9655,N_8847,N_8222);
nand U9656 (N_9656,N_8828,N_8614);
nor U9657 (N_9657,N_8499,N_8083);
or U9658 (N_9658,N_8104,N_8449);
or U9659 (N_9659,N_8082,N_8875);
and U9660 (N_9660,N_8162,N_8974);
or U9661 (N_9661,N_8539,N_8997);
nand U9662 (N_9662,N_8372,N_8929);
or U9663 (N_9663,N_8217,N_8653);
or U9664 (N_9664,N_8423,N_8289);
nand U9665 (N_9665,N_8174,N_8611);
and U9666 (N_9666,N_8884,N_8475);
and U9667 (N_9667,N_8740,N_8592);
nand U9668 (N_9668,N_8345,N_8880);
and U9669 (N_9669,N_8889,N_8286);
nand U9670 (N_9670,N_8917,N_8122);
or U9671 (N_9671,N_8664,N_8091);
and U9672 (N_9672,N_8813,N_8217);
nor U9673 (N_9673,N_8474,N_8825);
nand U9674 (N_9674,N_8628,N_8021);
nand U9675 (N_9675,N_8191,N_8036);
and U9676 (N_9676,N_8032,N_8237);
nand U9677 (N_9677,N_8031,N_8498);
and U9678 (N_9678,N_8867,N_8122);
nand U9679 (N_9679,N_8874,N_8402);
nand U9680 (N_9680,N_8864,N_8483);
nand U9681 (N_9681,N_8220,N_8908);
and U9682 (N_9682,N_8165,N_8389);
and U9683 (N_9683,N_8027,N_8675);
nor U9684 (N_9684,N_8889,N_8978);
nor U9685 (N_9685,N_8512,N_8939);
xnor U9686 (N_9686,N_8759,N_8884);
nor U9687 (N_9687,N_8220,N_8212);
nor U9688 (N_9688,N_8199,N_8264);
nand U9689 (N_9689,N_8080,N_8603);
and U9690 (N_9690,N_8513,N_8296);
nand U9691 (N_9691,N_8547,N_8154);
or U9692 (N_9692,N_8019,N_8993);
or U9693 (N_9693,N_8204,N_8017);
and U9694 (N_9694,N_8711,N_8776);
or U9695 (N_9695,N_8730,N_8717);
or U9696 (N_9696,N_8324,N_8802);
or U9697 (N_9697,N_8531,N_8073);
or U9698 (N_9698,N_8817,N_8690);
or U9699 (N_9699,N_8429,N_8376);
and U9700 (N_9700,N_8607,N_8458);
or U9701 (N_9701,N_8889,N_8452);
nand U9702 (N_9702,N_8879,N_8313);
or U9703 (N_9703,N_8785,N_8797);
or U9704 (N_9704,N_8642,N_8354);
or U9705 (N_9705,N_8033,N_8303);
nand U9706 (N_9706,N_8934,N_8083);
and U9707 (N_9707,N_8138,N_8069);
and U9708 (N_9708,N_8599,N_8939);
or U9709 (N_9709,N_8176,N_8662);
nand U9710 (N_9710,N_8328,N_8122);
and U9711 (N_9711,N_8052,N_8807);
nand U9712 (N_9712,N_8366,N_8211);
nand U9713 (N_9713,N_8251,N_8511);
or U9714 (N_9714,N_8542,N_8254);
and U9715 (N_9715,N_8027,N_8437);
and U9716 (N_9716,N_8765,N_8885);
or U9717 (N_9717,N_8448,N_8793);
nand U9718 (N_9718,N_8010,N_8248);
nand U9719 (N_9719,N_8333,N_8058);
nand U9720 (N_9720,N_8884,N_8127);
nor U9721 (N_9721,N_8566,N_8879);
and U9722 (N_9722,N_8349,N_8103);
and U9723 (N_9723,N_8300,N_8673);
nand U9724 (N_9724,N_8453,N_8823);
nor U9725 (N_9725,N_8851,N_8305);
or U9726 (N_9726,N_8783,N_8913);
nand U9727 (N_9727,N_8461,N_8974);
or U9728 (N_9728,N_8600,N_8155);
and U9729 (N_9729,N_8938,N_8253);
nand U9730 (N_9730,N_8802,N_8023);
and U9731 (N_9731,N_8555,N_8783);
nand U9732 (N_9732,N_8994,N_8479);
xor U9733 (N_9733,N_8204,N_8004);
nand U9734 (N_9734,N_8563,N_8793);
nor U9735 (N_9735,N_8434,N_8586);
or U9736 (N_9736,N_8590,N_8730);
nor U9737 (N_9737,N_8842,N_8201);
nand U9738 (N_9738,N_8324,N_8835);
nor U9739 (N_9739,N_8531,N_8360);
and U9740 (N_9740,N_8970,N_8247);
and U9741 (N_9741,N_8735,N_8915);
nor U9742 (N_9742,N_8949,N_8918);
and U9743 (N_9743,N_8302,N_8137);
and U9744 (N_9744,N_8209,N_8092);
nor U9745 (N_9745,N_8041,N_8944);
nor U9746 (N_9746,N_8356,N_8295);
nand U9747 (N_9747,N_8735,N_8382);
or U9748 (N_9748,N_8603,N_8441);
or U9749 (N_9749,N_8254,N_8061);
nand U9750 (N_9750,N_8139,N_8002);
and U9751 (N_9751,N_8969,N_8633);
and U9752 (N_9752,N_8888,N_8174);
and U9753 (N_9753,N_8521,N_8717);
or U9754 (N_9754,N_8702,N_8977);
xor U9755 (N_9755,N_8507,N_8512);
nor U9756 (N_9756,N_8899,N_8954);
and U9757 (N_9757,N_8666,N_8543);
or U9758 (N_9758,N_8050,N_8835);
and U9759 (N_9759,N_8349,N_8621);
nor U9760 (N_9760,N_8314,N_8614);
nor U9761 (N_9761,N_8641,N_8644);
or U9762 (N_9762,N_8893,N_8304);
nor U9763 (N_9763,N_8695,N_8329);
or U9764 (N_9764,N_8893,N_8185);
nand U9765 (N_9765,N_8911,N_8176);
and U9766 (N_9766,N_8019,N_8953);
nor U9767 (N_9767,N_8980,N_8061);
or U9768 (N_9768,N_8211,N_8914);
nand U9769 (N_9769,N_8623,N_8995);
nand U9770 (N_9770,N_8148,N_8490);
or U9771 (N_9771,N_8715,N_8228);
nand U9772 (N_9772,N_8050,N_8448);
nor U9773 (N_9773,N_8583,N_8829);
nor U9774 (N_9774,N_8545,N_8279);
and U9775 (N_9775,N_8816,N_8493);
and U9776 (N_9776,N_8526,N_8193);
nor U9777 (N_9777,N_8108,N_8316);
nand U9778 (N_9778,N_8569,N_8874);
nand U9779 (N_9779,N_8483,N_8149);
xor U9780 (N_9780,N_8918,N_8441);
or U9781 (N_9781,N_8450,N_8278);
nand U9782 (N_9782,N_8890,N_8416);
nor U9783 (N_9783,N_8286,N_8694);
and U9784 (N_9784,N_8927,N_8333);
and U9785 (N_9785,N_8480,N_8433);
or U9786 (N_9786,N_8245,N_8938);
or U9787 (N_9787,N_8905,N_8288);
and U9788 (N_9788,N_8163,N_8062);
or U9789 (N_9789,N_8079,N_8863);
or U9790 (N_9790,N_8007,N_8415);
nand U9791 (N_9791,N_8323,N_8281);
and U9792 (N_9792,N_8240,N_8925);
nand U9793 (N_9793,N_8454,N_8499);
or U9794 (N_9794,N_8819,N_8946);
xor U9795 (N_9795,N_8519,N_8222);
and U9796 (N_9796,N_8683,N_8537);
or U9797 (N_9797,N_8597,N_8029);
and U9798 (N_9798,N_8303,N_8756);
and U9799 (N_9799,N_8516,N_8986);
nand U9800 (N_9800,N_8308,N_8911);
and U9801 (N_9801,N_8353,N_8975);
nor U9802 (N_9802,N_8270,N_8043);
and U9803 (N_9803,N_8318,N_8334);
nand U9804 (N_9804,N_8641,N_8828);
nor U9805 (N_9805,N_8262,N_8291);
nor U9806 (N_9806,N_8487,N_8029);
and U9807 (N_9807,N_8866,N_8167);
nor U9808 (N_9808,N_8862,N_8436);
xor U9809 (N_9809,N_8435,N_8173);
nor U9810 (N_9810,N_8335,N_8905);
nand U9811 (N_9811,N_8472,N_8992);
nor U9812 (N_9812,N_8870,N_8539);
nor U9813 (N_9813,N_8978,N_8072);
or U9814 (N_9814,N_8338,N_8746);
nor U9815 (N_9815,N_8614,N_8397);
nand U9816 (N_9816,N_8305,N_8848);
or U9817 (N_9817,N_8128,N_8869);
nand U9818 (N_9818,N_8681,N_8161);
or U9819 (N_9819,N_8107,N_8872);
nand U9820 (N_9820,N_8910,N_8152);
or U9821 (N_9821,N_8153,N_8688);
nand U9822 (N_9822,N_8436,N_8096);
nand U9823 (N_9823,N_8393,N_8331);
nand U9824 (N_9824,N_8574,N_8014);
nor U9825 (N_9825,N_8494,N_8560);
and U9826 (N_9826,N_8292,N_8172);
nand U9827 (N_9827,N_8549,N_8242);
nand U9828 (N_9828,N_8591,N_8602);
nor U9829 (N_9829,N_8034,N_8963);
and U9830 (N_9830,N_8992,N_8634);
and U9831 (N_9831,N_8848,N_8891);
nor U9832 (N_9832,N_8781,N_8717);
or U9833 (N_9833,N_8141,N_8688);
or U9834 (N_9834,N_8017,N_8447);
nor U9835 (N_9835,N_8502,N_8975);
xnor U9836 (N_9836,N_8832,N_8302);
and U9837 (N_9837,N_8355,N_8418);
nand U9838 (N_9838,N_8823,N_8612);
and U9839 (N_9839,N_8860,N_8979);
or U9840 (N_9840,N_8728,N_8838);
or U9841 (N_9841,N_8510,N_8674);
xnor U9842 (N_9842,N_8726,N_8824);
or U9843 (N_9843,N_8061,N_8493);
and U9844 (N_9844,N_8214,N_8884);
nand U9845 (N_9845,N_8241,N_8322);
or U9846 (N_9846,N_8657,N_8981);
nand U9847 (N_9847,N_8169,N_8608);
nor U9848 (N_9848,N_8149,N_8907);
or U9849 (N_9849,N_8274,N_8371);
nor U9850 (N_9850,N_8264,N_8978);
nor U9851 (N_9851,N_8565,N_8825);
and U9852 (N_9852,N_8051,N_8497);
and U9853 (N_9853,N_8539,N_8259);
nor U9854 (N_9854,N_8070,N_8655);
nand U9855 (N_9855,N_8125,N_8453);
and U9856 (N_9856,N_8828,N_8627);
nand U9857 (N_9857,N_8420,N_8776);
and U9858 (N_9858,N_8792,N_8015);
xnor U9859 (N_9859,N_8794,N_8535);
nor U9860 (N_9860,N_8376,N_8227);
and U9861 (N_9861,N_8085,N_8702);
or U9862 (N_9862,N_8072,N_8262);
and U9863 (N_9863,N_8462,N_8968);
or U9864 (N_9864,N_8334,N_8289);
nand U9865 (N_9865,N_8264,N_8195);
nand U9866 (N_9866,N_8427,N_8809);
nand U9867 (N_9867,N_8996,N_8650);
and U9868 (N_9868,N_8899,N_8267);
or U9869 (N_9869,N_8198,N_8525);
or U9870 (N_9870,N_8760,N_8041);
and U9871 (N_9871,N_8670,N_8463);
and U9872 (N_9872,N_8291,N_8740);
and U9873 (N_9873,N_8679,N_8732);
nor U9874 (N_9874,N_8104,N_8358);
xor U9875 (N_9875,N_8694,N_8905);
nand U9876 (N_9876,N_8702,N_8653);
and U9877 (N_9877,N_8194,N_8871);
nor U9878 (N_9878,N_8211,N_8605);
nand U9879 (N_9879,N_8365,N_8459);
nand U9880 (N_9880,N_8605,N_8224);
or U9881 (N_9881,N_8152,N_8832);
xor U9882 (N_9882,N_8903,N_8649);
nor U9883 (N_9883,N_8313,N_8054);
xor U9884 (N_9884,N_8192,N_8930);
and U9885 (N_9885,N_8509,N_8719);
nand U9886 (N_9886,N_8608,N_8315);
or U9887 (N_9887,N_8131,N_8263);
nand U9888 (N_9888,N_8521,N_8228);
nand U9889 (N_9889,N_8541,N_8813);
and U9890 (N_9890,N_8476,N_8316);
nand U9891 (N_9891,N_8035,N_8922);
nor U9892 (N_9892,N_8776,N_8297);
or U9893 (N_9893,N_8797,N_8321);
nand U9894 (N_9894,N_8410,N_8320);
xor U9895 (N_9895,N_8980,N_8226);
nor U9896 (N_9896,N_8852,N_8524);
nand U9897 (N_9897,N_8809,N_8972);
and U9898 (N_9898,N_8976,N_8453);
and U9899 (N_9899,N_8584,N_8617);
nand U9900 (N_9900,N_8191,N_8442);
nand U9901 (N_9901,N_8765,N_8381);
and U9902 (N_9902,N_8765,N_8718);
nand U9903 (N_9903,N_8010,N_8988);
nand U9904 (N_9904,N_8034,N_8359);
nor U9905 (N_9905,N_8995,N_8800);
and U9906 (N_9906,N_8435,N_8084);
or U9907 (N_9907,N_8908,N_8045);
and U9908 (N_9908,N_8691,N_8833);
nand U9909 (N_9909,N_8136,N_8790);
or U9910 (N_9910,N_8806,N_8332);
nor U9911 (N_9911,N_8606,N_8583);
nand U9912 (N_9912,N_8339,N_8993);
nor U9913 (N_9913,N_8642,N_8062);
xnor U9914 (N_9914,N_8104,N_8540);
and U9915 (N_9915,N_8861,N_8614);
nor U9916 (N_9916,N_8259,N_8235);
or U9917 (N_9917,N_8715,N_8719);
nand U9918 (N_9918,N_8759,N_8951);
nor U9919 (N_9919,N_8010,N_8243);
nor U9920 (N_9920,N_8853,N_8894);
nand U9921 (N_9921,N_8023,N_8596);
nand U9922 (N_9922,N_8686,N_8731);
and U9923 (N_9923,N_8878,N_8466);
nand U9924 (N_9924,N_8604,N_8200);
or U9925 (N_9925,N_8702,N_8194);
or U9926 (N_9926,N_8634,N_8485);
and U9927 (N_9927,N_8307,N_8047);
nor U9928 (N_9928,N_8776,N_8972);
or U9929 (N_9929,N_8201,N_8260);
nor U9930 (N_9930,N_8860,N_8152);
nor U9931 (N_9931,N_8910,N_8387);
nor U9932 (N_9932,N_8200,N_8765);
nand U9933 (N_9933,N_8083,N_8190);
nand U9934 (N_9934,N_8995,N_8507);
and U9935 (N_9935,N_8956,N_8068);
nand U9936 (N_9936,N_8536,N_8153);
nor U9937 (N_9937,N_8368,N_8559);
and U9938 (N_9938,N_8130,N_8742);
or U9939 (N_9939,N_8308,N_8580);
or U9940 (N_9940,N_8842,N_8185);
and U9941 (N_9941,N_8696,N_8040);
nand U9942 (N_9942,N_8800,N_8798);
nand U9943 (N_9943,N_8182,N_8560);
and U9944 (N_9944,N_8469,N_8944);
nor U9945 (N_9945,N_8043,N_8042);
nand U9946 (N_9946,N_8814,N_8536);
or U9947 (N_9947,N_8446,N_8292);
or U9948 (N_9948,N_8061,N_8429);
and U9949 (N_9949,N_8583,N_8132);
nand U9950 (N_9950,N_8226,N_8057);
nand U9951 (N_9951,N_8988,N_8891);
or U9952 (N_9952,N_8023,N_8765);
nor U9953 (N_9953,N_8997,N_8598);
nand U9954 (N_9954,N_8714,N_8372);
nand U9955 (N_9955,N_8970,N_8400);
nor U9956 (N_9956,N_8935,N_8596);
and U9957 (N_9957,N_8164,N_8123);
and U9958 (N_9958,N_8147,N_8816);
nor U9959 (N_9959,N_8347,N_8171);
and U9960 (N_9960,N_8561,N_8828);
nor U9961 (N_9961,N_8481,N_8904);
and U9962 (N_9962,N_8605,N_8196);
or U9963 (N_9963,N_8047,N_8414);
or U9964 (N_9964,N_8858,N_8522);
or U9965 (N_9965,N_8716,N_8775);
or U9966 (N_9966,N_8167,N_8619);
nor U9967 (N_9967,N_8944,N_8952);
and U9968 (N_9968,N_8710,N_8554);
nand U9969 (N_9969,N_8853,N_8699);
or U9970 (N_9970,N_8969,N_8764);
nor U9971 (N_9971,N_8019,N_8190);
nor U9972 (N_9972,N_8097,N_8027);
and U9973 (N_9973,N_8387,N_8364);
and U9974 (N_9974,N_8457,N_8662);
and U9975 (N_9975,N_8254,N_8223);
or U9976 (N_9976,N_8236,N_8465);
or U9977 (N_9977,N_8511,N_8621);
nor U9978 (N_9978,N_8075,N_8475);
nand U9979 (N_9979,N_8509,N_8152);
nor U9980 (N_9980,N_8289,N_8664);
nor U9981 (N_9981,N_8475,N_8114);
or U9982 (N_9982,N_8513,N_8459);
nand U9983 (N_9983,N_8672,N_8937);
nor U9984 (N_9984,N_8212,N_8160);
and U9985 (N_9985,N_8890,N_8230);
and U9986 (N_9986,N_8822,N_8706);
or U9987 (N_9987,N_8521,N_8206);
nand U9988 (N_9988,N_8216,N_8441);
nor U9989 (N_9989,N_8043,N_8414);
and U9990 (N_9990,N_8000,N_8869);
nand U9991 (N_9991,N_8612,N_8787);
nand U9992 (N_9992,N_8221,N_8050);
nor U9993 (N_9993,N_8849,N_8137);
nor U9994 (N_9994,N_8131,N_8400);
nor U9995 (N_9995,N_8894,N_8339);
nand U9996 (N_9996,N_8693,N_8867);
and U9997 (N_9997,N_8374,N_8722);
nor U9998 (N_9998,N_8287,N_8799);
or U9999 (N_9999,N_8287,N_8777);
nand UO_0 (O_0,N_9859,N_9230);
or UO_1 (O_1,N_9048,N_9463);
nor UO_2 (O_2,N_9383,N_9284);
or UO_3 (O_3,N_9897,N_9535);
or UO_4 (O_4,N_9370,N_9121);
and UO_5 (O_5,N_9307,N_9496);
nor UO_6 (O_6,N_9014,N_9367);
and UO_7 (O_7,N_9570,N_9471);
or UO_8 (O_8,N_9693,N_9511);
nor UO_9 (O_9,N_9842,N_9641);
or UO_10 (O_10,N_9628,N_9372);
nand UO_11 (O_11,N_9928,N_9276);
nor UO_12 (O_12,N_9402,N_9504);
or UO_13 (O_13,N_9821,N_9484);
or UO_14 (O_14,N_9246,N_9186);
nor UO_15 (O_15,N_9938,N_9262);
and UO_16 (O_16,N_9459,N_9659);
or UO_17 (O_17,N_9783,N_9063);
nand UO_18 (O_18,N_9019,N_9267);
or UO_19 (O_19,N_9323,N_9984);
nor UO_20 (O_20,N_9639,N_9272);
nor UO_21 (O_21,N_9066,N_9444);
or UO_22 (O_22,N_9492,N_9971);
or UO_23 (O_23,N_9243,N_9024);
nor UO_24 (O_24,N_9830,N_9960);
and UO_25 (O_25,N_9438,N_9612);
and UO_26 (O_26,N_9348,N_9603);
or UO_27 (O_27,N_9039,N_9390);
or UO_28 (O_28,N_9685,N_9103);
xnor UO_29 (O_29,N_9137,N_9180);
nand UO_30 (O_30,N_9819,N_9923);
nor UO_31 (O_31,N_9599,N_9654);
nor UO_32 (O_32,N_9555,N_9507);
nand UO_33 (O_33,N_9715,N_9489);
nand UO_34 (O_34,N_9510,N_9907);
nor UO_35 (O_35,N_9857,N_9688);
nor UO_36 (O_36,N_9605,N_9889);
or UO_37 (O_37,N_9018,N_9170);
or UO_38 (O_38,N_9881,N_9860);
and UO_39 (O_39,N_9914,N_9544);
nor UO_40 (O_40,N_9041,N_9601);
xor UO_41 (O_41,N_9754,N_9271);
and UO_42 (O_42,N_9891,N_9211);
or UO_43 (O_43,N_9523,N_9855);
or UO_44 (O_44,N_9179,N_9485);
nor UO_45 (O_45,N_9849,N_9532);
or UO_46 (O_46,N_9616,N_9545);
nand UO_47 (O_47,N_9123,N_9106);
or UO_48 (O_48,N_9579,N_9957);
or UO_49 (O_49,N_9032,N_9518);
or UO_50 (O_50,N_9756,N_9665);
or UO_51 (O_51,N_9345,N_9217);
nor UO_52 (O_52,N_9576,N_9714);
nor UO_53 (O_53,N_9131,N_9983);
and UO_54 (O_54,N_9711,N_9038);
xor UO_55 (O_55,N_9139,N_9076);
or UO_56 (O_56,N_9514,N_9158);
and UO_57 (O_57,N_9780,N_9409);
nand UO_58 (O_58,N_9350,N_9245);
and UO_59 (O_59,N_9361,N_9051);
and UO_60 (O_60,N_9346,N_9846);
nand UO_61 (O_61,N_9719,N_9644);
xnor UO_62 (O_62,N_9304,N_9992);
and UO_63 (O_63,N_9253,N_9446);
or UO_64 (O_64,N_9672,N_9297);
and UO_65 (O_65,N_9132,N_9887);
nor UO_66 (O_66,N_9396,N_9606);
and UO_67 (O_67,N_9499,N_9764);
and UO_68 (O_68,N_9280,N_9306);
nor UO_69 (O_69,N_9582,N_9286);
or UO_70 (O_70,N_9493,N_9737);
nor UO_71 (O_71,N_9573,N_9153);
or UO_72 (O_72,N_9801,N_9144);
nand UO_73 (O_73,N_9427,N_9125);
and UO_74 (O_74,N_9317,N_9423);
and UO_75 (O_75,N_9909,N_9739);
or UO_76 (O_76,N_9084,N_9724);
or UO_77 (O_77,N_9017,N_9788);
or UO_78 (O_78,N_9160,N_9115);
or UO_79 (O_79,N_9791,N_9939);
nand UO_80 (O_80,N_9474,N_9070);
nand UO_81 (O_81,N_9255,N_9242);
nor UO_82 (O_82,N_9666,N_9344);
xnor UO_83 (O_83,N_9389,N_9833);
nor UO_84 (O_84,N_9210,N_9425);
or UO_85 (O_85,N_9716,N_9634);
or UO_86 (O_86,N_9454,N_9572);
nor UO_87 (O_87,N_9260,N_9723);
and UO_88 (O_88,N_9373,N_9966);
nor UO_89 (O_89,N_9352,N_9977);
xnor UO_90 (O_90,N_9093,N_9657);
nor UO_91 (O_91,N_9642,N_9406);
and UO_92 (O_92,N_9325,N_9809);
and UO_93 (O_93,N_9053,N_9356);
xnor UO_94 (O_94,N_9495,N_9234);
and UO_95 (O_95,N_9192,N_9730);
nor UO_96 (O_96,N_9519,N_9185);
or UO_97 (O_97,N_9633,N_9640);
or UO_98 (O_98,N_9962,N_9274);
nor UO_99 (O_99,N_9073,N_9589);
or UO_100 (O_100,N_9237,N_9945);
and UO_101 (O_101,N_9117,N_9422);
nor UO_102 (O_102,N_9216,N_9003);
and UO_103 (O_103,N_9335,N_9910);
and UO_104 (O_104,N_9786,N_9974);
and UO_105 (O_105,N_9126,N_9130);
or UO_106 (O_106,N_9200,N_9787);
or UO_107 (O_107,N_9840,N_9915);
nor UO_108 (O_108,N_9675,N_9162);
nand UO_109 (O_109,N_9655,N_9741);
nand UO_110 (O_110,N_9080,N_9177);
nand UO_111 (O_111,N_9903,N_9885);
nand UO_112 (O_112,N_9205,N_9526);
nand UO_113 (O_113,N_9434,N_9414);
nor UO_114 (O_114,N_9638,N_9671);
or UO_115 (O_115,N_9785,N_9790);
nand UO_116 (O_116,N_9827,N_9305);
and UO_117 (O_117,N_9293,N_9105);
or UO_118 (O_118,N_9109,N_9797);
and UO_119 (O_119,N_9173,N_9701);
or UO_120 (O_120,N_9021,N_9033);
and UO_121 (O_121,N_9759,N_9450);
nor UO_122 (O_122,N_9602,N_9278);
or UO_123 (O_123,N_9238,N_9298);
and UO_124 (O_124,N_9773,N_9886);
nand UO_125 (O_125,N_9733,N_9340);
or UO_126 (O_126,N_9023,N_9997);
or UO_127 (O_127,N_9037,N_9865);
nand UO_128 (O_128,N_9294,N_9405);
or UO_129 (O_129,N_9623,N_9822);
or UO_130 (O_130,N_9586,N_9175);
nor UO_131 (O_131,N_9696,N_9538);
nor UO_132 (O_132,N_9189,N_9228);
or UO_133 (O_133,N_9761,N_9445);
and UO_134 (O_134,N_9236,N_9858);
or UO_135 (O_135,N_9001,N_9101);
nor UO_136 (O_136,N_9895,N_9890);
or UO_137 (O_137,N_9751,N_9300);
nor UO_138 (O_138,N_9497,N_9154);
or UO_139 (O_139,N_9964,N_9631);
nand UO_140 (O_140,N_9922,N_9433);
and UO_141 (O_141,N_9698,N_9618);
nand UO_142 (O_142,N_9480,N_9810);
nor UO_143 (O_143,N_9678,N_9637);
nor UO_144 (O_144,N_9784,N_9184);
and UO_145 (O_145,N_9240,N_9250);
nand UO_146 (O_146,N_9580,N_9836);
and UO_147 (O_147,N_9443,N_9584);
nor UO_148 (O_148,N_9826,N_9967);
nand UO_149 (O_149,N_9442,N_9432);
nand UO_150 (O_150,N_9371,N_9904);
nor UO_151 (O_151,N_9662,N_9789);
or UO_152 (O_152,N_9202,N_9762);
nor UO_153 (O_153,N_9068,N_9525);
or UO_154 (O_154,N_9439,N_9086);
or UO_155 (O_155,N_9987,N_9428);
nor UO_156 (O_156,N_9447,N_9862);
and UO_157 (O_157,N_9851,N_9481);
nor UO_158 (O_158,N_9159,N_9869);
nand UO_159 (O_159,N_9385,N_9407);
nor UO_160 (O_160,N_9941,N_9506);
nor UO_161 (O_161,N_9558,N_9416);
or UO_162 (O_162,N_9172,N_9218);
nand UO_163 (O_163,N_9204,N_9883);
or UO_164 (O_164,N_9649,N_9387);
or UO_165 (O_165,N_9408,N_9709);
and UO_166 (O_166,N_9501,N_9148);
nor UO_167 (O_167,N_9430,N_9911);
or UO_168 (O_168,N_9248,N_9308);
or UO_169 (O_169,N_9046,N_9136);
or UO_170 (O_170,N_9884,N_9338);
and UO_171 (O_171,N_9798,N_9195);
nand UO_172 (O_172,N_9985,N_9295);
nor UO_173 (O_173,N_9866,N_9410);
and UO_174 (O_174,N_9333,N_9825);
or UO_175 (O_175,N_9533,N_9163);
and UO_176 (O_176,N_9000,N_9479);
and UO_177 (O_177,N_9948,N_9959);
nor UO_178 (O_178,N_9670,N_9712);
nor UO_179 (O_179,N_9134,N_9973);
and UO_180 (O_180,N_9475,N_9635);
or UO_181 (O_181,N_9074,N_9800);
nor UO_182 (O_182,N_9301,N_9980);
or UO_183 (O_183,N_9806,N_9913);
nand UO_184 (O_184,N_9691,N_9164);
nand UO_185 (O_185,N_9465,N_9950);
or UO_186 (O_186,N_9375,N_9477);
and UO_187 (O_187,N_9363,N_9660);
nand UO_188 (O_188,N_9156,N_9873);
and UO_189 (O_189,N_9081,N_9264);
or UO_190 (O_190,N_9088,N_9231);
nor UO_191 (O_191,N_9779,N_9169);
nor UO_192 (O_192,N_9401,N_9469);
nor UO_193 (O_193,N_9415,N_9607);
and UO_194 (O_194,N_9133,N_9976);
nor UO_195 (O_195,N_9285,N_9462);
or UO_196 (O_196,N_9986,N_9050);
nand UO_197 (O_197,N_9832,N_9355);
and UO_198 (O_198,N_9288,N_9774);
or UO_199 (O_199,N_9811,N_9968);
and UO_200 (O_200,N_9958,N_9850);
and UO_201 (O_201,N_9608,N_9328);
nand UO_202 (O_202,N_9878,N_9956);
nor UO_203 (O_203,N_9540,N_9682);
nor UO_204 (O_204,N_9040,N_9494);
or UO_205 (O_205,N_9282,N_9488);
nand UO_206 (O_206,N_9543,N_9632);
or UO_207 (O_207,N_9515,N_9888);
nand UO_208 (O_208,N_9279,N_9744);
nor UO_209 (O_209,N_9951,N_9690);
and UO_210 (O_210,N_9145,N_9007);
or UO_211 (O_211,N_9818,N_9176);
and UO_212 (O_212,N_9763,N_9843);
or UO_213 (O_213,N_9578,N_9547);
and UO_214 (O_214,N_9694,N_9542);
or UO_215 (O_215,N_9585,N_9440);
xnor UO_216 (O_216,N_9012,N_9235);
nand UO_217 (O_217,N_9567,N_9222);
or UO_218 (O_218,N_9880,N_9223);
or UO_219 (O_219,N_9766,N_9362);
and UO_220 (O_220,N_9557,N_9057);
nor UO_221 (O_221,N_9667,N_9291);
or UO_222 (O_222,N_9174,N_9892);
nand UO_223 (O_223,N_9005,N_9347);
nor UO_224 (O_224,N_9726,N_9368);
nor UO_225 (O_225,N_9208,N_9996);
or UO_226 (O_226,N_9326,N_9646);
nand UO_227 (O_227,N_9182,N_9729);
xor UO_228 (O_228,N_9482,N_9491);
nor UO_229 (O_229,N_9342,N_9932);
nand UO_230 (O_230,N_9838,N_9868);
nor UO_231 (O_231,N_9203,N_9871);
or UO_232 (O_232,N_9457,N_9815);
and UO_233 (O_233,N_9877,N_9487);
nor UO_234 (O_234,N_9949,N_9593);
and UO_235 (O_235,N_9676,N_9364);
nor UO_236 (O_236,N_9187,N_9856);
nand UO_237 (O_237,N_9717,N_9772);
nand UO_238 (O_238,N_9844,N_9219);
or UO_239 (O_239,N_9142,N_9935);
nor UO_240 (O_240,N_9527,N_9466);
or UO_241 (O_241,N_9513,N_9596);
nand UO_242 (O_242,N_9327,N_9930);
and UO_243 (O_243,N_9379,N_9359);
or UO_244 (O_244,N_9583,N_9963);
nor UO_245 (O_245,N_9096,N_9400);
and UO_246 (O_246,N_9102,N_9829);
or UO_247 (O_247,N_9703,N_9831);
nor UO_248 (O_248,N_9556,N_9686);
and UO_249 (O_249,N_9100,N_9718);
or UO_250 (O_250,N_9118,N_9942);
nand UO_251 (O_251,N_9995,N_9934);
nand UO_252 (O_252,N_9736,N_9095);
xor UO_253 (O_253,N_9214,N_9768);
or UO_254 (O_254,N_9498,N_9706);
or UO_255 (O_255,N_9357,N_9025);
or UO_256 (O_256,N_9517,N_9413);
or UO_257 (O_257,N_9529,N_9568);
nor UO_258 (O_258,N_9734,N_9699);
xnor UO_259 (O_259,N_9165,N_9059);
nor UO_260 (O_260,N_9331,N_9653);
and UO_261 (O_261,N_9728,N_9664);
or UO_262 (O_262,N_9738,N_9429);
nor UO_263 (O_263,N_9652,N_9448);
nand UO_264 (O_264,N_9929,N_9975);
nand UO_265 (O_265,N_9199,N_9550);
nand UO_266 (O_266,N_9104,N_9044);
and UO_267 (O_267,N_9943,N_9979);
or UO_268 (O_268,N_9075,N_9912);
nor UO_269 (O_269,N_9626,N_9876);
nand UO_270 (O_270,N_9680,N_9027);
nand UO_271 (O_271,N_9595,N_9029);
xnor UO_272 (O_272,N_9224,N_9324);
nand UO_273 (O_273,N_9417,N_9872);
nand UO_274 (O_274,N_9321,N_9770);
nand UO_275 (O_275,N_9534,N_9269);
or UO_276 (O_276,N_9455,N_9263);
and UO_277 (O_277,N_9178,N_9314);
xor UO_278 (O_278,N_9157,N_9955);
or UO_279 (O_279,N_9839,N_9099);
and UO_280 (O_280,N_9055,N_9658);
and UO_281 (O_281,N_9735,N_9266);
nand UO_282 (O_282,N_9502,N_9970);
and UO_283 (O_283,N_9918,N_9648);
nand UO_284 (O_284,N_9509,N_9311);
nor UO_285 (O_285,N_9569,N_9536);
nand UO_286 (O_286,N_9380,N_9581);
nor UO_287 (O_287,N_9135,N_9114);
and UO_288 (O_288,N_9707,N_9229);
nor UO_289 (O_289,N_9225,N_9767);
xnor UO_290 (O_290,N_9852,N_9150);
nor UO_291 (O_291,N_9061,N_9643);
nor UO_292 (O_292,N_9587,N_9171);
and UO_293 (O_293,N_9702,N_9194);
nor UO_294 (O_294,N_9537,N_9470);
nand UO_295 (O_295,N_9988,N_9745);
nor UO_296 (O_296,N_9814,N_9151);
or UO_297 (O_297,N_9619,N_9874);
nand UO_298 (O_298,N_9393,N_9054);
and UO_299 (O_299,N_9590,N_9899);
nand UO_300 (O_300,N_9392,N_9908);
nand UO_301 (O_301,N_9065,N_9813);
or UO_302 (O_302,N_9207,N_9879);
nor UO_303 (O_303,N_9853,N_9281);
xnor UO_304 (O_304,N_9742,N_9931);
nand UO_305 (O_305,N_9900,N_9620);
xnor UO_306 (O_306,N_9622,N_9574);
nand UO_307 (O_307,N_9817,N_9467);
and UO_308 (O_308,N_9064,N_9528);
and UO_309 (O_309,N_9270,N_9399);
or UO_310 (O_310,N_9588,N_9917);
nand UO_311 (O_311,N_9720,N_9337);
nand UO_312 (O_312,N_9140,N_9863);
nand UO_313 (O_313,N_9905,N_9369);
nor UO_314 (O_314,N_9265,N_9722);
or UO_315 (O_315,N_9227,N_9010);
nor UO_316 (O_316,N_9206,N_9760);
xor UO_317 (O_317,N_9365,N_9743);
and UO_318 (O_318,N_9559,N_9894);
or UO_319 (O_319,N_9629,N_9336);
nor UO_320 (O_320,N_9087,N_9116);
nor UO_321 (O_321,N_9149,N_9841);
or UO_322 (O_322,N_9188,N_9615);
nand UO_323 (O_323,N_9875,N_9847);
nor UO_324 (O_324,N_9468,N_9167);
nand UO_325 (O_325,N_9777,N_9113);
xor UO_326 (O_326,N_9677,N_9656);
and UO_327 (O_327,N_9600,N_9028);
xor UO_328 (O_328,N_9940,N_9530);
or UO_329 (O_329,N_9577,N_9244);
and UO_330 (O_330,N_9056,N_9072);
or UO_331 (O_331,N_9143,N_9757);
nor UO_332 (O_332,N_9112,N_9473);
or UO_333 (O_333,N_9315,N_9110);
nor UO_334 (O_334,N_9820,N_9034);
nor UO_335 (O_335,N_9564,N_9896);
nor UO_336 (O_336,N_9845,N_9681);
nand UO_337 (O_337,N_9376,N_9412);
nand UO_338 (O_338,N_9394,N_9343);
nor UO_339 (O_339,N_9740,N_9009);
or UO_340 (O_340,N_9503,N_9299);
and UO_341 (O_341,N_9047,N_9122);
nand UO_342 (O_342,N_9378,N_9598);
and UO_343 (O_343,N_9239,N_9226);
xor UO_344 (O_344,N_9531,N_9097);
and UO_345 (O_345,N_9478,N_9727);
or UO_346 (O_346,N_9614,N_9036);
and UO_347 (O_347,N_9837,N_9998);
nand UO_348 (O_348,N_9098,N_9661);
nand UO_349 (O_349,N_9566,N_9289);
nor UO_350 (O_350,N_9043,N_9085);
nand UO_351 (O_351,N_9746,N_9391);
nor UO_352 (O_352,N_9561,N_9927);
nor UO_353 (O_353,N_9312,N_9209);
and UO_354 (O_354,N_9627,N_9549);
nor UO_355 (O_355,N_9403,N_9259);
nand UO_356 (O_356,N_9092,N_9329);
nor UO_357 (O_357,N_9546,N_9953);
or UO_358 (O_358,N_9360,N_9252);
and UO_359 (O_359,N_9898,N_9591);
nand UO_360 (O_360,N_9453,N_9094);
and UO_361 (O_361,N_9381,N_9674);
or UO_362 (O_362,N_9476,N_9944);
nor UO_363 (O_363,N_9554,N_9552);
nand UO_364 (O_364,N_9366,N_9058);
and UO_365 (O_365,N_9981,N_9794);
nor UO_366 (O_366,N_9524,N_9647);
or UO_367 (O_367,N_9421,N_9435);
and UO_368 (O_368,N_9650,N_9349);
or UO_369 (O_369,N_9700,N_9141);
nand UO_370 (O_370,N_9775,N_9418);
or UO_371 (O_371,N_9936,N_9330);
nor UO_372 (O_372,N_9273,N_9309);
nor UO_373 (O_373,N_9750,N_9748);
and UO_374 (O_374,N_9420,N_9120);
nand UO_375 (O_375,N_9002,N_9351);
nand UO_376 (O_376,N_9937,N_9213);
nor UO_377 (O_377,N_9395,N_9864);
or UO_378 (O_378,N_9926,N_9424);
and UO_379 (O_379,N_9198,N_9256);
and UO_380 (O_380,N_9919,N_9322);
or UO_381 (O_381,N_9008,N_9991);
nand UO_382 (O_382,N_9969,N_9548);
nand UO_383 (O_383,N_9013,N_9020);
or UO_384 (O_384,N_9316,N_9212);
and UO_385 (O_385,N_9334,N_9804);
and UO_386 (O_386,N_9030,N_9332);
nor UO_387 (O_387,N_9521,N_9999);
nand UO_388 (O_388,N_9490,N_9769);
or UO_389 (O_389,N_9341,N_9695);
and UO_390 (O_390,N_9386,N_9310);
or UO_391 (O_391,N_9834,N_9906);
nand UO_392 (O_392,N_9052,N_9778);
nand UO_393 (O_393,N_9138,N_9249);
or UO_394 (O_394,N_9689,N_9077);
nand UO_395 (O_395,N_9196,N_9796);
or UO_396 (O_396,N_9426,N_9456);
nand UO_397 (O_397,N_9708,N_9035);
nor UO_398 (O_398,N_9609,N_9848);
nand UO_399 (O_399,N_9683,N_9684);
or UO_400 (O_400,N_9181,N_9083);
nand UO_401 (O_401,N_9129,N_9516);
nand UO_402 (O_402,N_9079,N_9802);
and UO_403 (O_403,N_9500,N_9725);
or UO_404 (O_404,N_9215,N_9128);
nand UO_405 (O_405,N_9374,N_9464);
nand UO_406 (O_406,N_9107,N_9233);
nor UO_407 (O_407,N_9303,N_9042);
and UO_408 (O_408,N_9867,N_9771);
nand UO_409 (O_409,N_9776,N_9431);
and UO_410 (O_410,N_9449,N_9460);
nand UO_411 (O_411,N_9965,N_9902);
nor UO_412 (O_412,N_9071,N_9006);
nor UO_413 (O_413,N_9508,N_9982);
or UO_414 (O_414,N_9015,N_9563);
or UO_415 (O_415,N_9067,N_9713);
and UO_416 (O_416,N_9803,N_9697);
xnor UO_417 (O_417,N_9283,N_9512);
and UO_418 (O_418,N_9078,N_9625);
nand UO_419 (O_419,N_9782,N_9292);
nor UO_420 (O_420,N_9990,N_9382);
or UO_421 (O_421,N_9011,N_9320);
and UO_422 (O_422,N_9404,N_9946);
xor UO_423 (O_423,N_9108,N_9947);
or UO_424 (O_424,N_9565,N_9630);
and UO_425 (O_425,N_9539,N_9069);
xnor UO_426 (O_426,N_9679,N_9755);
and UO_427 (O_427,N_9155,N_9916);
nor UO_428 (O_428,N_9663,N_9854);
or UO_429 (O_429,N_9287,N_9978);
or UO_430 (O_430,N_9925,N_9994);
xor UO_431 (O_431,N_9232,N_9765);
or UO_432 (O_432,N_9835,N_9621);
nor UO_433 (O_433,N_9520,N_9472);
and UO_434 (O_434,N_9193,N_9045);
or UO_435 (O_435,N_9617,N_9452);
and UO_436 (O_436,N_9793,N_9870);
and UO_437 (O_437,N_9220,N_9636);
or UO_438 (O_438,N_9749,N_9384);
and UO_439 (O_439,N_9575,N_9592);
nor UO_440 (O_440,N_9277,N_9247);
nor UO_441 (O_441,N_9687,N_9183);
or UO_442 (O_442,N_9339,N_9673);
nand UO_443 (O_443,N_9313,N_9275);
and UO_444 (O_444,N_9828,N_9026);
or UO_445 (O_445,N_9824,N_9799);
nor UO_446 (O_446,N_9060,N_9319);
and UO_447 (O_447,N_9451,N_9721);
or UO_448 (O_448,N_9091,N_9704);
nand UO_449 (O_449,N_9354,N_9016);
nand UO_450 (O_450,N_9611,N_9146);
nand UO_451 (O_451,N_9597,N_9221);
nor UO_452 (O_452,N_9388,N_9419);
nor UO_453 (O_453,N_9124,N_9082);
or UO_454 (O_454,N_9111,N_9004);
or UO_455 (O_455,N_9358,N_9254);
nor UO_456 (O_456,N_9377,N_9645);
nor UO_457 (O_457,N_9522,N_9553);
or UO_458 (O_458,N_9753,N_9732);
nor UO_459 (O_459,N_9747,N_9901);
nand UO_460 (O_460,N_9920,N_9437);
and UO_461 (O_461,N_9483,N_9551);
nor UO_462 (O_462,N_9152,N_9961);
nand UO_463 (O_463,N_9090,N_9692);
and UO_464 (O_464,N_9807,N_9812);
nor UO_465 (O_465,N_9921,N_9651);
and UO_466 (O_466,N_9168,N_9486);
nor UO_467 (O_467,N_9808,N_9290);
or UO_468 (O_468,N_9166,N_9792);
nor UO_469 (O_469,N_9710,N_9823);
nand UO_470 (O_470,N_9604,N_9258);
nor UO_471 (O_471,N_9261,N_9562);
nand UO_472 (O_472,N_9397,N_9560);
nor UO_473 (O_473,N_9398,N_9624);
nand UO_474 (O_474,N_9952,N_9571);
or UO_475 (O_475,N_9731,N_9147);
nor UO_476 (O_476,N_9805,N_9594);
nor UO_477 (O_477,N_9861,N_9241);
nand UO_478 (O_478,N_9924,N_9954);
nand UO_479 (O_479,N_9461,N_9752);
xor UO_480 (O_480,N_9296,N_9972);
nor UO_481 (O_481,N_9089,N_9893);
and UO_482 (O_482,N_9302,N_9318);
xnor UO_483 (O_483,N_9882,N_9062);
nor UO_484 (O_484,N_9161,N_9441);
or UO_485 (O_485,N_9758,N_9197);
nor UO_486 (O_486,N_9668,N_9031);
or UO_487 (O_487,N_9049,N_9816);
nand UO_488 (O_488,N_9795,N_9268);
and UO_489 (O_489,N_9933,N_9781);
and UO_490 (O_490,N_9705,N_9190);
or UO_491 (O_491,N_9127,N_9613);
nand UO_492 (O_492,N_9022,N_9505);
or UO_493 (O_493,N_9989,N_9610);
nor UO_494 (O_494,N_9436,N_9993);
or UO_495 (O_495,N_9191,N_9411);
or UO_496 (O_496,N_9669,N_9458);
or UO_497 (O_497,N_9353,N_9201);
nand UO_498 (O_498,N_9541,N_9257);
nor UO_499 (O_499,N_9251,N_9119);
nand UO_500 (O_500,N_9977,N_9584);
nor UO_501 (O_501,N_9732,N_9027);
or UO_502 (O_502,N_9251,N_9455);
nor UO_503 (O_503,N_9197,N_9612);
and UO_504 (O_504,N_9750,N_9414);
nand UO_505 (O_505,N_9837,N_9514);
or UO_506 (O_506,N_9125,N_9137);
nor UO_507 (O_507,N_9655,N_9830);
nor UO_508 (O_508,N_9420,N_9134);
xor UO_509 (O_509,N_9411,N_9527);
and UO_510 (O_510,N_9723,N_9746);
and UO_511 (O_511,N_9358,N_9044);
xnor UO_512 (O_512,N_9946,N_9367);
and UO_513 (O_513,N_9958,N_9288);
and UO_514 (O_514,N_9551,N_9158);
or UO_515 (O_515,N_9247,N_9485);
nand UO_516 (O_516,N_9853,N_9623);
nand UO_517 (O_517,N_9589,N_9517);
nand UO_518 (O_518,N_9800,N_9540);
or UO_519 (O_519,N_9832,N_9688);
or UO_520 (O_520,N_9243,N_9836);
nor UO_521 (O_521,N_9083,N_9797);
and UO_522 (O_522,N_9402,N_9973);
nor UO_523 (O_523,N_9187,N_9507);
or UO_524 (O_524,N_9243,N_9878);
or UO_525 (O_525,N_9509,N_9998);
and UO_526 (O_526,N_9148,N_9412);
nor UO_527 (O_527,N_9392,N_9299);
nor UO_528 (O_528,N_9630,N_9437);
or UO_529 (O_529,N_9328,N_9758);
nor UO_530 (O_530,N_9200,N_9106);
nor UO_531 (O_531,N_9629,N_9165);
nand UO_532 (O_532,N_9062,N_9506);
xor UO_533 (O_533,N_9232,N_9333);
nand UO_534 (O_534,N_9575,N_9691);
and UO_535 (O_535,N_9782,N_9743);
and UO_536 (O_536,N_9219,N_9330);
and UO_537 (O_537,N_9197,N_9429);
nand UO_538 (O_538,N_9208,N_9115);
or UO_539 (O_539,N_9063,N_9767);
nor UO_540 (O_540,N_9827,N_9360);
nand UO_541 (O_541,N_9878,N_9014);
and UO_542 (O_542,N_9387,N_9733);
nor UO_543 (O_543,N_9934,N_9515);
and UO_544 (O_544,N_9541,N_9514);
nor UO_545 (O_545,N_9033,N_9592);
nor UO_546 (O_546,N_9789,N_9443);
or UO_547 (O_547,N_9894,N_9977);
or UO_548 (O_548,N_9192,N_9150);
and UO_549 (O_549,N_9620,N_9481);
and UO_550 (O_550,N_9913,N_9406);
nor UO_551 (O_551,N_9859,N_9342);
or UO_552 (O_552,N_9504,N_9621);
xnor UO_553 (O_553,N_9011,N_9978);
and UO_554 (O_554,N_9179,N_9166);
or UO_555 (O_555,N_9781,N_9853);
nand UO_556 (O_556,N_9206,N_9355);
or UO_557 (O_557,N_9279,N_9383);
nand UO_558 (O_558,N_9769,N_9208);
nand UO_559 (O_559,N_9236,N_9165);
and UO_560 (O_560,N_9755,N_9292);
nor UO_561 (O_561,N_9102,N_9506);
and UO_562 (O_562,N_9266,N_9167);
or UO_563 (O_563,N_9459,N_9277);
nor UO_564 (O_564,N_9958,N_9289);
nor UO_565 (O_565,N_9920,N_9537);
or UO_566 (O_566,N_9020,N_9457);
nor UO_567 (O_567,N_9892,N_9743);
xnor UO_568 (O_568,N_9517,N_9677);
and UO_569 (O_569,N_9978,N_9968);
nand UO_570 (O_570,N_9303,N_9168);
and UO_571 (O_571,N_9997,N_9183);
or UO_572 (O_572,N_9303,N_9858);
or UO_573 (O_573,N_9780,N_9943);
nand UO_574 (O_574,N_9211,N_9066);
nor UO_575 (O_575,N_9501,N_9525);
nor UO_576 (O_576,N_9080,N_9133);
nor UO_577 (O_577,N_9660,N_9681);
nand UO_578 (O_578,N_9761,N_9379);
nand UO_579 (O_579,N_9991,N_9394);
nand UO_580 (O_580,N_9532,N_9083);
nor UO_581 (O_581,N_9191,N_9622);
and UO_582 (O_582,N_9689,N_9885);
nand UO_583 (O_583,N_9938,N_9494);
nand UO_584 (O_584,N_9974,N_9709);
or UO_585 (O_585,N_9298,N_9131);
or UO_586 (O_586,N_9882,N_9535);
or UO_587 (O_587,N_9368,N_9231);
nand UO_588 (O_588,N_9365,N_9294);
and UO_589 (O_589,N_9248,N_9442);
and UO_590 (O_590,N_9645,N_9230);
and UO_591 (O_591,N_9078,N_9167);
nor UO_592 (O_592,N_9035,N_9226);
or UO_593 (O_593,N_9685,N_9797);
or UO_594 (O_594,N_9421,N_9473);
and UO_595 (O_595,N_9979,N_9827);
nor UO_596 (O_596,N_9723,N_9272);
nand UO_597 (O_597,N_9281,N_9920);
nand UO_598 (O_598,N_9848,N_9389);
nand UO_599 (O_599,N_9989,N_9237);
or UO_600 (O_600,N_9896,N_9766);
nand UO_601 (O_601,N_9374,N_9621);
and UO_602 (O_602,N_9630,N_9795);
or UO_603 (O_603,N_9210,N_9468);
nand UO_604 (O_604,N_9523,N_9844);
or UO_605 (O_605,N_9639,N_9294);
and UO_606 (O_606,N_9561,N_9462);
or UO_607 (O_607,N_9601,N_9116);
or UO_608 (O_608,N_9921,N_9313);
nor UO_609 (O_609,N_9132,N_9455);
and UO_610 (O_610,N_9042,N_9868);
nor UO_611 (O_611,N_9957,N_9994);
and UO_612 (O_612,N_9889,N_9217);
nor UO_613 (O_613,N_9230,N_9670);
nor UO_614 (O_614,N_9218,N_9858);
xnor UO_615 (O_615,N_9111,N_9947);
or UO_616 (O_616,N_9669,N_9813);
nand UO_617 (O_617,N_9645,N_9353);
nor UO_618 (O_618,N_9183,N_9708);
or UO_619 (O_619,N_9710,N_9795);
and UO_620 (O_620,N_9495,N_9083);
nand UO_621 (O_621,N_9934,N_9944);
or UO_622 (O_622,N_9960,N_9788);
and UO_623 (O_623,N_9181,N_9978);
nand UO_624 (O_624,N_9042,N_9466);
nor UO_625 (O_625,N_9521,N_9125);
nor UO_626 (O_626,N_9019,N_9003);
nor UO_627 (O_627,N_9969,N_9739);
nor UO_628 (O_628,N_9242,N_9838);
xnor UO_629 (O_629,N_9920,N_9262);
or UO_630 (O_630,N_9721,N_9702);
or UO_631 (O_631,N_9641,N_9988);
nor UO_632 (O_632,N_9269,N_9784);
or UO_633 (O_633,N_9672,N_9463);
and UO_634 (O_634,N_9056,N_9919);
and UO_635 (O_635,N_9932,N_9297);
nand UO_636 (O_636,N_9768,N_9319);
and UO_637 (O_637,N_9450,N_9548);
nor UO_638 (O_638,N_9389,N_9746);
and UO_639 (O_639,N_9654,N_9440);
xnor UO_640 (O_640,N_9850,N_9504);
nor UO_641 (O_641,N_9286,N_9971);
or UO_642 (O_642,N_9363,N_9214);
or UO_643 (O_643,N_9406,N_9401);
nor UO_644 (O_644,N_9652,N_9259);
and UO_645 (O_645,N_9747,N_9373);
or UO_646 (O_646,N_9487,N_9452);
nor UO_647 (O_647,N_9542,N_9676);
nor UO_648 (O_648,N_9272,N_9754);
and UO_649 (O_649,N_9831,N_9096);
nand UO_650 (O_650,N_9136,N_9440);
and UO_651 (O_651,N_9181,N_9443);
nand UO_652 (O_652,N_9761,N_9044);
nand UO_653 (O_653,N_9654,N_9084);
nand UO_654 (O_654,N_9864,N_9928);
xor UO_655 (O_655,N_9836,N_9967);
nor UO_656 (O_656,N_9173,N_9497);
and UO_657 (O_657,N_9932,N_9098);
nand UO_658 (O_658,N_9632,N_9128);
nand UO_659 (O_659,N_9911,N_9079);
or UO_660 (O_660,N_9263,N_9383);
and UO_661 (O_661,N_9857,N_9778);
nor UO_662 (O_662,N_9541,N_9943);
and UO_663 (O_663,N_9273,N_9762);
and UO_664 (O_664,N_9653,N_9259);
or UO_665 (O_665,N_9783,N_9485);
nand UO_666 (O_666,N_9513,N_9986);
nor UO_667 (O_667,N_9787,N_9991);
nor UO_668 (O_668,N_9975,N_9693);
nand UO_669 (O_669,N_9868,N_9860);
or UO_670 (O_670,N_9931,N_9807);
nor UO_671 (O_671,N_9286,N_9550);
nor UO_672 (O_672,N_9756,N_9153);
xor UO_673 (O_673,N_9736,N_9469);
or UO_674 (O_674,N_9932,N_9094);
nor UO_675 (O_675,N_9252,N_9313);
and UO_676 (O_676,N_9810,N_9745);
nor UO_677 (O_677,N_9793,N_9644);
nand UO_678 (O_678,N_9573,N_9528);
nor UO_679 (O_679,N_9833,N_9254);
or UO_680 (O_680,N_9179,N_9002);
or UO_681 (O_681,N_9183,N_9587);
and UO_682 (O_682,N_9034,N_9095);
and UO_683 (O_683,N_9843,N_9346);
nor UO_684 (O_684,N_9792,N_9592);
nand UO_685 (O_685,N_9070,N_9321);
nand UO_686 (O_686,N_9522,N_9040);
nor UO_687 (O_687,N_9093,N_9277);
nor UO_688 (O_688,N_9593,N_9452);
or UO_689 (O_689,N_9596,N_9091);
and UO_690 (O_690,N_9297,N_9828);
xnor UO_691 (O_691,N_9717,N_9153);
or UO_692 (O_692,N_9714,N_9860);
and UO_693 (O_693,N_9776,N_9775);
nor UO_694 (O_694,N_9666,N_9794);
nor UO_695 (O_695,N_9869,N_9174);
and UO_696 (O_696,N_9139,N_9481);
and UO_697 (O_697,N_9549,N_9500);
or UO_698 (O_698,N_9439,N_9844);
or UO_699 (O_699,N_9828,N_9132);
or UO_700 (O_700,N_9622,N_9639);
xnor UO_701 (O_701,N_9721,N_9458);
and UO_702 (O_702,N_9408,N_9407);
or UO_703 (O_703,N_9813,N_9658);
and UO_704 (O_704,N_9223,N_9065);
and UO_705 (O_705,N_9654,N_9401);
or UO_706 (O_706,N_9270,N_9963);
nand UO_707 (O_707,N_9108,N_9021);
or UO_708 (O_708,N_9575,N_9727);
nand UO_709 (O_709,N_9551,N_9830);
nand UO_710 (O_710,N_9841,N_9163);
nand UO_711 (O_711,N_9972,N_9144);
and UO_712 (O_712,N_9830,N_9924);
nand UO_713 (O_713,N_9090,N_9626);
or UO_714 (O_714,N_9584,N_9107);
or UO_715 (O_715,N_9201,N_9690);
nand UO_716 (O_716,N_9313,N_9109);
nand UO_717 (O_717,N_9377,N_9444);
or UO_718 (O_718,N_9500,N_9327);
or UO_719 (O_719,N_9819,N_9271);
or UO_720 (O_720,N_9218,N_9803);
nand UO_721 (O_721,N_9558,N_9136);
nand UO_722 (O_722,N_9998,N_9545);
nand UO_723 (O_723,N_9450,N_9925);
nor UO_724 (O_724,N_9051,N_9601);
and UO_725 (O_725,N_9771,N_9995);
nand UO_726 (O_726,N_9768,N_9204);
and UO_727 (O_727,N_9611,N_9715);
nand UO_728 (O_728,N_9269,N_9696);
and UO_729 (O_729,N_9867,N_9144);
and UO_730 (O_730,N_9458,N_9097);
nor UO_731 (O_731,N_9921,N_9455);
or UO_732 (O_732,N_9670,N_9531);
and UO_733 (O_733,N_9009,N_9823);
nand UO_734 (O_734,N_9215,N_9873);
and UO_735 (O_735,N_9829,N_9379);
nand UO_736 (O_736,N_9654,N_9190);
nor UO_737 (O_737,N_9763,N_9182);
or UO_738 (O_738,N_9847,N_9548);
and UO_739 (O_739,N_9764,N_9724);
and UO_740 (O_740,N_9011,N_9762);
and UO_741 (O_741,N_9947,N_9073);
nor UO_742 (O_742,N_9332,N_9182);
and UO_743 (O_743,N_9374,N_9047);
xor UO_744 (O_744,N_9618,N_9179);
xnor UO_745 (O_745,N_9655,N_9086);
or UO_746 (O_746,N_9615,N_9157);
and UO_747 (O_747,N_9769,N_9547);
xnor UO_748 (O_748,N_9825,N_9092);
and UO_749 (O_749,N_9572,N_9516);
or UO_750 (O_750,N_9651,N_9778);
nor UO_751 (O_751,N_9965,N_9053);
nand UO_752 (O_752,N_9865,N_9537);
and UO_753 (O_753,N_9387,N_9157);
or UO_754 (O_754,N_9241,N_9494);
or UO_755 (O_755,N_9927,N_9063);
and UO_756 (O_756,N_9607,N_9988);
nand UO_757 (O_757,N_9004,N_9400);
or UO_758 (O_758,N_9672,N_9220);
nor UO_759 (O_759,N_9908,N_9095);
and UO_760 (O_760,N_9292,N_9990);
nor UO_761 (O_761,N_9467,N_9065);
nand UO_762 (O_762,N_9902,N_9213);
nor UO_763 (O_763,N_9440,N_9444);
or UO_764 (O_764,N_9819,N_9059);
and UO_765 (O_765,N_9031,N_9446);
nand UO_766 (O_766,N_9563,N_9185);
nor UO_767 (O_767,N_9930,N_9739);
nor UO_768 (O_768,N_9116,N_9913);
and UO_769 (O_769,N_9570,N_9523);
nand UO_770 (O_770,N_9246,N_9052);
and UO_771 (O_771,N_9329,N_9945);
nor UO_772 (O_772,N_9099,N_9662);
or UO_773 (O_773,N_9459,N_9406);
nor UO_774 (O_774,N_9318,N_9246);
xnor UO_775 (O_775,N_9183,N_9954);
nand UO_776 (O_776,N_9548,N_9758);
or UO_777 (O_777,N_9686,N_9466);
or UO_778 (O_778,N_9998,N_9602);
and UO_779 (O_779,N_9785,N_9455);
or UO_780 (O_780,N_9241,N_9513);
xnor UO_781 (O_781,N_9755,N_9843);
or UO_782 (O_782,N_9269,N_9907);
nor UO_783 (O_783,N_9162,N_9560);
nor UO_784 (O_784,N_9270,N_9838);
and UO_785 (O_785,N_9595,N_9472);
nor UO_786 (O_786,N_9184,N_9004);
or UO_787 (O_787,N_9655,N_9110);
nand UO_788 (O_788,N_9489,N_9447);
nand UO_789 (O_789,N_9216,N_9821);
nand UO_790 (O_790,N_9180,N_9716);
or UO_791 (O_791,N_9834,N_9740);
nor UO_792 (O_792,N_9793,N_9413);
nand UO_793 (O_793,N_9398,N_9322);
nand UO_794 (O_794,N_9723,N_9110);
nand UO_795 (O_795,N_9521,N_9243);
and UO_796 (O_796,N_9941,N_9298);
or UO_797 (O_797,N_9573,N_9161);
or UO_798 (O_798,N_9654,N_9443);
or UO_799 (O_799,N_9341,N_9893);
and UO_800 (O_800,N_9053,N_9299);
nor UO_801 (O_801,N_9712,N_9334);
nand UO_802 (O_802,N_9031,N_9045);
or UO_803 (O_803,N_9975,N_9776);
nand UO_804 (O_804,N_9886,N_9324);
nor UO_805 (O_805,N_9464,N_9867);
or UO_806 (O_806,N_9819,N_9262);
nand UO_807 (O_807,N_9835,N_9946);
or UO_808 (O_808,N_9006,N_9727);
and UO_809 (O_809,N_9102,N_9075);
nor UO_810 (O_810,N_9525,N_9245);
or UO_811 (O_811,N_9125,N_9478);
nand UO_812 (O_812,N_9353,N_9660);
nand UO_813 (O_813,N_9748,N_9287);
and UO_814 (O_814,N_9847,N_9940);
or UO_815 (O_815,N_9136,N_9577);
or UO_816 (O_816,N_9193,N_9888);
nor UO_817 (O_817,N_9249,N_9230);
nor UO_818 (O_818,N_9989,N_9412);
nand UO_819 (O_819,N_9168,N_9367);
nand UO_820 (O_820,N_9933,N_9389);
nand UO_821 (O_821,N_9516,N_9575);
nor UO_822 (O_822,N_9519,N_9528);
or UO_823 (O_823,N_9237,N_9861);
nand UO_824 (O_824,N_9547,N_9105);
or UO_825 (O_825,N_9400,N_9187);
nor UO_826 (O_826,N_9546,N_9645);
nand UO_827 (O_827,N_9157,N_9740);
nand UO_828 (O_828,N_9508,N_9163);
or UO_829 (O_829,N_9325,N_9691);
nor UO_830 (O_830,N_9850,N_9369);
nand UO_831 (O_831,N_9509,N_9791);
nand UO_832 (O_832,N_9440,N_9450);
nand UO_833 (O_833,N_9644,N_9134);
xor UO_834 (O_834,N_9002,N_9096);
nand UO_835 (O_835,N_9290,N_9307);
nand UO_836 (O_836,N_9551,N_9733);
or UO_837 (O_837,N_9042,N_9563);
and UO_838 (O_838,N_9368,N_9672);
and UO_839 (O_839,N_9776,N_9843);
and UO_840 (O_840,N_9777,N_9558);
nand UO_841 (O_841,N_9561,N_9807);
and UO_842 (O_842,N_9013,N_9182);
nor UO_843 (O_843,N_9293,N_9318);
xor UO_844 (O_844,N_9552,N_9370);
or UO_845 (O_845,N_9674,N_9296);
or UO_846 (O_846,N_9639,N_9543);
nand UO_847 (O_847,N_9493,N_9416);
nor UO_848 (O_848,N_9543,N_9828);
and UO_849 (O_849,N_9119,N_9978);
or UO_850 (O_850,N_9850,N_9538);
nor UO_851 (O_851,N_9601,N_9724);
or UO_852 (O_852,N_9501,N_9919);
or UO_853 (O_853,N_9316,N_9376);
nand UO_854 (O_854,N_9867,N_9548);
nand UO_855 (O_855,N_9095,N_9584);
nor UO_856 (O_856,N_9194,N_9833);
xor UO_857 (O_857,N_9689,N_9318);
or UO_858 (O_858,N_9968,N_9114);
and UO_859 (O_859,N_9552,N_9568);
or UO_860 (O_860,N_9400,N_9760);
nand UO_861 (O_861,N_9294,N_9482);
nor UO_862 (O_862,N_9493,N_9732);
nand UO_863 (O_863,N_9438,N_9148);
nor UO_864 (O_864,N_9953,N_9240);
xnor UO_865 (O_865,N_9501,N_9779);
nand UO_866 (O_866,N_9498,N_9417);
nor UO_867 (O_867,N_9075,N_9422);
nand UO_868 (O_868,N_9867,N_9177);
nand UO_869 (O_869,N_9201,N_9193);
nand UO_870 (O_870,N_9790,N_9340);
nor UO_871 (O_871,N_9233,N_9325);
or UO_872 (O_872,N_9412,N_9219);
or UO_873 (O_873,N_9547,N_9562);
nor UO_874 (O_874,N_9786,N_9494);
nand UO_875 (O_875,N_9918,N_9921);
nand UO_876 (O_876,N_9150,N_9560);
and UO_877 (O_877,N_9225,N_9388);
and UO_878 (O_878,N_9780,N_9729);
nor UO_879 (O_879,N_9869,N_9823);
and UO_880 (O_880,N_9647,N_9513);
and UO_881 (O_881,N_9828,N_9638);
nand UO_882 (O_882,N_9377,N_9681);
and UO_883 (O_883,N_9751,N_9976);
and UO_884 (O_884,N_9417,N_9660);
nand UO_885 (O_885,N_9252,N_9123);
nor UO_886 (O_886,N_9382,N_9945);
and UO_887 (O_887,N_9666,N_9480);
and UO_888 (O_888,N_9340,N_9146);
or UO_889 (O_889,N_9929,N_9273);
nand UO_890 (O_890,N_9041,N_9011);
nand UO_891 (O_891,N_9402,N_9121);
and UO_892 (O_892,N_9934,N_9505);
xor UO_893 (O_893,N_9475,N_9135);
or UO_894 (O_894,N_9921,N_9790);
nor UO_895 (O_895,N_9717,N_9413);
or UO_896 (O_896,N_9915,N_9364);
and UO_897 (O_897,N_9982,N_9421);
nor UO_898 (O_898,N_9276,N_9252);
and UO_899 (O_899,N_9803,N_9830);
nor UO_900 (O_900,N_9440,N_9631);
and UO_901 (O_901,N_9052,N_9232);
xor UO_902 (O_902,N_9692,N_9182);
nand UO_903 (O_903,N_9797,N_9188);
xnor UO_904 (O_904,N_9424,N_9427);
nand UO_905 (O_905,N_9513,N_9484);
nand UO_906 (O_906,N_9673,N_9573);
nand UO_907 (O_907,N_9720,N_9575);
or UO_908 (O_908,N_9065,N_9209);
nand UO_909 (O_909,N_9617,N_9935);
nand UO_910 (O_910,N_9506,N_9675);
xnor UO_911 (O_911,N_9680,N_9839);
nor UO_912 (O_912,N_9557,N_9822);
nor UO_913 (O_913,N_9874,N_9551);
nand UO_914 (O_914,N_9900,N_9038);
and UO_915 (O_915,N_9699,N_9380);
or UO_916 (O_916,N_9599,N_9129);
or UO_917 (O_917,N_9650,N_9369);
nand UO_918 (O_918,N_9341,N_9002);
and UO_919 (O_919,N_9334,N_9905);
nand UO_920 (O_920,N_9214,N_9220);
or UO_921 (O_921,N_9863,N_9254);
or UO_922 (O_922,N_9893,N_9054);
nor UO_923 (O_923,N_9543,N_9476);
and UO_924 (O_924,N_9384,N_9144);
nand UO_925 (O_925,N_9729,N_9232);
nand UO_926 (O_926,N_9994,N_9652);
nor UO_927 (O_927,N_9361,N_9762);
nor UO_928 (O_928,N_9230,N_9557);
or UO_929 (O_929,N_9375,N_9399);
nor UO_930 (O_930,N_9301,N_9446);
nand UO_931 (O_931,N_9493,N_9189);
or UO_932 (O_932,N_9483,N_9268);
nor UO_933 (O_933,N_9976,N_9335);
nor UO_934 (O_934,N_9513,N_9546);
nand UO_935 (O_935,N_9795,N_9539);
and UO_936 (O_936,N_9322,N_9652);
nor UO_937 (O_937,N_9651,N_9672);
or UO_938 (O_938,N_9336,N_9172);
and UO_939 (O_939,N_9615,N_9416);
nor UO_940 (O_940,N_9264,N_9338);
nand UO_941 (O_941,N_9505,N_9810);
and UO_942 (O_942,N_9109,N_9691);
nor UO_943 (O_943,N_9742,N_9248);
nand UO_944 (O_944,N_9614,N_9878);
and UO_945 (O_945,N_9356,N_9307);
nor UO_946 (O_946,N_9608,N_9460);
nor UO_947 (O_947,N_9852,N_9698);
nor UO_948 (O_948,N_9494,N_9156);
nor UO_949 (O_949,N_9672,N_9946);
and UO_950 (O_950,N_9987,N_9194);
and UO_951 (O_951,N_9538,N_9378);
nor UO_952 (O_952,N_9103,N_9130);
and UO_953 (O_953,N_9275,N_9684);
nand UO_954 (O_954,N_9393,N_9971);
nand UO_955 (O_955,N_9201,N_9987);
nand UO_956 (O_956,N_9593,N_9809);
or UO_957 (O_957,N_9530,N_9996);
nand UO_958 (O_958,N_9030,N_9862);
and UO_959 (O_959,N_9135,N_9936);
nand UO_960 (O_960,N_9215,N_9668);
nand UO_961 (O_961,N_9856,N_9990);
or UO_962 (O_962,N_9759,N_9242);
and UO_963 (O_963,N_9955,N_9021);
nand UO_964 (O_964,N_9818,N_9071);
xor UO_965 (O_965,N_9346,N_9610);
nor UO_966 (O_966,N_9030,N_9482);
or UO_967 (O_967,N_9260,N_9376);
and UO_968 (O_968,N_9476,N_9105);
nor UO_969 (O_969,N_9257,N_9863);
nor UO_970 (O_970,N_9892,N_9553);
or UO_971 (O_971,N_9166,N_9871);
and UO_972 (O_972,N_9594,N_9888);
or UO_973 (O_973,N_9073,N_9232);
and UO_974 (O_974,N_9263,N_9965);
and UO_975 (O_975,N_9917,N_9478);
nand UO_976 (O_976,N_9716,N_9681);
nor UO_977 (O_977,N_9552,N_9110);
nor UO_978 (O_978,N_9486,N_9626);
nor UO_979 (O_979,N_9222,N_9992);
and UO_980 (O_980,N_9426,N_9623);
nand UO_981 (O_981,N_9737,N_9261);
nand UO_982 (O_982,N_9503,N_9471);
or UO_983 (O_983,N_9544,N_9697);
and UO_984 (O_984,N_9228,N_9884);
nand UO_985 (O_985,N_9987,N_9641);
nor UO_986 (O_986,N_9894,N_9852);
nand UO_987 (O_987,N_9637,N_9511);
nand UO_988 (O_988,N_9720,N_9112);
and UO_989 (O_989,N_9890,N_9242);
nor UO_990 (O_990,N_9637,N_9308);
nand UO_991 (O_991,N_9833,N_9666);
nand UO_992 (O_992,N_9025,N_9065);
nand UO_993 (O_993,N_9907,N_9337);
and UO_994 (O_994,N_9105,N_9552);
nor UO_995 (O_995,N_9273,N_9039);
or UO_996 (O_996,N_9059,N_9642);
and UO_997 (O_997,N_9147,N_9754);
nand UO_998 (O_998,N_9106,N_9769);
nor UO_999 (O_999,N_9835,N_9693);
nand UO_1000 (O_1000,N_9397,N_9375);
nand UO_1001 (O_1001,N_9140,N_9062);
and UO_1002 (O_1002,N_9832,N_9927);
nor UO_1003 (O_1003,N_9782,N_9182);
nor UO_1004 (O_1004,N_9413,N_9150);
nor UO_1005 (O_1005,N_9902,N_9561);
and UO_1006 (O_1006,N_9650,N_9300);
and UO_1007 (O_1007,N_9258,N_9694);
or UO_1008 (O_1008,N_9216,N_9723);
nor UO_1009 (O_1009,N_9883,N_9252);
or UO_1010 (O_1010,N_9269,N_9549);
and UO_1011 (O_1011,N_9762,N_9213);
or UO_1012 (O_1012,N_9900,N_9601);
nand UO_1013 (O_1013,N_9161,N_9658);
or UO_1014 (O_1014,N_9674,N_9686);
nand UO_1015 (O_1015,N_9419,N_9306);
and UO_1016 (O_1016,N_9968,N_9846);
nand UO_1017 (O_1017,N_9790,N_9253);
or UO_1018 (O_1018,N_9031,N_9586);
and UO_1019 (O_1019,N_9798,N_9268);
nand UO_1020 (O_1020,N_9350,N_9976);
nand UO_1021 (O_1021,N_9881,N_9188);
or UO_1022 (O_1022,N_9700,N_9958);
or UO_1023 (O_1023,N_9207,N_9602);
or UO_1024 (O_1024,N_9250,N_9106);
or UO_1025 (O_1025,N_9639,N_9349);
or UO_1026 (O_1026,N_9217,N_9835);
or UO_1027 (O_1027,N_9603,N_9545);
nand UO_1028 (O_1028,N_9806,N_9396);
and UO_1029 (O_1029,N_9285,N_9131);
and UO_1030 (O_1030,N_9500,N_9020);
nor UO_1031 (O_1031,N_9465,N_9776);
nand UO_1032 (O_1032,N_9609,N_9529);
or UO_1033 (O_1033,N_9626,N_9202);
and UO_1034 (O_1034,N_9872,N_9941);
nand UO_1035 (O_1035,N_9874,N_9647);
nor UO_1036 (O_1036,N_9259,N_9094);
or UO_1037 (O_1037,N_9132,N_9372);
nor UO_1038 (O_1038,N_9365,N_9339);
and UO_1039 (O_1039,N_9818,N_9888);
or UO_1040 (O_1040,N_9749,N_9435);
or UO_1041 (O_1041,N_9587,N_9935);
and UO_1042 (O_1042,N_9518,N_9168);
xnor UO_1043 (O_1043,N_9319,N_9905);
nand UO_1044 (O_1044,N_9791,N_9920);
nor UO_1045 (O_1045,N_9847,N_9723);
nor UO_1046 (O_1046,N_9084,N_9179);
and UO_1047 (O_1047,N_9126,N_9808);
nor UO_1048 (O_1048,N_9760,N_9303);
xor UO_1049 (O_1049,N_9352,N_9188);
or UO_1050 (O_1050,N_9066,N_9968);
and UO_1051 (O_1051,N_9820,N_9662);
and UO_1052 (O_1052,N_9947,N_9339);
or UO_1053 (O_1053,N_9314,N_9353);
and UO_1054 (O_1054,N_9660,N_9722);
nor UO_1055 (O_1055,N_9043,N_9450);
nor UO_1056 (O_1056,N_9644,N_9351);
nand UO_1057 (O_1057,N_9632,N_9169);
or UO_1058 (O_1058,N_9993,N_9767);
and UO_1059 (O_1059,N_9464,N_9328);
nor UO_1060 (O_1060,N_9372,N_9699);
and UO_1061 (O_1061,N_9349,N_9445);
and UO_1062 (O_1062,N_9365,N_9048);
and UO_1063 (O_1063,N_9292,N_9661);
nand UO_1064 (O_1064,N_9589,N_9729);
or UO_1065 (O_1065,N_9468,N_9339);
and UO_1066 (O_1066,N_9987,N_9859);
or UO_1067 (O_1067,N_9381,N_9387);
nand UO_1068 (O_1068,N_9975,N_9611);
nor UO_1069 (O_1069,N_9260,N_9038);
or UO_1070 (O_1070,N_9089,N_9856);
nor UO_1071 (O_1071,N_9428,N_9229);
nand UO_1072 (O_1072,N_9897,N_9718);
or UO_1073 (O_1073,N_9186,N_9922);
nor UO_1074 (O_1074,N_9909,N_9850);
nand UO_1075 (O_1075,N_9677,N_9635);
or UO_1076 (O_1076,N_9277,N_9621);
and UO_1077 (O_1077,N_9023,N_9844);
or UO_1078 (O_1078,N_9347,N_9547);
nand UO_1079 (O_1079,N_9233,N_9910);
nor UO_1080 (O_1080,N_9033,N_9921);
or UO_1081 (O_1081,N_9598,N_9765);
nand UO_1082 (O_1082,N_9177,N_9730);
nor UO_1083 (O_1083,N_9946,N_9714);
or UO_1084 (O_1084,N_9768,N_9983);
nand UO_1085 (O_1085,N_9757,N_9261);
nand UO_1086 (O_1086,N_9091,N_9940);
and UO_1087 (O_1087,N_9083,N_9836);
or UO_1088 (O_1088,N_9902,N_9751);
and UO_1089 (O_1089,N_9366,N_9078);
or UO_1090 (O_1090,N_9062,N_9705);
and UO_1091 (O_1091,N_9189,N_9360);
and UO_1092 (O_1092,N_9583,N_9142);
nand UO_1093 (O_1093,N_9307,N_9520);
nand UO_1094 (O_1094,N_9295,N_9698);
or UO_1095 (O_1095,N_9426,N_9648);
nand UO_1096 (O_1096,N_9433,N_9726);
nor UO_1097 (O_1097,N_9715,N_9411);
nor UO_1098 (O_1098,N_9783,N_9127);
nand UO_1099 (O_1099,N_9681,N_9966);
and UO_1100 (O_1100,N_9016,N_9477);
and UO_1101 (O_1101,N_9018,N_9852);
nand UO_1102 (O_1102,N_9236,N_9406);
and UO_1103 (O_1103,N_9699,N_9219);
nand UO_1104 (O_1104,N_9371,N_9214);
and UO_1105 (O_1105,N_9387,N_9228);
or UO_1106 (O_1106,N_9183,N_9188);
nor UO_1107 (O_1107,N_9413,N_9871);
and UO_1108 (O_1108,N_9515,N_9326);
nor UO_1109 (O_1109,N_9630,N_9687);
nor UO_1110 (O_1110,N_9167,N_9295);
and UO_1111 (O_1111,N_9962,N_9035);
nor UO_1112 (O_1112,N_9162,N_9064);
or UO_1113 (O_1113,N_9539,N_9521);
and UO_1114 (O_1114,N_9736,N_9729);
and UO_1115 (O_1115,N_9317,N_9873);
nor UO_1116 (O_1116,N_9732,N_9716);
or UO_1117 (O_1117,N_9847,N_9536);
nand UO_1118 (O_1118,N_9820,N_9884);
xor UO_1119 (O_1119,N_9864,N_9080);
or UO_1120 (O_1120,N_9548,N_9482);
and UO_1121 (O_1121,N_9473,N_9744);
and UO_1122 (O_1122,N_9395,N_9570);
or UO_1123 (O_1123,N_9338,N_9466);
or UO_1124 (O_1124,N_9421,N_9597);
and UO_1125 (O_1125,N_9113,N_9690);
nand UO_1126 (O_1126,N_9731,N_9016);
and UO_1127 (O_1127,N_9071,N_9787);
and UO_1128 (O_1128,N_9031,N_9321);
or UO_1129 (O_1129,N_9983,N_9375);
nand UO_1130 (O_1130,N_9483,N_9203);
nand UO_1131 (O_1131,N_9077,N_9595);
or UO_1132 (O_1132,N_9408,N_9893);
and UO_1133 (O_1133,N_9526,N_9851);
or UO_1134 (O_1134,N_9458,N_9630);
nand UO_1135 (O_1135,N_9982,N_9098);
nor UO_1136 (O_1136,N_9234,N_9132);
nand UO_1137 (O_1137,N_9110,N_9403);
nand UO_1138 (O_1138,N_9431,N_9960);
nand UO_1139 (O_1139,N_9484,N_9817);
and UO_1140 (O_1140,N_9682,N_9440);
nand UO_1141 (O_1141,N_9257,N_9219);
nand UO_1142 (O_1142,N_9551,N_9399);
or UO_1143 (O_1143,N_9348,N_9698);
nor UO_1144 (O_1144,N_9847,N_9102);
nand UO_1145 (O_1145,N_9335,N_9686);
and UO_1146 (O_1146,N_9712,N_9828);
nand UO_1147 (O_1147,N_9730,N_9922);
nor UO_1148 (O_1148,N_9200,N_9164);
nand UO_1149 (O_1149,N_9696,N_9079);
and UO_1150 (O_1150,N_9808,N_9296);
and UO_1151 (O_1151,N_9288,N_9409);
nor UO_1152 (O_1152,N_9177,N_9108);
nand UO_1153 (O_1153,N_9007,N_9140);
xor UO_1154 (O_1154,N_9196,N_9335);
nor UO_1155 (O_1155,N_9067,N_9211);
nor UO_1156 (O_1156,N_9838,N_9284);
nand UO_1157 (O_1157,N_9559,N_9385);
and UO_1158 (O_1158,N_9097,N_9653);
nand UO_1159 (O_1159,N_9155,N_9477);
nand UO_1160 (O_1160,N_9814,N_9425);
or UO_1161 (O_1161,N_9050,N_9884);
or UO_1162 (O_1162,N_9100,N_9504);
or UO_1163 (O_1163,N_9119,N_9637);
and UO_1164 (O_1164,N_9177,N_9875);
nand UO_1165 (O_1165,N_9073,N_9812);
or UO_1166 (O_1166,N_9218,N_9217);
nor UO_1167 (O_1167,N_9618,N_9696);
nand UO_1168 (O_1168,N_9608,N_9872);
nand UO_1169 (O_1169,N_9075,N_9582);
nor UO_1170 (O_1170,N_9516,N_9976);
nand UO_1171 (O_1171,N_9409,N_9319);
nor UO_1172 (O_1172,N_9430,N_9173);
or UO_1173 (O_1173,N_9659,N_9528);
or UO_1174 (O_1174,N_9326,N_9680);
nor UO_1175 (O_1175,N_9923,N_9145);
nand UO_1176 (O_1176,N_9991,N_9322);
and UO_1177 (O_1177,N_9277,N_9784);
or UO_1178 (O_1178,N_9832,N_9904);
or UO_1179 (O_1179,N_9403,N_9919);
and UO_1180 (O_1180,N_9820,N_9539);
nor UO_1181 (O_1181,N_9457,N_9482);
nor UO_1182 (O_1182,N_9396,N_9353);
or UO_1183 (O_1183,N_9239,N_9103);
or UO_1184 (O_1184,N_9084,N_9656);
and UO_1185 (O_1185,N_9868,N_9491);
or UO_1186 (O_1186,N_9054,N_9437);
nor UO_1187 (O_1187,N_9457,N_9288);
nor UO_1188 (O_1188,N_9671,N_9618);
nor UO_1189 (O_1189,N_9932,N_9773);
nand UO_1190 (O_1190,N_9485,N_9774);
nand UO_1191 (O_1191,N_9386,N_9242);
nor UO_1192 (O_1192,N_9532,N_9825);
or UO_1193 (O_1193,N_9219,N_9163);
nand UO_1194 (O_1194,N_9877,N_9965);
or UO_1195 (O_1195,N_9758,N_9008);
or UO_1196 (O_1196,N_9082,N_9990);
or UO_1197 (O_1197,N_9562,N_9265);
and UO_1198 (O_1198,N_9890,N_9437);
and UO_1199 (O_1199,N_9167,N_9498);
nor UO_1200 (O_1200,N_9415,N_9659);
or UO_1201 (O_1201,N_9659,N_9156);
nand UO_1202 (O_1202,N_9351,N_9188);
nand UO_1203 (O_1203,N_9935,N_9801);
and UO_1204 (O_1204,N_9736,N_9953);
nand UO_1205 (O_1205,N_9527,N_9076);
or UO_1206 (O_1206,N_9147,N_9971);
nand UO_1207 (O_1207,N_9882,N_9021);
and UO_1208 (O_1208,N_9758,N_9815);
or UO_1209 (O_1209,N_9431,N_9466);
nand UO_1210 (O_1210,N_9902,N_9956);
nand UO_1211 (O_1211,N_9857,N_9168);
nor UO_1212 (O_1212,N_9383,N_9287);
or UO_1213 (O_1213,N_9889,N_9350);
nand UO_1214 (O_1214,N_9753,N_9815);
and UO_1215 (O_1215,N_9515,N_9484);
and UO_1216 (O_1216,N_9483,N_9053);
and UO_1217 (O_1217,N_9680,N_9672);
nor UO_1218 (O_1218,N_9008,N_9528);
and UO_1219 (O_1219,N_9138,N_9369);
nor UO_1220 (O_1220,N_9416,N_9556);
nand UO_1221 (O_1221,N_9651,N_9733);
and UO_1222 (O_1222,N_9727,N_9905);
nand UO_1223 (O_1223,N_9841,N_9263);
or UO_1224 (O_1224,N_9420,N_9759);
or UO_1225 (O_1225,N_9108,N_9488);
nand UO_1226 (O_1226,N_9744,N_9384);
nor UO_1227 (O_1227,N_9424,N_9062);
and UO_1228 (O_1228,N_9638,N_9274);
and UO_1229 (O_1229,N_9913,N_9508);
and UO_1230 (O_1230,N_9911,N_9706);
and UO_1231 (O_1231,N_9552,N_9579);
or UO_1232 (O_1232,N_9284,N_9658);
and UO_1233 (O_1233,N_9100,N_9650);
or UO_1234 (O_1234,N_9433,N_9645);
nand UO_1235 (O_1235,N_9044,N_9102);
nand UO_1236 (O_1236,N_9508,N_9333);
nor UO_1237 (O_1237,N_9479,N_9184);
or UO_1238 (O_1238,N_9733,N_9852);
and UO_1239 (O_1239,N_9668,N_9814);
or UO_1240 (O_1240,N_9539,N_9666);
or UO_1241 (O_1241,N_9242,N_9258);
nor UO_1242 (O_1242,N_9298,N_9235);
and UO_1243 (O_1243,N_9684,N_9913);
and UO_1244 (O_1244,N_9068,N_9996);
or UO_1245 (O_1245,N_9369,N_9874);
nand UO_1246 (O_1246,N_9811,N_9000);
and UO_1247 (O_1247,N_9959,N_9839);
nand UO_1248 (O_1248,N_9817,N_9048);
and UO_1249 (O_1249,N_9494,N_9915);
and UO_1250 (O_1250,N_9018,N_9030);
and UO_1251 (O_1251,N_9904,N_9580);
and UO_1252 (O_1252,N_9195,N_9302);
nand UO_1253 (O_1253,N_9829,N_9283);
or UO_1254 (O_1254,N_9059,N_9724);
nor UO_1255 (O_1255,N_9336,N_9026);
nor UO_1256 (O_1256,N_9437,N_9556);
nand UO_1257 (O_1257,N_9410,N_9703);
and UO_1258 (O_1258,N_9392,N_9844);
and UO_1259 (O_1259,N_9811,N_9570);
and UO_1260 (O_1260,N_9628,N_9679);
nand UO_1261 (O_1261,N_9993,N_9189);
and UO_1262 (O_1262,N_9654,N_9195);
nand UO_1263 (O_1263,N_9703,N_9279);
nor UO_1264 (O_1264,N_9488,N_9682);
or UO_1265 (O_1265,N_9630,N_9138);
nand UO_1266 (O_1266,N_9114,N_9903);
nor UO_1267 (O_1267,N_9709,N_9081);
or UO_1268 (O_1268,N_9557,N_9841);
nor UO_1269 (O_1269,N_9966,N_9367);
nand UO_1270 (O_1270,N_9105,N_9807);
nand UO_1271 (O_1271,N_9952,N_9044);
nor UO_1272 (O_1272,N_9183,N_9490);
nand UO_1273 (O_1273,N_9370,N_9710);
nand UO_1274 (O_1274,N_9598,N_9508);
or UO_1275 (O_1275,N_9542,N_9227);
or UO_1276 (O_1276,N_9902,N_9230);
nand UO_1277 (O_1277,N_9565,N_9778);
and UO_1278 (O_1278,N_9730,N_9914);
nand UO_1279 (O_1279,N_9217,N_9099);
nand UO_1280 (O_1280,N_9520,N_9516);
or UO_1281 (O_1281,N_9835,N_9556);
nor UO_1282 (O_1282,N_9555,N_9475);
or UO_1283 (O_1283,N_9382,N_9383);
xnor UO_1284 (O_1284,N_9783,N_9444);
nor UO_1285 (O_1285,N_9343,N_9643);
nand UO_1286 (O_1286,N_9708,N_9462);
nand UO_1287 (O_1287,N_9160,N_9661);
nand UO_1288 (O_1288,N_9944,N_9384);
nand UO_1289 (O_1289,N_9509,N_9977);
nor UO_1290 (O_1290,N_9615,N_9590);
and UO_1291 (O_1291,N_9689,N_9421);
nand UO_1292 (O_1292,N_9386,N_9748);
or UO_1293 (O_1293,N_9590,N_9620);
or UO_1294 (O_1294,N_9634,N_9986);
and UO_1295 (O_1295,N_9751,N_9346);
and UO_1296 (O_1296,N_9482,N_9365);
and UO_1297 (O_1297,N_9916,N_9052);
nand UO_1298 (O_1298,N_9695,N_9530);
and UO_1299 (O_1299,N_9396,N_9584);
or UO_1300 (O_1300,N_9024,N_9295);
nor UO_1301 (O_1301,N_9922,N_9559);
and UO_1302 (O_1302,N_9677,N_9212);
and UO_1303 (O_1303,N_9719,N_9350);
and UO_1304 (O_1304,N_9908,N_9569);
and UO_1305 (O_1305,N_9442,N_9240);
nor UO_1306 (O_1306,N_9138,N_9056);
nand UO_1307 (O_1307,N_9324,N_9576);
xnor UO_1308 (O_1308,N_9996,N_9615);
nand UO_1309 (O_1309,N_9762,N_9435);
and UO_1310 (O_1310,N_9753,N_9166);
nor UO_1311 (O_1311,N_9425,N_9924);
or UO_1312 (O_1312,N_9784,N_9067);
nor UO_1313 (O_1313,N_9022,N_9955);
nor UO_1314 (O_1314,N_9283,N_9672);
nor UO_1315 (O_1315,N_9124,N_9841);
or UO_1316 (O_1316,N_9763,N_9589);
and UO_1317 (O_1317,N_9706,N_9712);
nor UO_1318 (O_1318,N_9796,N_9709);
nor UO_1319 (O_1319,N_9478,N_9084);
nand UO_1320 (O_1320,N_9759,N_9593);
nand UO_1321 (O_1321,N_9289,N_9334);
or UO_1322 (O_1322,N_9852,N_9467);
and UO_1323 (O_1323,N_9722,N_9843);
nor UO_1324 (O_1324,N_9639,N_9982);
nor UO_1325 (O_1325,N_9271,N_9092);
and UO_1326 (O_1326,N_9399,N_9930);
and UO_1327 (O_1327,N_9688,N_9952);
and UO_1328 (O_1328,N_9860,N_9988);
nor UO_1329 (O_1329,N_9502,N_9328);
or UO_1330 (O_1330,N_9139,N_9917);
and UO_1331 (O_1331,N_9764,N_9161);
and UO_1332 (O_1332,N_9104,N_9112);
nand UO_1333 (O_1333,N_9708,N_9859);
nand UO_1334 (O_1334,N_9572,N_9288);
or UO_1335 (O_1335,N_9595,N_9569);
nand UO_1336 (O_1336,N_9656,N_9004);
or UO_1337 (O_1337,N_9876,N_9068);
or UO_1338 (O_1338,N_9402,N_9944);
nand UO_1339 (O_1339,N_9493,N_9094);
nand UO_1340 (O_1340,N_9750,N_9866);
and UO_1341 (O_1341,N_9737,N_9504);
nand UO_1342 (O_1342,N_9414,N_9720);
and UO_1343 (O_1343,N_9970,N_9618);
or UO_1344 (O_1344,N_9802,N_9638);
or UO_1345 (O_1345,N_9763,N_9203);
nor UO_1346 (O_1346,N_9286,N_9891);
nand UO_1347 (O_1347,N_9183,N_9021);
and UO_1348 (O_1348,N_9770,N_9571);
or UO_1349 (O_1349,N_9705,N_9812);
nand UO_1350 (O_1350,N_9197,N_9381);
nor UO_1351 (O_1351,N_9772,N_9375);
nand UO_1352 (O_1352,N_9860,N_9609);
and UO_1353 (O_1353,N_9421,N_9950);
or UO_1354 (O_1354,N_9248,N_9078);
xor UO_1355 (O_1355,N_9507,N_9087);
nor UO_1356 (O_1356,N_9242,N_9888);
or UO_1357 (O_1357,N_9599,N_9990);
nand UO_1358 (O_1358,N_9962,N_9218);
nand UO_1359 (O_1359,N_9041,N_9679);
xor UO_1360 (O_1360,N_9817,N_9551);
and UO_1361 (O_1361,N_9623,N_9383);
or UO_1362 (O_1362,N_9455,N_9522);
nor UO_1363 (O_1363,N_9937,N_9874);
and UO_1364 (O_1364,N_9367,N_9812);
and UO_1365 (O_1365,N_9062,N_9640);
nand UO_1366 (O_1366,N_9520,N_9534);
nor UO_1367 (O_1367,N_9085,N_9849);
nand UO_1368 (O_1368,N_9261,N_9019);
nand UO_1369 (O_1369,N_9030,N_9114);
or UO_1370 (O_1370,N_9379,N_9389);
nand UO_1371 (O_1371,N_9909,N_9831);
or UO_1372 (O_1372,N_9044,N_9898);
nand UO_1373 (O_1373,N_9444,N_9816);
or UO_1374 (O_1374,N_9111,N_9673);
nand UO_1375 (O_1375,N_9690,N_9184);
nand UO_1376 (O_1376,N_9445,N_9590);
and UO_1377 (O_1377,N_9866,N_9544);
or UO_1378 (O_1378,N_9570,N_9463);
nand UO_1379 (O_1379,N_9456,N_9395);
and UO_1380 (O_1380,N_9446,N_9851);
nand UO_1381 (O_1381,N_9560,N_9898);
or UO_1382 (O_1382,N_9454,N_9891);
nand UO_1383 (O_1383,N_9425,N_9267);
and UO_1384 (O_1384,N_9684,N_9390);
nor UO_1385 (O_1385,N_9591,N_9107);
nand UO_1386 (O_1386,N_9557,N_9756);
nand UO_1387 (O_1387,N_9394,N_9631);
and UO_1388 (O_1388,N_9490,N_9371);
or UO_1389 (O_1389,N_9054,N_9474);
and UO_1390 (O_1390,N_9231,N_9854);
and UO_1391 (O_1391,N_9247,N_9932);
nor UO_1392 (O_1392,N_9995,N_9483);
nor UO_1393 (O_1393,N_9715,N_9265);
or UO_1394 (O_1394,N_9298,N_9324);
nand UO_1395 (O_1395,N_9339,N_9911);
or UO_1396 (O_1396,N_9028,N_9557);
nor UO_1397 (O_1397,N_9092,N_9008);
and UO_1398 (O_1398,N_9494,N_9003);
nor UO_1399 (O_1399,N_9771,N_9098);
nand UO_1400 (O_1400,N_9516,N_9395);
or UO_1401 (O_1401,N_9693,N_9944);
or UO_1402 (O_1402,N_9754,N_9522);
nand UO_1403 (O_1403,N_9314,N_9471);
nand UO_1404 (O_1404,N_9255,N_9930);
nand UO_1405 (O_1405,N_9652,N_9077);
and UO_1406 (O_1406,N_9578,N_9488);
nand UO_1407 (O_1407,N_9192,N_9928);
nor UO_1408 (O_1408,N_9941,N_9853);
or UO_1409 (O_1409,N_9668,N_9510);
or UO_1410 (O_1410,N_9170,N_9606);
or UO_1411 (O_1411,N_9703,N_9087);
nor UO_1412 (O_1412,N_9162,N_9413);
or UO_1413 (O_1413,N_9965,N_9797);
nand UO_1414 (O_1414,N_9711,N_9968);
xor UO_1415 (O_1415,N_9141,N_9793);
nor UO_1416 (O_1416,N_9367,N_9599);
nand UO_1417 (O_1417,N_9047,N_9277);
and UO_1418 (O_1418,N_9566,N_9412);
nor UO_1419 (O_1419,N_9068,N_9537);
or UO_1420 (O_1420,N_9391,N_9228);
and UO_1421 (O_1421,N_9109,N_9560);
or UO_1422 (O_1422,N_9823,N_9368);
and UO_1423 (O_1423,N_9264,N_9135);
and UO_1424 (O_1424,N_9983,N_9361);
nand UO_1425 (O_1425,N_9720,N_9748);
or UO_1426 (O_1426,N_9545,N_9795);
and UO_1427 (O_1427,N_9602,N_9856);
xor UO_1428 (O_1428,N_9729,N_9242);
nand UO_1429 (O_1429,N_9468,N_9157);
or UO_1430 (O_1430,N_9435,N_9614);
and UO_1431 (O_1431,N_9926,N_9341);
nor UO_1432 (O_1432,N_9059,N_9097);
or UO_1433 (O_1433,N_9118,N_9588);
and UO_1434 (O_1434,N_9877,N_9481);
or UO_1435 (O_1435,N_9508,N_9004);
or UO_1436 (O_1436,N_9029,N_9053);
nor UO_1437 (O_1437,N_9838,N_9189);
nand UO_1438 (O_1438,N_9974,N_9481);
or UO_1439 (O_1439,N_9162,N_9532);
and UO_1440 (O_1440,N_9932,N_9541);
nand UO_1441 (O_1441,N_9647,N_9617);
or UO_1442 (O_1442,N_9141,N_9858);
or UO_1443 (O_1443,N_9575,N_9902);
and UO_1444 (O_1444,N_9451,N_9901);
and UO_1445 (O_1445,N_9763,N_9370);
or UO_1446 (O_1446,N_9598,N_9412);
and UO_1447 (O_1447,N_9009,N_9289);
nor UO_1448 (O_1448,N_9152,N_9241);
nand UO_1449 (O_1449,N_9849,N_9225);
nand UO_1450 (O_1450,N_9049,N_9960);
and UO_1451 (O_1451,N_9774,N_9400);
nor UO_1452 (O_1452,N_9619,N_9233);
and UO_1453 (O_1453,N_9473,N_9614);
nand UO_1454 (O_1454,N_9709,N_9512);
or UO_1455 (O_1455,N_9356,N_9239);
nand UO_1456 (O_1456,N_9629,N_9169);
nand UO_1457 (O_1457,N_9959,N_9932);
or UO_1458 (O_1458,N_9858,N_9143);
or UO_1459 (O_1459,N_9178,N_9201);
nand UO_1460 (O_1460,N_9172,N_9464);
xor UO_1461 (O_1461,N_9586,N_9486);
and UO_1462 (O_1462,N_9766,N_9762);
and UO_1463 (O_1463,N_9439,N_9435);
xnor UO_1464 (O_1464,N_9109,N_9555);
and UO_1465 (O_1465,N_9861,N_9706);
nor UO_1466 (O_1466,N_9419,N_9885);
and UO_1467 (O_1467,N_9330,N_9439);
nand UO_1468 (O_1468,N_9688,N_9379);
xnor UO_1469 (O_1469,N_9378,N_9444);
nand UO_1470 (O_1470,N_9708,N_9751);
nand UO_1471 (O_1471,N_9509,N_9414);
and UO_1472 (O_1472,N_9200,N_9342);
and UO_1473 (O_1473,N_9742,N_9787);
and UO_1474 (O_1474,N_9893,N_9039);
nor UO_1475 (O_1475,N_9319,N_9088);
or UO_1476 (O_1476,N_9569,N_9586);
and UO_1477 (O_1477,N_9817,N_9501);
or UO_1478 (O_1478,N_9410,N_9296);
and UO_1479 (O_1479,N_9531,N_9113);
and UO_1480 (O_1480,N_9954,N_9636);
nand UO_1481 (O_1481,N_9413,N_9414);
and UO_1482 (O_1482,N_9496,N_9368);
or UO_1483 (O_1483,N_9475,N_9504);
nor UO_1484 (O_1484,N_9440,N_9645);
and UO_1485 (O_1485,N_9715,N_9374);
nand UO_1486 (O_1486,N_9397,N_9985);
or UO_1487 (O_1487,N_9198,N_9413);
and UO_1488 (O_1488,N_9442,N_9580);
and UO_1489 (O_1489,N_9649,N_9302);
nand UO_1490 (O_1490,N_9061,N_9575);
or UO_1491 (O_1491,N_9763,N_9900);
or UO_1492 (O_1492,N_9957,N_9420);
and UO_1493 (O_1493,N_9642,N_9516);
nand UO_1494 (O_1494,N_9247,N_9482);
nand UO_1495 (O_1495,N_9673,N_9933);
nor UO_1496 (O_1496,N_9164,N_9779);
nor UO_1497 (O_1497,N_9515,N_9132);
nor UO_1498 (O_1498,N_9906,N_9164);
or UO_1499 (O_1499,N_9852,N_9989);
endmodule