module basic_500_3000_500_60_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
xor U0 (N_0,In_20,In_102);
xnor U1 (N_1,In_130,In_351);
nand U2 (N_2,In_462,In_443);
or U3 (N_3,In_84,In_136);
and U4 (N_4,In_425,In_1);
or U5 (N_5,In_192,In_196);
and U6 (N_6,In_430,In_170);
nand U7 (N_7,In_458,In_202);
xnor U8 (N_8,In_143,In_244);
xor U9 (N_9,In_495,In_68);
and U10 (N_10,In_426,In_375);
nor U11 (N_11,In_14,In_228);
or U12 (N_12,In_121,In_257);
nor U13 (N_13,In_156,In_155);
xnor U14 (N_14,In_493,In_201);
or U15 (N_15,In_492,In_129);
and U16 (N_16,In_22,In_62);
and U17 (N_17,In_260,In_75);
nand U18 (N_18,In_127,In_447);
or U19 (N_19,In_453,In_281);
nor U20 (N_20,In_176,In_388);
and U21 (N_21,In_498,In_463);
and U22 (N_22,In_397,In_165);
and U23 (N_23,In_284,In_308);
and U24 (N_24,In_368,In_496);
or U25 (N_25,In_317,In_67);
nor U26 (N_26,In_344,In_103);
or U27 (N_27,In_26,In_210);
nor U28 (N_28,In_51,In_389);
or U29 (N_29,In_421,In_441);
xor U30 (N_30,In_36,In_262);
nor U31 (N_31,In_60,In_207);
xnor U32 (N_32,In_444,In_174);
nand U33 (N_33,In_96,In_229);
nor U34 (N_34,In_213,In_348);
nand U35 (N_35,In_97,In_374);
xnor U36 (N_36,In_399,In_474);
or U37 (N_37,In_195,In_34);
and U38 (N_38,In_172,In_57);
nand U39 (N_39,In_190,In_298);
xnor U40 (N_40,In_25,In_381);
or U41 (N_41,In_413,In_488);
xor U42 (N_42,In_6,In_332);
or U43 (N_43,In_232,In_132);
nand U44 (N_44,In_52,In_433);
nor U45 (N_45,In_261,In_47);
or U46 (N_46,In_114,In_414);
nor U47 (N_47,In_352,In_149);
nand U48 (N_48,In_442,In_289);
nand U49 (N_49,In_99,In_146);
or U50 (N_50,In_341,In_40);
and U51 (N_51,In_336,In_116);
or U52 (N_52,N_7,In_98);
xor U53 (N_53,In_320,In_445);
xnor U54 (N_54,In_459,In_131);
nor U55 (N_55,In_358,In_247);
and U56 (N_56,In_88,In_391);
xnor U57 (N_57,In_226,In_119);
and U58 (N_58,In_386,In_70);
nand U59 (N_59,In_206,In_380);
nor U60 (N_60,In_71,In_392);
xor U61 (N_61,In_489,In_145);
nor U62 (N_62,In_328,In_407);
xnor U63 (N_63,In_243,In_385);
nand U64 (N_64,In_301,In_265);
or U65 (N_65,In_299,In_266);
nor U66 (N_66,In_58,In_59);
or U67 (N_67,In_187,In_66);
nand U68 (N_68,In_471,In_377);
nor U69 (N_69,In_238,In_152);
nor U70 (N_70,In_168,In_258);
nor U71 (N_71,N_5,In_406);
or U72 (N_72,N_17,In_420);
or U73 (N_73,In_241,In_282);
and U74 (N_74,In_74,In_429);
nand U75 (N_75,In_38,In_402);
or U76 (N_76,In_360,In_365);
nand U77 (N_77,In_147,In_248);
nand U78 (N_78,In_113,N_37);
xor U79 (N_79,In_315,N_22);
and U80 (N_80,In_55,In_109);
nand U81 (N_81,In_366,In_126);
nand U82 (N_82,In_294,In_218);
xor U83 (N_83,In_154,In_356);
nor U84 (N_84,In_461,In_200);
nor U85 (N_85,In_321,In_82);
and U86 (N_86,In_259,In_390);
and U87 (N_87,In_279,In_69);
or U88 (N_88,In_403,In_65);
nand U89 (N_89,In_27,In_111);
nand U90 (N_90,In_189,In_456);
or U91 (N_91,In_92,In_475);
or U92 (N_92,In_337,In_4);
nand U93 (N_93,In_237,In_467);
nor U94 (N_94,N_49,In_494);
nand U95 (N_95,In_326,In_45);
nand U96 (N_96,N_18,N_46);
or U97 (N_97,In_292,In_423);
or U98 (N_98,In_437,In_411);
nand U99 (N_99,In_269,In_184);
or U100 (N_100,In_8,N_90);
or U101 (N_101,N_1,In_303);
nand U102 (N_102,In_327,N_3);
and U103 (N_103,In_466,In_353);
xnor U104 (N_104,In_482,In_280);
xnor U105 (N_105,N_68,In_80);
nand U106 (N_106,N_86,In_329);
or U107 (N_107,In_387,N_71);
nand U108 (N_108,In_177,In_86);
nand U109 (N_109,In_295,In_63);
nand U110 (N_110,In_370,In_138);
and U111 (N_111,In_340,N_74);
and U112 (N_112,In_164,In_29);
or U113 (N_113,N_95,In_204);
nand U114 (N_114,In_50,In_7);
or U115 (N_115,In_49,In_401);
nand U116 (N_116,In_450,In_77);
and U117 (N_117,In_311,In_212);
nor U118 (N_118,N_55,N_34);
and U119 (N_119,In_240,N_67);
nor U120 (N_120,In_438,In_137);
nand U121 (N_121,In_185,In_322);
nor U122 (N_122,In_373,In_118);
nor U123 (N_123,In_44,N_36);
and U124 (N_124,In_231,N_52);
xnor U125 (N_125,N_10,N_72);
or U126 (N_126,In_215,In_427);
nand U127 (N_127,In_393,In_287);
xnor U128 (N_128,N_65,N_2);
nand U129 (N_129,N_24,In_361);
and U130 (N_130,In_179,In_251);
nand U131 (N_131,In_225,In_300);
or U132 (N_132,In_197,In_150);
xor U133 (N_133,N_87,In_307);
nand U134 (N_134,In_46,N_33);
nand U135 (N_135,In_349,In_53);
nor U136 (N_136,In_404,In_408);
or U137 (N_137,In_452,In_424);
xnor U138 (N_138,N_83,In_419);
nor U139 (N_139,N_75,N_97);
nor U140 (N_140,In_310,In_305);
and U141 (N_141,In_478,In_335);
and U142 (N_142,In_64,N_93);
nor U143 (N_143,In_128,In_276);
and U144 (N_144,In_314,In_448);
nand U145 (N_145,In_440,In_338);
and U146 (N_146,In_472,In_319);
or U147 (N_147,N_57,In_333);
xnor U148 (N_148,In_357,In_30);
or U149 (N_149,In_270,In_283);
nor U150 (N_150,N_119,N_32);
or U151 (N_151,N_47,In_108);
xor U152 (N_152,In_33,In_249);
nand U153 (N_153,In_93,N_107);
nand U154 (N_154,In_431,N_133);
and U155 (N_155,In_306,In_94);
nor U156 (N_156,N_130,In_85);
and U157 (N_157,In_369,N_63);
or U158 (N_158,In_334,In_476);
xnor U159 (N_159,N_113,N_15);
or U160 (N_160,In_87,N_134);
nor U161 (N_161,In_372,In_123);
or U162 (N_162,In_73,N_85);
nand U163 (N_163,In_78,In_479);
xnor U164 (N_164,In_21,N_42);
nand U165 (N_165,N_135,In_417);
nor U166 (N_166,In_37,N_105);
nor U167 (N_167,In_48,In_439);
or U168 (N_168,N_13,N_144);
and U169 (N_169,In_346,N_124);
nand U170 (N_170,In_139,In_10);
or U171 (N_171,In_160,N_111);
nor U172 (N_172,In_0,N_127);
or U173 (N_173,In_362,In_39);
nor U174 (N_174,N_51,N_120);
nor U175 (N_175,N_138,In_454);
nand U176 (N_176,In_480,In_436);
and U177 (N_177,In_290,In_418);
nor U178 (N_178,N_145,N_28);
and U179 (N_179,In_394,In_81);
nand U180 (N_180,N_30,N_35);
nand U181 (N_181,N_62,In_432);
and U182 (N_182,In_24,In_239);
nor U183 (N_183,In_455,In_378);
and U184 (N_184,In_91,N_140);
nand U185 (N_185,In_151,In_460);
nand U186 (N_186,In_41,In_167);
or U187 (N_187,In_297,In_120);
xor U188 (N_188,In_485,In_469);
and U189 (N_189,In_487,In_106);
nor U190 (N_190,In_457,In_79);
and U191 (N_191,In_293,In_263);
nand U192 (N_192,In_203,N_27);
and U193 (N_193,In_112,In_219);
nor U194 (N_194,In_140,In_400);
and U195 (N_195,In_18,N_45);
or U196 (N_196,In_209,In_468);
nand U197 (N_197,In_451,In_9);
nor U198 (N_198,N_136,In_199);
nor U199 (N_199,In_43,In_288);
or U200 (N_200,In_31,N_160);
nor U201 (N_201,N_38,N_158);
xnor U202 (N_202,N_16,N_195);
or U203 (N_203,In_465,In_235);
xor U204 (N_204,N_64,N_0);
nor U205 (N_205,In_233,In_144);
nand U206 (N_206,N_26,In_278);
or U207 (N_207,N_94,In_182);
nand U208 (N_208,N_80,N_54);
nor U209 (N_209,N_141,In_323);
and U210 (N_210,In_23,In_312);
xnor U211 (N_211,N_70,N_9);
and U212 (N_212,N_188,In_271);
nor U213 (N_213,In_224,In_83);
and U214 (N_214,In_256,In_234);
or U215 (N_215,In_347,N_50);
and U216 (N_216,In_17,N_194);
nand U217 (N_217,In_286,In_19);
and U218 (N_218,In_175,In_161);
xnor U219 (N_219,N_132,In_110);
nand U220 (N_220,In_221,In_296);
xor U221 (N_221,In_169,N_175);
nand U222 (N_222,In_350,In_250);
or U223 (N_223,N_154,N_76);
and U224 (N_224,In_28,N_29);
xnor U225 (N_225,In_194,N_155);
and U226 (N_226,In_267,N_12);
xor U227 (N_227,In_236,In_343);
xor U228 (N_228,In_90,N_79);
or U229 (N_229,N_149,N_123);
and U230 (N_230,In_355,In_302);
nand U231 (N_231,In_217,In_148);
and U232 (N_232,N_125,N_108);
nor U233 (N_233,In_227,In_470);
nand U234 (N_234,In_324,In_483);
or U235 (N_235,In_273,N_176);
nand U236 (N_236,N_131,N_59);
nand U237 (N_237,N_147,In_473);
nor U238 (N_238,In_122,In_412);
nor U239 (N_239,In_13,In_277);
or U240 (N_240,N_117,N_43);
and U241 (N_241,In_422,N_143);
nand U242 (N_242,In_274,N_106);
and U243 (N_243,In_216,In_331);
xor U244 (N_244,N_21,In_354);
xnor U245 (N_245,In_379,N_6);
or U246 (N_246,N_4,N_181);
and U247 (N_247,In_61,N_150);
nor U248 (N_248,N_166,N_19);
nand U249 (N_249,In_383,N_137);
nor U250 (N_250,N_161,In_5);
or U251 (N_251,N_239,N_204);
nand U252 (N_252,N_179,In_107);
xor U253 (N_253,In_464,N_217);
xor U254 (N_254,In_499,In_124);
xnor U255 (N_255,N_234,In_434);
or U256 (N_256,N_248,N_193);
or U257 (N_257,In_325,N_172);
and U258 (N_258,N_128,N_157);
xor U259 (N_259,N_225,N_218);
nand U260 (N_260,In_125,N_58);
and U261 (N_261,N_199,N_103);
and U262 (N_262,In_198,N_249);
xor U263 (N_263,In_264,In_481);
xor U264 (N_264,N_84,N_220);
and U265 (N_265,In_376,N_182);
nor U266 (N_266,In_76,N_99);
nor U267 (N_267,In_268,In_491);
or U268 (N_268,In_398,In_446);
or U269 (N_269,In_115,In_32);
xnor U270 (N_270,In_316,In_95);
or U271 (N_271,N_228,In_72);
or U272 (N_272,N_196,In_410);
nor U273 (N_273,N_78,N_48);
xnor U274 (N_274,N_142,N_198);
nor U275 (N_275,N_209,In_180);
nor U276 (N_276,N_39,In_382);
and U277 (N_277,N_114,In_428);
or U278 (N_278,N_243,N_109);
and U279 (N_279,N_23,In_313);
or U280 (N_280,N_214,N_183);
and U281 (N_281,In_371,In_158);
or U282 (N_282,In_181,In_211);
and U283 (N_283,In_220,N_186);
xor U284 (N_284,N_213,N_192);
and U285 (N_285,In_157,In_100);
xnor U286 (N_286,N_98,N_205);
or U287 (N_287,In_395,N_92);
and U288 (N_288,In_272,N_245);
or U289 (N_289,In_166,N_241);
xnor U290 (N_290,N_210,N_14);
and U291 (N_291,N_118,N_216);
nor U292 (N_292,N_153,N_115);
nor U293 (N_293,N_231,In_497);
nor U294 (N_294,In_104,In_242);
or U295 (N_295,N_100,In_384);
xnor U296 (N_296,N_41,N_20);
and U297 (N_297,N_44,N_236);
and U298 (N_298,In_153,N_201);
nand U299 (N_299,N_116,N_156);
or U300 (N_300,N_206,N_298);
and U301 (N_301,In_142,N_223);
or U302 (N_302,In_409,N_233);
nor U303 (N_303,N_256,In_162);
or U304 (N_304,N_282,N_173);
and U305 (N_305,N_263,In_178);
and U306 (N_306,N_180,N_191);
or U307 (N_307,In_214,N_290);
xnor U308 (N_308,N_238,N_81);
and U309 (N_309,N_292,In_183);
nand U310 (N_310,N_274,N_276);
nor U311 (N_311,In_133,In_117);
xor U312 (N_312,N_89,N_8);
xnor U313 (N_313,N_221,N_289);
nor U314 (N_314,In_3,N_227);
nor U315 (N_315,N_178,N_184);
nand U316 (N_316,N_82,N_247);
and U317 (N_317,In_253,N_163);
xnor U318 (N_318,In_364,N_104);
or U319 (N_319,In_435,N_271);
and U320 (N_320,N_185,N_200);
nor U321 (N_321,In_405,N_171);
xor U322 (N_322,N_129,In_230);
or U323 (N_323,N_40,N_61);
nor U324 (N_324,N_31,N_283);
nor U325 (N_325,N_284,N_294);
nand U326 (N_326,N_164,N_257);
nand U327 (N_327,In_291,N_258);
nand U328 (N_328,N_25,N_229);
or U329 (N_329,In_367,N_286);
nand U330 (N_330,N_56,N_169);
xnor U331 (N_331,N_268,N_212);
or U332 (N_332,In_309,In_135);
xor U333 (N_333,In_252,In_339);
and U334 (N_334,N_224,N_159);
xnor U335 (N_335,In_56,In_191);
and U336 (N_336,N_165,N_237);
or U337 (N_337,N_146,N_207);
nor U338 (N_338,N_177,In_186);
nor U339 (N_339,N_272,N_190);
nand U340 (N_340,In_35,N_297);
xnor U341 (N_341,N_168,N_270);
nand U342 (N_342,In_415,N_91);
or U343 (N_343,In_396,N_287);
nand U344 (N_344,N_11,In_304);
or U345 (N_345,N_232,N_202);
or U346 (N_346,In_359,N_250);
xnor U347 (N_347,In_101,N_264);
or U348 (N_348,In_449,N_255);
xor U349 (N_349,In_12,N_152);
nor U350 (N_350,N_279,N_267);
or U351 (N_351,In_193,N_328);
and U352 (N_352,N_262,N_208);
xor U353 (N_353,N_312,N_295);
nor U354 (N_354,N_299,N_110);
xor U355 (N_355,N_322,N_317);
xnor U356 (N_356,In_345,N_242);
or U357 (N_357,N_189,In_484);
nand U358 (N_358,N_318,N_174);
or U359 (N_359,N_344,N_162);
nand U360 (N_360,N_309,In_330);
nand U361 (N_361,N_261,N_341);
nand U362 (N_362,N_246,N_337);
nor U363 (N_363,N_230,N_333);
and U364 (N_364,N_313,In_141);
nor U365 (N_365,N_269,In_477);
xor U366 (N_366,In_105,N_323);
nor U367 (N_367,N_88,N_251);
or U368 (N_368,N_307,N_266);
and U369 (N_369,N_336,N_167);
nor U370 (N_370,N_219,N_170);
or U371 (N_371,N_347,N_260);
nor U372 (N_372,In_486,N_112);
xor U373 (N_373,In_11,N_329);
nor U374 (N_374,N_296,In_255);
or U375 (N_375,N_222,N_197);
nor U376 (N_376,N_281,In_342);
or U377 (N_377,N_122,N_327);
or U378 (N_378,In_54,N_325);
nand U379 (N_379,N_148,In_285);
xnor U380 (N_380,In_173,N_240);
xor U381 (N_381,N_215,In_254);
nor U382 (N_382,N_339,In_188);
or U383 (N_383,N_265,N_340);
xor U384 (N_384,In_205,N_300);
and U385 (N_385,N_308,In_159);
nand U386 (N_386,N_293,N_303);
nor U387 (N_387,N_321,In_2);
and U388 (N_388,N_291,N_139);
or U389 (N_389,In_208,N_343);
xnor U390 (N_390,In_171,N_342);
xnor U391 (N_391,N_330,N_244);
nor U392 (N_392,N_253,In_246);
xnor U393 (N_393,N_316,In_42);
nand U394 (N_394,In_363,N_126);
xor U395 (N_395,In_89,In_134);
and U396 (N_396,N_346,In_163);
or U397 (N_397,N_310,N_302);
xor U398 (N_398,N_102,N_334);
and U399 (N_399,N_338,In_16);
or U400 (N_400,In_15,N_362);
xnor U401 (N_401,N_96,N_315);
xor U402 (N_402,In_223,In_275);
nand U403 (N_403,N_384,N_226);
and U404 (N_404,N_211,N_306);
xor U405 (N_405,N_349,N_288);
or U406 (N_406,In_416,In_222);
nand U407 (N_407,N_350,N_389);
or U408 (N_408,N_368,N_371);
or U409 (N_409,N_335,N_348);
xnor U410 (N_410,N_311,N_331);
nand U411 (N_411,N_355,N_332);
xor U412 (N_412,N_387,N_363);
or U413 (N_413,N_278,N_121);
xnor U414 (N_414,N_259,N_353);
or U415 (N_415,N_390,N_320);
xor U416 (N_416,N_385,N_361);
nand U417 (N_417,N_396,N_66);
nor U418 (N_418,N_369,N_394);
and U419 (N_419,N_395,N_382);
and U420 (N_420,N_203,N_301);
and U421 (N_421,In_245,N_356);
nand U422 (N_422,In_490,N_357);
nor U423 (N_423,N_386,N_354);
and U424 (N_424,N_366,N_324);
xnor U425 (N_425,N_73,N_364);
or U426 (N_426,N_373,N_235);
or U427 (N_427,N_254,N_280);
and U428 (N_428,N_359,N_358);
xor U429 (N_429,N_69,N_374);
and U430 (N_430,N_345,N_365);
nor U431 (N_431,N_383,N_351);
nand U432 (N_432,N_275,In_318);
nor U433 (N_433,N_273,N_252);
nand U434 (N_434,N_319,N_399);
nand U435 (N_435,N_372,N_304);
nor U436 (N_436,N_392,N_378);
xnor U437 (N_437,N_367,N_397);
and U438 (N_438,N_352,N_380);
nor U439 (N_439,N_305,N_381);
xor U440 (N_440,N_375,N_60);
nand U441 (N_441,N_314,N_360);
and U442 (N_442,N_370,N_398);
nand U443 (N_443,N_326,N_376);
xnor U444 (N_444,N_53,N_151);
or U445 (N_445,N_277,N_393);
or U446 (N_446,N_388,N_101);
xnor U447 (N_447,N_187,N_379);
and U448 (N_448,N_377,N_285);
and U449 (N_449,N_77,N_391);
or U450 (N_450,N_443,N_421);
or U451 (N_451,N_403,N_442);
nor U452 (N_452,N_446,N_412);
xor U453 (N_453,N_433,N_447);
nand U454 (N_454,N_423,N_405);
xor U455 (N_455,N_411,N_425);
or U456 (N_456,N_400,N_424);
nor U457 (N_457,N_407,N_436);
or U458 (N_458,N_435,N_408);
nor U459 (N_459,N_416,N_429);
and U460 (N_460,N_441,N_437);
xor U461 (N_461,N_445,N_402);
and U462 (N_462,N_427,N_413);
nor U463 (N_463,N_414,N_419);
or U464 (N_464,N_449,N_418);
nor U465 (N_465,N_420,N_422);
or U466 (N_466,N_409,N_434);
or U467 (N_467,N_430,N_426);
xor U468 (N_468,N_444,N_417);
or U469 (N_469,N_415,N_410);
nor U470 (N_470,N_432,N_404);
xnor U471 (N_471,N_401,N_438);
and U472 (N_472,N_428,N_448);
nand U473 (N_473,N_406,N_431);
nand U474 (N_474,N_440,N_439);
or U475 (N_475,N_447,N_445);
nand U476 (N_476,N_435,N_422);
nor U477 (N_477,N_437,N_411);
nand U478 (N_478,N_435,N_421);
xnor U479 (N_479,N_412,N_436);
or U480 (N_480,N_412,N_425);
or U481 (N_481,N_427,N_423);
xor U482 (N_482,N_411,N_447);
or U483 (N_483,N_449,N_406);
and U484 (N_484,N_420,N_426);
nand U485 (N_485,N_400,N_446);
or U486 (N_486,N_429,N_407);
nor U487 (N_487,N_402,N_443);
or U488 (N_488,N_432,N_411);
or U489 (N_489,N_406,N_421);
nor U490 (N_490,N_430,N_424);
nor U491 (N_491,N_424,N_407);
and U492 (N_492,N_446,N_411);
xnor U493 (N_493,N_415,N_449);
or U494 (N_494,N_421,N_415);
nor U495 (N_495,N_400,N_441);
and U496 (N_496,N_407,N_414);
nand U497 (N_497,N_449,N_447);
xnor U498 (N_498,N_432,N_425);
nor U499 (N_499,N_403,N_443);
or U500 (N_500,N_483,N_456);
and U501 (N_501,N_455,N_479);
and U502 (N_502,N_485,N_465);
xnor U503 (N_503,N_487,N_469);
nor U504 (N_504,N_488,N_494);
and U505 (N_505,N_463,N_477);
or U506 (N_506,N_478,N_460);
and U507 (N_507,N_473,N_492);
nand U508 (N_508,N_474,N_450);
xor U509 (N_509,N_495,N_464);
nor U510 (N_510,N_475,N_458);
and U511 (N_511,N_471,N_467);
xnor U512 (N_512,N_454,N_470);
xnor U513 (N_513,N_451,N_498);
nor U514 (N_514,N_466,N_468);
or U515 (N_515,N_459,N_462);
xor U516 (N_516,N_493,N_481);
nor U517 (N_517,N_497,N_489);
nand U518 (N_518,N_480,N_486);
and U519 (N_519,N_476,N_452);
xnor U520 (N_520,N_490,N_484);
nand U521 (N_521,N_491,N_457);
nand U522 (N_522,N_453,N_499);
and U523 (N_523,N_472,N_461);
nand U524 (N_524,N_482,N_496);
xor U525 (N_525,N_485,N_493);
nand U526 (N_526,N_466,N_465);
or U527 (N_527,N_475,N_457);
and U528 (N_528,N_480,N_495);
nor U529 (N_529,N_493,N_478);
or U530 (N_530,N_463,N_480);
nand U531 (N_531,N_454,N_484);
and U532 (N_532,N_471,N_495);
nor U533 (N_533,N_451,N_462);
nand U534 (N_534,N_468,N_465);
xor U535 (N_535,N_492,N_477);
xor U536 (N_536,N_454,N_476);
xnor U537 (N_537,N_451,N_491);
nor U538 (N_538,N_477,N_473);
xor U539 (N_539,N_485,N_464);
nand U540 (N_540,N_473,N_475);
or U541 (N_541,N_468,N_486);
and U542 (N_542,N_474,N_457);
xor U543 (N_543,N_464,N_490);
nor U544 (N_544,N_471,N_484);
or U545 (N_545,N_463,N_460);
and U546 (N_546,N_459,N_450);
nand U547 (N_547,N_497,N_486);
xor U548 (N_548,N_453,N_464);
and U549 (N_549,N_472,N_489);
nor U550 (N_550,N_521,N_546);
or U551 (N_551,N_543,N_538);
and U552 (N_552,N_501,N_503);
nand U553 (N_553,N_545,N_532);
or U554 (N_554,N_518,N_502);
nor U555 (N_555,N_504,N_515);
nand U556 (N_556,N_530,N_500);
nor U557 (N_557,N_513,N_549);
nand U558 (N_558,N_508,N_547);
nor U559 (N_559,N_539,N_548);
nand U560 (N_560,N_528,N_510);
nand U561 (N_561,N_511,N_512);
xnor U562 (N_562,N_540,N_535);
nor U563 (N_563,N_542,N_523);
and U564 (N_564,N_533,N_536);
or U565 (N_565,N_541,N_516);
nor U566 (N_566,N_529,N_527);
or U567 (N_567,N_506,N_505);
or U568 (N_568,N_509,N_519);
and U569 (N_569,N_537,N_531);
nor U570 (N_570,N_534,N_507);
or U571 (N_571,N_526,N_514);
and U572 (N_572,N_520,N_517);
or U573 (N_573,N_522,N_525);
or U574 (N_574,N_524,N_544);
nor U575 (N_575,N_508,N_509);
nor U576 (N_576,N_536,N_526);
nand U577 (N_577,N_545,N_537);
or U578 (N_578,N_536,N_545);
or U579 (N_579,N_502,N_531);
xor U580 (N_580,N_508,N_516);
nor U581 (N_581,N_516,N_501);
nor U582 (N_582,N_533,N_543);
nor U583 (N_583,N_517,N_543);
or U584 (N_584,N_529,N_531);
xor U585 (N_585,N_547,N_500);
nand U586 (N_586,N_542,N_538);
nor U587 (N_587,N_520,N_518);
or U588 (N_588,N_549,N_515);
and U589 (N_589,N_506,N_523);
nand U590 (N_590,N_522,N_501);
and U591 (N_591,N_533,N_534);
and U592 (N_592,N_530,N_548);
or U593 (N_593,N_501,N_504);
and U594 (N_594,N_544,N_537);
and U595 (N_595,N_509,N_502);
nand U596 (N_596,N_529,N_501);
and U597 (N_597,N_520,N_539);
and U598 (N_598,N_514,N_508);
and U599 (N_599,N_500,N_543);
nand U600 (N_600,N_565,N_596);
or U601 (N_601,N_586,N_578);
nor U602 (N_602,N_572,N_598);
nand U603 (N_603,N_568,N_550);
nand U604 (N_604,N_571,N_567);
nor U605 (N_605,N_594,N_551);
xnor U606 (N_606,N_580,N_584);
nand U607 (N_607,N_561,N_570);
nand U608 (N_608,N_559,N_597);
nor U609 (N_609,N_573,N_556);
and U610 (N_610,N_569,N_564);
and U611 (N_611,N_591,N_555);
or U612 (N_612,N_579,N_566);
nor U613 (N_613,N_552,N_588);
nor U614 (N_614,N_585,N_593);
nor U615 (N_615,N_595,N_587);
xor U616 (N_616,N_563,N_558);
nor U617 (N_617,N_560,N_592);
or U618 (N_618,N_577,N_557);
xor U619 (N_619,N_590,N_581);
xnor U620 (N_620,N_553,N_574);
nor U621 (N_621,N_562,N_599);
and U622 (N_622,N_576,N_582);
or U623 (N_623,N_589,N_583);
and U624 (N_624,N_554,N_575);
xnor U625 (N_625,N_575,N_561);
and U626 (N_626,N_576,N_568);
or U627 (N_627,N_597,N_596);
nor U628 (N_628,N_554,N_579);
xnor U629 (N_629,N_576,N_569);
nor U630 (N_630,N_578,N_552);
xor U631 (N_631,N_586,N_595);
nor U632 (N_632,N_596,N_595);
and U633 (N_633,N_597,N_598);
nand U634 (N_634,N_569,N_584);
nor U635 (N_635,N_567,N_563);
nor U636 (N_636,N_571,N_584);
and U637 (N_637,N_582,N_564);
nor U638 (N_638,N_550,N_570);
nor U639 (N_639,N_557,N_550);
xor U640 (N_640,N_599,N_576);
nand U641 (N_641,N_560,N_567);
nand U642 (N_642,N_587,N_561);
and U643 (N_643,N_556,N_594);
nand U644 (N_644,N_580,N_570);
nand U645 (N_645,N_582,N_583);
or U646 (N_646,N_567,N_590);
nor U647 (N_647,N_553,N_581);
nand U648 (N_648,N_561,N_581);
or U649 (N_649,N_552,N_590);
and U650 (N_650,N_620,N_648);
and U651 (N_651,N_637,N_621);
nand U652 (N_652,N_601,N_638);
and U653 (N_653,N_639,N_615);
nor U654 (N_654,N_635,N_636);
xor U655 (N_655,N_600,N_611);
or U656 (N_656,N_641,N_645);
nand U657 (N_657,N_628,N_629);
and U658 (N_658,N_610,N_646);
xnor U659 (N_659,N_607,N_619);
xor U660 (N_660,N_647,N_644);
and U661 (N_661,N_618,N_613);
and U662 (N_662,N_632,N_631);
and U663 (N_663,N_627,N_623);
nand U664 (N_664,N_633,N_625);
xnor U665 (N_665,N_617,N_606);
or U666 (N_666,N_624,N_608);
and U667 (N_667,N_616,N_609);
or U668 (N_668,N_643,N_614);
xor U669 (N_669,N_626,N_605);
xnor U670 (N_670,N_622,N_604);
nand U671 (N_671,N_602,N_649);
and U672 (N_672,N_612,N_640);
or U673 (N_673,N_630,N_642);
xnor U674 (N_674,N_603,N_634);
or U675 (N_675,N_630,N_617);
nand U676 (N_676,N_640,N_645);
or U677 (N_677,N_642,N_627);
or U678 (N_678,N_648,N_643);
nand U679 (N_679,N_631,N_649);
or U680 (N_680,N_607,N_649);
xnor U681 (N_681,N_637,N_618);
xor U682 (N_682,N_611,N_628);
nor U683 (N_683,N_645,N_615);
nand U684 (N_684,N_621,N_615);
xor U685 (N_685,N_600,N_610);
nand U686 (N_686,N_647,N_629);
nor U687 (N_687,N_647,N_626);
nor U688 (N_688,N_634,N_627);
nand U689 (N_689,N_619,N_605);
or U690 (N_690,N_646,N_608);
xnor U691 (N_691,N_644,N_616);
or U692 (N_692,N_618,N_632);
or U693 (N_693,N_608,N_619);
and U694 (N_694,N_620,N_631);
and U695 (N_695,N_639,N_636);
or U696 (N_696,N_635,N_603);
nor U697 (N_697,N_619,N_643);
and U698 (N_698,N_648,N_630);
and U699 (N_699,N_630,N_606);
or U700 (N_700,N_696,N_652);
xnor U701 (N_701,N_663,N_661);
or U702 (N_702,N_678,N_670);
nor U703 (N_703,N_680,N_658);
nand U704 (N_704,N_651,N_699);
and U705 (N_705,N_650,N_677);
nor U706 (N_706,N_665,N_659);
and U707 (N_707,N_686,N_681);
nor U708 (N_708,N_692,N_697);
nor U709 (N_709,N_657,N_683);
nand U710 (N_710,N_656,N_685);
and U711 (N_711,N_674,N_682);
xor U712 (N_712,N_698,N_655);
nand U713 (N_713,N_653,N_666);
and U714 (N_714,N_679,N_684);
and U715 (N_715,N_675,N_654);
nand U716 (N_716,N_691,N_673);
nand U717 (N_717,N_695,N_688);
xor U718 (N_718,N_668,N_689);
xor U719 (N_719,N_687,N_664);
nand U720 (N_720,N_667,N_690);
nor U721 (N_721,N_671,N_694);
nand U722 (N_722,N_672,N_669);
or U723 (N_723,N_693,N_676);
nor U724 (N_724,N_660,N_662);
xor U725 (N_725,N_659,N_690);
xnor U726 (N_726,N_697,N_656);
or U727 (N_727,N_654,N_670);
xnor U728 (N_728,N_667,N_678);
xnor U729 (N_729,N_652,N_666);
xor U730 (N_730,N_680,N_691);
and U731 (N_731,N_692,N_650);
nand U732 (N_732,N_698,N_657);
nor U733 (N_733,N_653,N_668);
and U734 (N_734,N_669,N_683);
or U735 (N_735,N_679,N_676);
nand U736 (N_736,N_653,N_651);
or U737 (N_737,N_698,N_690);
xnor U738 (N_738,N_669,N_662);
nor U739 (N_739,N_690,N_650);
nand U740 (N_740,N_677,N_694);
and U741 (N_741,N_690,N_678);
or U742 (N_742,N_678,N_657);
and U743 (N_743,N_662,N_683);
nor U744 (N_744,N_655,N_680);
or U745 (N_745,N_662,N_693);
or U746 (N_746,N_682,N_664);
nand U747 (N_747,N_693,N_681);
xnor U748 (N_748,N_679,N_667);
xor U749 (N_749,N_698,N_695);
nor U750 (N_750,N_742,N_717);
xor U751 (N_751,N_746,N_745);
and U752 (N_752,N_728,N_738);
nand U753 (N_753,N_747,N_722);
nor U754 (N_754,N_741,N_739);
xnor U755 (N_755,N_749,N_735);
nand U756 (N_756,N_740,N_707);
or U757 (N_757,N_726,N_748);
xor U758 (N_758,N_714,N_743);
xnor U759 (N_759,N_711,N_701);
or U760 (N_760,N_709,N_704);
or U761 (N_761,N_718,N_702);
or U762 (N_762,N_725,N_719);
nor U763 (N_763,N_734,N_744);
nand U764 (N_764,N_703,N_731);
nand U765 (N_765,N_723,N_732);
and U766 (N_766,N_713,N_705);
or U767 (N_767,N_710,N_712);
xor U768 (N_768,N_708,N_706);
and U769 (N_769,N_720,N_737);
or U770 (N_770,N_715,N_721);
nor U771 (N_771,N_700,N_724);
xnor U772 (N_772,N_729,N_736);
or U773 (N_773,N_727,N_730);
and U774 (N_774,N_716,N_733);
nor U775 (N_775,N_715,N_710);
or U776 (N_776,N_728,N_701);
nor U777 (N_777,N_727,N_713);
nand U778 (N_778,N_748,N_715);
xnor U779 (N_779,N_724,N_709);
nand U780 (N_780,N_714,N_721);
or U781 (N_781,N_707,N_702);
or U782 (N_782,N_737,N_719);
and U783 (N_783,N_712,N_714);
nand U784 (N_784,N_739,N_737);
nor U785 (N_785,N_744,N_716);
nand U786 (N_786,N_709,N_705);
nand U787 (N_787,N_742,N_740);
or U788 (N_788,N_733,N_712);
nand U789 (N_789,N_709,N_721);
or U790 (N_790,N_731,N_706);
and U791 (N_791,N_716,N_707);
nor U792 (N_792,N_745,N_700);
or U793 (N_793,N_715,N_702);
nor U794 (N_794,N_737,N_724);
or U795 (N_795,N_702,N_726);
or U796 (N_796,N_715,N_701);
nor U797 (N_797,N_722,N_745);
xnor U798 (N_798,N_713,N_707);
and U799 (N_799,N_706,N_742);
or U800 (N_800,N_753,N_764);
and U801 (N_801,N_773,N_785);
nor U802 (N_802,N_755,N_771);
and U803 (N_803,N_770,N_784);
nand U804 (N_804,N_761,N_766);
nor U805 (N_805,N_786,N_776);
or U806 (N_806,N_798,N_769);
and U807 (N_807,N_774,N_762);
and U808 (N_808,N_772,N_758);
or U809 (N_809,N_781,N_754);
and U810 (N_810,N_794,N_789);
or U811 (N_811,N_778,N_795);
and U812 (N_812,N_779,N_780);
and U813 (N_813,N_756,N_775);
or U814 (N_814,N_782,N_783);
nand U815 (N_815,N_757,N_790);
nand U816 (N_816,N_767,N_793);
nand U817 (N_817,N_751,N_792);
or U818 (N_818,N_750,N_791);
xnor U819 (N_819,N_787,N_759);
nand U820 (N_820,N_763,N_765);
nand U821 (N_821,N_797,N_768);
or U822 (N_822,N_788,N_777);
xnor U823 (N_823,N_752,N_799);
or U824 (N_824,N_760,N_796);
xnor U825 (N_825,N_771,N_775);
and U826 (N_826,N_765,N_797);
nor U827 (N_827,N_782,N_785);
xor U828 (N_828,N_777,N_774);
or U829 (N_829,N_761,N_793);
or U830 (N_830,N_779,N_751);
xnor U831 (N_831,N_794,N_752);
nor U832 (N_832,N_791,N_772);
nor U833 (N_833,N_772,N_760);
nor U834 (N_834,N_757,N_797);
nor U835 (N_835,N_773,N_790);
xnor U836 (N_836,N_755,N_784);
and U837 (N_837,N_750,N_786);
xnor U838 (N_838,N_785,N_765);
and U839 (N_839,N_780,N_778);
and U840 (N_840,N_761,N_780);
or U841 (N_841,N_776,N_775);
and U842 (N_842,N_775,N_772);
or U843 (N_843,N_776,N_764);
and U844 (N_844,N_771,N_776);
nor U845 (N_845,N_769,N_764);
nor U846 (N_846,N_797,N_798);
and U847 (N_847,N_788,N_753);
or U848 (N_848,N_775,N_788);
or U849 (N_849,N_758,N_779);
or U850 (N_850,N_809,N_826);
xor U851 (N_851,N_835,N_807);
nand U852 (N_852,N_811,N_830);
nor U853 (N_853,N_847,N_805);
nand U854 (N_854,N_819,N_829);
nand U855 (N_855,N_832,N_848);
nor U856 (N_856,N_803,N_817);
xor U857 (N_857,N_846,N_831);
or U858 (N_858,N_849,N_838);
nand U859 (N_859,N_816,N_800);
nand U860 (N_860,N_837,N_808);
xnor U861 (N_861,N_842,N_825);
or U862 (N_862,N_841,N_828);
nor U863 (N_863,N_812,N_810);
nand U864 (N_864,N_802,N_844);
xnor U865 (N_865,N_815,N_821);
xnor U866 (N_866,N_827,N_820);
nor U867 (N_867,N_801,N_814);
nor U868 (N_868,N_836,N_839);
and U869 (N_869,N_804,N_813);
or U870 (N_870,N_845,N_822);
and U871 (N_871,N_823,N_843);
nand U872 (N_872,N_840,N_834);
nand U873 (N_873,N_818,N_824);
or U874 (N_874,N_806,N_833);
nor U875 (N_875,N_849,N_840);
or U876 (N_876,N_800,N_843);
nand U877 (N_877,N_826,N_832);
nor U878 (N_878,N_806,N_848);
nor U879 (N_879,N_808,N_829);
nor U880 (N_880,N_821,N_822);
xor U881 (N_881,N_814,N_804);
nor U882 (N_882,N_824,N_842);
or U883 (N_883,N_822,N_806);
nand U884 (N_884,N_833,N_828);
and U885 (N_885,N_819,N_821);
xor U886 (N_886,N_822,N_805);
nor U887 (N_887,N_849,N_841);
nand U888 (N_888,N_802,N_823);
nor U889 (N_889,N_819,N_818);
nand U890 (N_890,N_846,N_803);
or U891 (N_891,N_823,N_831);
nand U892 (N_892,N_826,N_831);
and U893 (N_893,N_803,N_811);
and U894 (N_894,N_801,N_849);
or U895 (N_895,N_823,N_826);
nor U896 (N_896,N_846,N_844);
and U897 (N_897,N_824,N_802);
nor U898 (N_898,N_833,N_848);
nand U899 (N_899,N_815,N_847);
or U900 (N_900,N_861,N_856);
or U901 (N_901,N_860,N_878);
and U902 (N_902,N_872,N_851);
xor U903 (N_903,N_873,N_852);
xor U904 (N_904,N_870,N_897);
xnor U905 (N_905,N_893,N_865);
and U906 (N_906,N_862,N_894);
nand U907 (N_907,N_855,N_881);
or U908 (N_908,N_876,N_884);
nand U909 (N_909,N_880,N_875);
and U910 (N_910,N_890,N_863);
nand U911 (N_911,N_899,N_891);
xnor U912 (N_912,N_871,N_874);
nor U913 (N_913,N_858,N_857);
xnor U914 (N_914,N_859,N_877);
or U915 (N_915,N_889,N_886);
nor U916 (N_916,N_892,N_868);
xnor U917 (N_917,N_885,N_895);
or U918 (N_918,N_869,N_883);
nor U919 (N_919,N_887,N_850);
and U920 (N_920,N_867,N_853);
xnor U921 (N_921,N_864,N_854);
xnor U922 (N_922,N_888,N_896);
nor U923 (N_923,N_866,N_898);
or U924 (N_924,N_879,N_882);
xor U925 (N_925,N_884,N_881);
and U926 (N_926,N_884,N_861);
or U927 (N_927,N_887,N_886);
nand U928 (N_928,N_890,N_894);
nor U929 (N_929,N_894,N_888);
and U930 (N_930,N_856,N_897);
or U931 (N_931,N_868,N_889);
or U932 (N_932,N_859,N_882);
nor U933 (N_933,N_891,N_851);
xnor U934 (N_934,N_857,N_865);
or U935 (N_935,N_862,N_860);
and U936 (N_936,N_888,N_886);
or U937 (N_937,N_850,N_858);
or U938 (N_938,N_883,N_870);
or U939 (N_939,N_887,N_881);
and U940 (N_940,N_890,N_886);
xnor U941 (N_941,N_894,N_876);
and U942 (N_942,N_858,N_864);
nor U943 (N_943,N_861,N_875);
nor U944 (N_944,N_874,N_895);
nor U945 (N_945,N_897,N_865);
or U946 (N_946,N_897,N_867);
or U947 (N_947,N_893,N_866);
nor U948 (N_948,N_867,N_858);
nand U949 (N_949,N_855,N_894);
or U950 (N_950,N_909,N_948);
and U951 (N_951,N_933,N_913);
nand U952 (N_952,N_905,N_946);
nor U953 (N_953,N_920,N_947);
nand U954 (N_954,N_907,N_900);
xnor U955 (N_955,N_904,N_937);
xnor U956 (N_956,N_914,N_919);
nor U957 (N_957,N_936,N_922);
nand U958 (N_958,N_911,N_910);
and U959 (N_959,N_925,N_942);
nand U960 (N_960,N_912,N_926);
nor U961 (N_961,N_934,N_916);
nor U962 (N_962,N_903,N_929);
nor U963 (N_963,N_923,N_906);
nor U964 (N_964,N_930,N_917);
nand U965 (N_965,N_939,N_949);
xnor U966 (N_966,N_943,N_908);
and U967 (N_967,N_931,N_945);
nor U968 (N_968,N_940,N_938);
or U969 (N_969,N_924,N_944);
nor U970 (N_970,N_928,N_927);
nor U971 (N_971,N_935,N_941);
or U972 (N_972,N_902,N_915);
nor U973 (N_973,N_932,N_921);
xnor U974 (N_974,N_901,N_918);
or U975 (N_975,N_929,N_925);
or U976 (N_976,N_949,N_930);
or U977 (N_977,N_907,N_927);
nand U978 (N_978,N_915,N_943);
and U979 (N_979,N_908,N_941);
nor U980 (N_980,N_926,N_931);
nor U981 (N_981,N_934,N_929);
or U982 (N_982,N_940,N_904);
xnor U983 (N_983,N_939,N_932);
nand U984 (N_984,N_908,N_902);
and U985 (N_985,N_917,N_922);
or U986 (N_986,N_927,N_938);
nor U987 (N_987,N_924,N_934);
nor U988 (N_988,N_931,N_912);
nor U989 (N_989,N_922,N_932);
or U990 (N_990,N_917,N_924);
nor U991 (N_991,N_906,N_907);
nand U992 (N_992,N_948,N_934);
nand U993 (N_993,N_905,N_927);
nor U994 (N_994,N_910,N_909);
xor U995 (N_995,N_920,N_932);
and U996 (N_996,N_908,N_940);
and U997 (N_997,N_939,N_947);
xor U998 (N_998,N_913,N_916);
and U999 (N_999,N_909,N_913);
or U1000 (N_1000,N_988,N_985);
and U1001 (N_1001,N_981,N_986);
xnor U1002 (N_1002,N_987,N_974);
nor U1003 (N_1003,N_982,N_993);
nand U1004 (N_1004,N_965,N_967);
and U1005 (N_1005,N_956,N_971);
and U1006 (N_1006,N_963,N_961);
and U1007 (N_1007,N_951,N_970);
or U1008 (N_1008,N_990,N_962);
nand U1009 (N_1009,N_999,N_973);
nand U1010 (N_1010,N_955,N_998);
and U1011 (N_1011,N_972,N_954);
and U1012 (N_1012,N_968,N_979);
nor U1013 (N_1013,N_959,N_957);
nor U1014 (N_1014,N_976,N_989);
nand U1015 (N_1015,N_980,N_969);
or U1016 (N_1016,N_958,N_994);
and U1017 (N_1017,N_997,N_983);
and U1018 (N_1018,N_975,N_996);
xnor U1019 (N_1019,N_966,N_984);
nor U1020 (N_1020,N_952,N_950);
and U1021 (N_1021,N_960,N_992);
and U1022 (N_1022,N_991,N_953);
nand U1023 (N_1023,N_995,N_977);
and U1024 (N_1024,N_964,N_978);
xnor U1025 (N_1025,N_984,N_962);
xnor U1026 (N_1026,N_993,N_966);
and U1027 (N_1027,N_969,N_978);
nor U1028 (N_1028,N_987,N_986);
xor U1029 (N_1029,N_978,N_961);
xnor U1030 (N_1030,N_982,N_973);
xor U1031 (N_1031,N_992,N_951);
nand U1032 (N_1032,N_969,N_997);
xor U1033 (N_1033,N_997,N_957);
nor U1034 (N_1034,N_975,N_962);
and U1035 (N_1035,N_967,N_962);
xor U1036 (N_1036,N_951,N_954);
and U1037 (N_1037,N_976,N_963);
xor U1038 (N_1038,N_999,N_952);
xnor U1039 (N_1039,N_953,N_983);
nor U1040 (N_1040,N_997,N_968);
or U1041 (N_1041,N_961,N_960);
or U1042 (N_1042,N_954,N_959);
and U1043 (N_1043,N_954,N_998);
nor U1044 (N_1044,N_954,N_963);
xor U1045 (N_1045,N_980,N_989);
xor U1046 (N_1046,N_978,N_997);
and U1047 (N_1047,N_966,N_961);
and U1048 (N_1048,N_968,N_976);
xnor U1049 (N_1049,N_956,N_986);
nand U1050 (N_1050,N_1039,N_1033);
nor U1051 (N_1051,N_1030,N_1048);
xor U1052 (N_1052,N_1043,N_1000);
and U1053 (N_1053,N_1013,N_1004);
nand U1054 (N_1054,N_1027,N_1010);
nand U1055 (N_1055,N_1008,N_1035);
nand U1056 (N_1056,N_1003,N_1037);
nand U1057 (N_1057,N_1022,N_1042);
and U1058 (N_1058,N_1024,N_1005);
or U1059 (N_1059,N_1028,N_1040);
xnor U1060 (N_1060,N_1045,N_1007);
xor U1061 (N_1061,N_1046,N_1009);
xor U1062 (N_1062,N_1014,N_1019);
nand U1063 (N_1063,N_1034,N_1018);
nand U1064 (N_1064,N_1029,N_1049);
xnor U1065 (N_1065,N_1047,N_1002);
nand U1066 (N_1066,N_1015,N_1017);
nor U1067 (N_1067,N_1023,N_1031);
nor U1068 (N_1068,N_1026,N_1036);
or U1069 (N_1069,N_1041,N_1006);
nor U1070 (N_1070,N_1011,N_1038);
xnor U1071 (N_1071,N_1044,N_1001);
and U1072 (N_1072,N_1032,N_1025);
nor U1073 (N_1073,N_1020,N_1021);
or U1074 (N_1074,N_1016,N_1012);
nand U1075 (N_1075,N_1024,N_1000);
nor U1076 (N_1076,N_1006,N_1044);
nor U1077 (N_1077,N_1004,N_1026);
xor U1078 (N_1078,N_1042,N_1025);
nand U1079 (N_1079,N_1009,N_1008);
xnor U1080 (N_1080,N_1020,N_1011);
nand U1081 (N_1081,N_1004,N_1037);
nand U1082 (N_1082,N_1028,N_1004);
and U1083 (N_1083,N_1019,N_1049);
nand U1084 (N_1084,N_1032,N_1026);
and U1085 (N_1085,N_1036,N_1018);
or U1086 (N_1086,N_1017,N_1044);
and U1087 (N_1087,N_1003,N_1047);
and U1088 (N_1088,N_1012,N_1021);
or U1089 (N_1089,N_1049,N_1008);
nor U1090 (N_1090,N_1004,N_1015);
nor U1091 (N_1091,N_1048,N_1040);
or U1092 (N_1092,N_1025,N_1012);
nor U1093 (N_1093,N_1024,N_1017);
and U1094 (N_1094,N_1044,N_1008);
and U1095 (N_1095,N_1027,N_1015);
nand U1096 (N_1096,N_1023,N_1039);
nand U1097 (N_1097,N_1006,N_1037);
nand U1098 (N_1098,N_1017,N_1022);
xnor U1099 (N_1099,N_1034,N_1008);
nor U1100 (N_1100,N_1067,N_1079);
nand U1101 (N_1101,N_1090,N_1092);
nor U1102 (N_1102,N_1064,N_1056);
or U1103 (N_1103,N_1053,N_1088);
nand U1104 (N_1104,N_1097,N_1096);
or U1105 (N_1105,N_1061,N_1069);
or U1106 (N_1106,N_1052,N_1055);
xnor U1107 (N_1107,N_1060,N_1082);
nand U1108 (N_1108,N_1099,N_1072);
nand U1109 (N_1109,N_1095,N_1068);
and U1110 (N_1110,N_1065,N_1084);
nor U1111 (N_1111,N_1091,N_1080);
nor U1112 (N_1112,N_1071,N_1062);
nand U1113 (N_1113,N_1058,N_1086);
nor U1114 (N_1114,N_1057,N_1051);
and U1115 (N_1115,N_1085,N_1098);
and U1116 (N_1116,N_1066,N_1059);
nand U1117 (N_1117,N_1054,N_1087);
and U1118 (N_1118,N_1063,N_1074);
or U1119 (N_1119,N_1081,N_1094);
nor U1120 (N_1120,N_1073,N_1050);
nor U1121 (N_1121,N_1070,N_1093);
nand U1122 (N_1122,N_1076,N_1078);
and U1123 (N_1123,N_1089,N_1075);
nand U1124 (N_1124,N_1077,N_1083);
and U1125 (N_1125,N_1096,N_1071);
or U1126 (N_1126,N_1081,N_1079);
or U1127 (N_1127,N_1075,N_1062);
and U1128 (N_1128,N_1077,N_1068);
nand U1129 (N_1129,N_1062,N_1088);
and U1130 (N_1130,N_1050,N_1060);
and U1131 (N_1131,N_1083,N_1055);
or U1132 (N_1132,N_1089,N_1055);
or U1133 (N_1133,N_1076,N_1063);
or U1134 (N_1134,N_1069,N_1064);
or U1135 (N_1135,N_1060,N_1076);
nor U1136 (N_1136,N_1097,N_1084);
xor U1137 (N_1137,N_1091,N_1053);
nand U1138 (N_1138,N_1079,N_1083);
xor U1139 (N_1139,N_1085,N_1093);
or U1140 (N_1140,N_1078,N_1092);
nand U1141 (N_1141,N_1074,N_1086);
or U1142 (N_1142,N_1069,N_1080);
xnor U1143 (N_1143,N_1071,N_1075);
nand U1144 (N_1144,N_1099,N_1067);
nand U1145 (N_1145,N_1066,N_1093);
xor U1146 (N_1146,N_1089,N_1080);
nand U1147 (N_1147,N_1071,N_1088);
and U1148 (N_1148,N_1084,N_1088);
or U1149 (N_1149,N_1084,N_1062);
or U1150 (N_1150,N_1105,N_1120);
xor U1151 (N_1151,N_1116,N_1126);
and U1152 (N_1152,N_1131,N_1140);
xnor U1153 (N_1153,N_1135,N_1113);
or U1154 (N_1154,N_1117,N_1111);
nor U1155 (N_1155,N_1143,N_1118);
or U1156 (N_1156,N_1108,N_1149);
nor U1157 (N_1157,N_1130,N_1115);
nand U1158 (N_1158,N_1139,N_1132);
and U1159 (N_1159,N_1144,N_1128);
or U1160 (N_1160,N_1141,N_1134);
and U1161 (N_1161,N_1122,N_1123);
or U1162 (N_1162,N_1138,N_1104);
nor U1163 (N_1163,N_1106,N_1125);
xnor U1164 (N_1164,N_1136,N_1146);
nor U1165 (N_1165,N_1114,N_1119);
nor U1166 (N_1166,N_1103,N_1100);
or U1167 (N_1167,N_1129,N_1147);
and U1168 (N_1168,N_1124,N_1137);
xor U1169 (N_1169,N_1127,N_1101);
and U1170 (N_1170,N_1109,N_1102);
nand U1171 (N_1171,N_1133,N_1121);
or U1172 (N_1172,N_1107,N_1112);
nand U1173 (N_1173,N_1145,N_1110);
xor U1174 (N_1174,N_1148,N_1142);
nand U1175 (N_1175,N_1126,N_1104);
nand U1176 (N_1176,N_1100,N_1116);
xor U1177 (N_1177,N_1120,N_1148);
xor U1178 (N_1178,N_1101,N_1102);
xnor U1179 (N_1179,N_1128,N_1108);
nor U1180 (N_1180,N_1103,N_1146);
nand U1181 (N_1181,N_1112,N_1146);
xnor U1182 (N_1182,N_1102,N_1130);
and U1183 (N_1183,N_1137,N_1145);
xor U1184 (N_1184,N_1119,N_1127);
nor U1185 (N_1185,N_1103,N_1106);
nor U1186 (N_1186,N_1107,N_1139);
xor U1187 (N_1187,N_1124,N_1144);
nand U1188 (N_1188,N_1118,N_1111);
nor U1189 (N_1189,N_1117,N_1107);
or U1190 (N_1190,N_1147,N_1136);
and U1191 (N_1191,N_1136,N_1131);
or U1192 (N_1192,N_1112,N_1120);
nand U1193 (N_1193,N_1132,N_1135);
or U1194 (N_1194,N_1125,N_1113);
and U1195 (N_1195,N_1114,N_1123);
nor U1196 (N_1196,N_1110,N_1133);
xor U1197 (N_1197,N_1114,N_1104);
or U1198 (N_1198,N_1141,N_1136);
and U1199 (N_1199,N_1120,N_1126);
nand U1200 (N_1200,N_1179,N_1192);
or U1201 (N_1201,N_1177,N_1185);
or U1202 (N_1202,N_1159,N_1152);
or U1203 (N_1203,N_1194,N_1154);
nor U1204 (N_1204,N_1164,N_1163);
xor U1205 (N_1205,N_1161,N_1174);
xnor U1206 (N_1206,N_1189,N_1196);
nand U1207 (N_1207,N_1190,N_1187);
or U1208 (N_1208,N_1198,N_1184);
nand U1209 (N_1209,N_1180,N_1170);
and U1210 (N_1210,N_1168,N_1181);
nor U1211 (N_1211,N_1166,N_1157);
xor U1212 (N_1212,N_1167,N_1175);
and U1213 (N_1213,N_1199,N_1195);
and U1214 (N_1214,N_1188,N_1156);
and U1215 (N_1215,N_1165,N_1178);
nor U1216 (N_1216,N_1191,N_1197);
and U1217 (N_1217,N_1182,N_1169);
xnor U1218 (N_1218,N_1160,N_1162);
and U1219 (N_1219,N_1171,N_1150);
xnor U1220 (N_1220,N_1155,N_1176);
xor U1221 (N_1221,N_1183,N_1173);
nor U1222 (N_1222,N_1158,N_1193);
xor U1223 (N_1223,N_1172,N_1186);
xor U1224 (N_1224,N_1151,N_1153);
nor U1225 (N_1225,N_1157,N_1156);
nor U1226 (N_1226,N_1188,N_1177);
nand U1227 (N_1227,N_1180,N_1181);
and U1228 (N_1228,N_1152,N_1176);
nand U1229 (N_1229,N_1184,N_1191);
xnor U1230 (N_1230,N_1192,N_1159);
or U1231 (N_1231,N_1190,N_1184);
nor U1232 (N_1232,N_1158,N_1156);
nand U1233 (N_1233,N_1181,N_1194);
xor U1234 (N_1234,N_1196,N_1172);
nor U1235 (N_1235,N_1184,N_1169);
xnor U1236 (N_1236,N_1190,N_1168);
nand U1237 (N_1237,N_1155,N_1169);
nor U1238 (N_1238,N_1181,N_1173);
nor U1239 (N_1239,N_1156,N_1189);
or U1240 (N_1240,N_1189,N_1158);
and U1241 (N_1241,N_1167,N_1194);
and U1242 (N_1242,N_1157,N_1190);
and U1243 (N_1243,N_1181,N_1172);
nand U1244 (N_1244,N_1164,N_1151);
and U1245 (N_1245,N_1198,N_1160);
xnor U1246 (N_1246,N_1198,N_1189);
xor U1247 (N_1247,N_1164,N_1154);
nor U1248 (N_1248,N_1165,N_1156);
xnor U1249 (N_1249,N_1186,N_1170);
or U1250 (N_1250,N_1243,N_1213);
nand U1251 (N_1251,N_1208,N_1230);
xor U1252 (N_1252,N_1238,N_1220);
and U1253 (N_1253,N_1216,N_1221);
nor U1254 (N_1254,N_1234,N_1210);
xnor U1255 (N_1255,N_1241,N_1217);
nand U1256 (N_1256,N_1203,N_1248);
or U1257 (N_1257,N_1209,N_1246);
xnor U1258 (N_1258,N_1247,N_1204);
nor U1259 (N_1259,N_1228,N_1202);
nor U1260 (N_1260,N_1244,N_1219);
and U1261 (N_1261,N_1235,N_1214);
nor U1262 (N_1262,N_1201,N_1242);
xor U1263 (N_1263,N_1239,N_1237);
nor U1264 (N_1264,N_1233,N_1211);
nor U1265 (N_1265,N_1229,N_1222);
or U1266 (N_1266,N_1207,N_1245);
or U1267 (N_1267,N_1249,N_1200);
nor U1268 (N_1268,N_1240,N_1227);
nor U1269 (N_1269,N_1232,N_1218);
nor U1270 (N_1270,N_1226,N_1212);
and U1271 (N_1271,N_1236,N_1205);
xnor U1272 (N_1272,N_1224,N_1215);
nor U1273 (N_1273,N_1223,N_1206);
or U1274 (N_1274,N_1231,N_1225);
nand U1275 (N_1275,N_1229,N_1204);
xor U1276 (N_1276,N_1236,N_1227);
or U1277 (N_1277,N_1202,N_1226);
xnor U1278 (N_1278,N_1208,N_1231);
and U1279 (N_1279,N_1243,N_1239);
and U1280 (N_1280,N_1204,N_1218);
or U1281 (N_1281,N_1237,N_1245);
nand U1282 (N_1282,N_1212,N_1215);
xor U1283 (N_1283,N_1230,N_1229);
and U1284 (N_1284,N_1228,N_1239);
xor U1285 (N_1285,N_1201,N_1241);
nand U1286 (N_1286,N_1205,N_1207);
and U1287 (N_1287,N_1249,N_1201);
or U1288 (N_1288,N_1227,N_1211);
and U1289 (N_1289,N_1206,N_1228);
and U1290 (N_1290,N_1243,N_1211);
nor U1291 (N_1291,N_1208,N_1237);
or U1292 (N_1292,N_1223,N_1203);
xnor U1293 (N_1293,N_1242,N_1205);
xnor U1294 (N_1294,N_1238,N_1236);
nand U1295 (N_1295,N_1236,N_1210);
xnor U1296 (N_1296,N_1231,N_1210);
nand U1297 (N_1297,N_1217,N_1224);
and U1298 (N_1298,N_1228,N_1213);
nor U1299 (N_1299,N_1226,N_1238);
and U1300 (N_1300,N_1267,N_1290);
xnor U1301 (N_1301,N_1254,N_1272);
nor U1302 (N_1302,N_1264,N_1261);
xor U1303 (N_1303,N_1262,N_1291);
or U1304 (N_1304,N_1256,N_1278);
xnor U1305 (N_1305,N_1285,N_1295);
nor U1306 (N_1306,N_1279,N_1269);
or U1307 (N_1307,N_1299,N_1266);
nor U1308 (N_1308,N_1287,N_1268);
xor U1309 (N_1309,N_1280,N_1296);
or U1310 (N_1310,N_1251,N_1271);
nand U1311 (N_1311,N_1255,N_1252);
and U1312 (N_1312,N_1253,N_1258);
and U1313 (N_1313,N_1286,N_1260);
nor U1314 (N_1314,N_1283,N_1281);
nor U1315 (N_1315,N_1259,N_1288);
nor U1316 (N_1316,N_1257,N_1263);
or U1317 (N_1317,N_1297,N_1270);
xnor U1318 (N_1318,N_1265,N_1274);
nor U1319 (N_1319,N_1289,N_1294);
nand U1320 (N_1320,N_1284,N_1273);
nand U1321 (N_1321,N_1292,N_1293);
and U1322 (N_1322,N_1250,N_1298);
and U1323 (N_1323,N_1275,N_1277);
and U1324 (N_1324,N_1276,N_1282);
nor U1325 (N_1325,N_1286,N_1263);
or U1326 (N_1326,N_1281,N_1270);
xnor U1327 (N_1327,N_1253,N_1255);
and U1328 (N_1328,N_1257,N_1273);
nand U1329 (N_1329,N_1276,N_1263);
xor U1330 (N_1330,N_1262,N_1289);
nor U1331 (N_1331,N_1280,N_1254);
and U1332 (N_1332,N_1274,N_1283);
or U1333 (N_1333,N_1293,N_1291);
and U1334 (N_1334,N_1289,N_1259);
and U1335 (N_1335,N_1275,N_1291);
and U1336 (N_1336,N_1270,N_1299);
nor U1337 (N_1337,N_1276,N_1280);
xnor U1338 (N_1338,N_1287,N_1275);
and U1339 (N_1339,N_1258,N_1269);
or U1340 (N_1340,N_1273,N_1252);
nand U1341 (N_1341,N_1287,N_1252);
and U1342 (N_1342,N_1274,N_1252);
or U1343 (N_1343,N_1284,N_1256);
nor U1344 (N_1344,N_1258,N_1264);
xnor U1345 (N_1345,N_1299,N_1272);
or U1346 (N_1346,N_1259,N_1264);
nand U1347 (N_1347,N_1260,N_1288);
nand U1348 (N_1348,N_1257,N_1267);
and U1349 (N_1349,N_1264,N_1281);
xor U1350 (N_1350,N_1314,N_1304);
nand U1351 (N_1351,N_1323,N_1306);
xor U1352 (N_1352,N_1305,N_1335);
xor U1353 (N_1353,N_1331,N_1345);
and U1354 (N_1354,N_1321,N_1346);
or U1355 (N_1355,N_1339,N_1329);
and U1356 (N_1356,N_1317,N_1332);
nand U1357 (N_1357,N_1312,N_1324);
nor U1358 (N_1358,N_1327,N_1300);
or U1359 (N_1359,N_1319,N_1307);
nor U1360 (N_1360,N_1349,N_1313);
nor U1361 (N_1361,N_1344,N_1303);
nand U1362 (N_1362,N_1310,N_1309);
xor U1363 (N_1363,N_1318,N_1315);
or U1364 (N_1364,N_1334,N_1340);
nand U1365 (N_1365,N_1326,N_1325);
nor U1366 (N_1366,N_1320,N_1348);
nand U1367 (N_1367,N_1316,N_1322);
nor U1368 (N_1368,N_1347,N_1333);
and U1369 (N_1369,N_1342,N_1341);
nor U1370 (N_1370,N_1336,N_1328);
nand U1371 (N_1371,N_1311,N_1308);
or U1372 (N_1372,N_1301,N_1330);
nand U1373 (N_1373,N_1302,N_1337);
and U1374 (N_1374,N_1343,N_1338);
nand U1375 (N_1375,N_1316,N_1302);
or U1376 (N_1376,N_1345,N_1309);
xor U1377 (N_1377,N_1343,N_1323);
nor U1378 (N_1378,N_1346,N_1306);
and U1379 (N_1379,N_1339,N_1334);
or U1380 (N_1380,N_1313,N_1342);
xor U1381 (N_1381,N_1319,N_1347);
xnor U1382 (N_1382,N_1346,N_1336);
nor U1383 (N_1383,N_1337,N_1335);
or U1384 (N_1384,N_1339,N_1349);
or U1385 (N_1385,N_1304,N_1311);
and U1386 (N_1386,N_1318,N_1303);
nor U1387 (N_1387,N_1308,N_1346);
nand U1388 (N_1388,N_1338,N_1305);
xor U1389 (N_1389,N_1306,N_1303);
and U1390 (N_1390,N_1322,N_1326);
xor U1391 (N_1391,N_1335,N_1330);
xnor U1392 (N_1392,N_1340,N_1325);
or U1393 (N_1393,N_1300,N_1306);
nand U1394 (N_1394,N_1335,N_1346);
xnor U1395 (N_1395,N_1302,N_1346);
nor U1396 (N_1396,N_1349,N_1323);
nor U1397 (N_1397,N_1324,N_1300);
and U1398 (N_1398,N_1349,N_1328);
or U1399 (N_1399,N_1314,N_1305);
nor U1400 (N_1400,N_1368,N_1376);
and U1401 (N_1401,N_1384,N_1350);
or U1402 (N_1402,N_1358,N_1390);
nand U1403 (N_1403,N_1365,N_1383);
xnor U1404 (N_1404,N_1370,N_1369);
or U1405 (N_1405,N_1373,N_1357);
xor U1406 (N_1406,N_1379,N_1378);
nor U1407 (N_1407,N_1386,N_1374);
nand U1408 (N_1408,N_1388,N_1351);
xnor U1409 (N_1409,N_1385,N_1391);
nand U1410 (N_1410,N_1364,N_1389);
nor U1411 (N_1411,N_1360,N_1381);
nand U1412 (N_1412,N_1356,N_1362);
and U1413 (N_1413,N_1392,N_1393);
nand U1414 (N_1414,N_1363,N_1375);
and U1415 (N_1415,N_1387,N_1354);
nand U1416 (N_1416,N_1353,N_1398);
xor U1417 (N_1417,N_1377,N_1397);
nor U1418 (N_1418,N_1352,N_1367);
nand U1419 (N_1419,N_1399,N_1366);
nand U1420 (N_1420,N_1394,N_1371);
nor U1421 (N_1421,N_1396,N_1355);
xnor U1422 (N_1422,N_1372,N_1395);
xnor U1423 (N_1423,N_1361,N_1382);
nor U1424 (N_1424,N_1380,N_1359);
nor U1425 (N_1425,N_1363,N_1388);
nand U1426 (N_1426,N_1392,N_1380);
nand U1427 (N_1427,N_1394,N_1356);
nand U1428 (N_1428,N_1357,N_1395);
nor U1429 (N_1429,N_1388,N_1382);
nor U1430 (N_1430,N_1360,N_1351);
or U1431 (N_1431,N_1394,N_1361);
or U1432 (N_1432,N_1396,N_1398);
nand U1433 (N_1433,N_1389,N_1397);
or U1434 (N_1434,N_1362,N_1392);
nor U1435 (N_1435,N_1370,N_1360);
nand U1436 (N_1436,N_1382,N_1368);
or U1437 (N_1437,N_1368,N_1365);
nand U1438 (N_1438,N_1390,N_1382);
and U1439 (N_1439,N_1397,N_1373);
nand U1440 (N_1440,N_1350,N_1377);
xor U1441 (N_1441,N_1382,N_1357);
or U1442 (N_1442,N_1362,N_1352);
xnor U1443 (N_1443,N_1361,N_1379);
and U1444 (N_1444,N_1376,N_1366);
nand U1445 (N_1445,N_1350,N_1397);
and U1446 (N_1446,N_1389,N_1386);
and U1447 (N_1447,N_1370,N_1352);
xor U1448 (N_1448,N_1388,N_1377);
nand U1449 (N_1449,N_1398,N_1364);
or U1450 (N_1450,N_1406,N_1423);
nor U1451 (N_1451,N_1433,N_1449);
and U1452 (N_1452,N_1413,N_1430);
xnor U1453 (N_1453,N_1422,N_1442);
nand U1454 (N_1454,N_1418,N_1437);
or U1455 (N_1455,N_1428,N_1446);
nand U1456 (N_1456,N_1403,N_1447);
xor U1457 (N_1457,N_1414,N_1436);
nor U1458 (N_1458,N_1426,N_1431);
or U1459 (N_1459,N_1432,N_1401);
xor U1460 (N_1460,N_1438,N_1408);
nand U1461 (N_1461,N_1441,N_1435);
or U1462 (N_1462,N_1444,N_1443);
and U1463 (N_1463,N_1440,N_1410);
or U1464 (N_1464,N_1411,N_1417);
xnor U1465 (N_1465,N_1421,N_1416);
nand U1466 (N_1466,N_1425,N_1420);
nand U1467 (N_1467,N_1409,N_1427);
and U1468 (N_1468,N_1402,N_1424);
nor U1469 (N_1469,N_1412,N_1448);
xor U1470 (N_1470,N_1404,N_1405);
xor U1471 (N_1471,N_1429,N_1439);
nand U1472 (N_1472,N_1419,N_1400);
and U1473 (N_1473,N_1407,N_1415);
and U1474 (N_1474,N_1445,N_1434);
nand U1475 (N_1475,N_1413,N_1425);
xor U1476 (N_1476,N_1449,N_1437);
and U1477 (N_1477,N_1413,N_1445);
and U1478 (N_1478,N_1404,N_1442);
or U1479 (N_1479,N_1446,N_1416);
nor U1480 (N_1480,N_1437,N_1412);
and U1481 (N_1481,N_1436,N_1418);
nand U1482 (N_1482,N_1431,N_1448);
and U1483 (N_1483,N_1435,N_1425);
xor U1484 (N_1484,N_1402,N_1410);
xnor U1485 (N_1485,N_1417,N_1449);
nor U1486 (N_1486,N_1440,N_1431);
or U1487 (N_1487,N_1440,N_1428);
nor U1488 (N_1488,N_1439,N_1430);
nor U1489 (N_1489,N_1406,N_1442);
xor U1490 (N_1490,N_1401,N_1443);
and U1491 (N_1491,N_1443,N_1409);
nand U1492 (N_1492,N_1442,N_1445);
nand U1493 (N_1493,N_1432,N_1439);
nor U1494 (N_1494,N_1424,N_1411);
nor U1495 (N_1495,N_1404,N_1425);
nor U1496 (N_1496,N_1449,N_1411);
or U1497 (N_1497,N_1401,N_1414);
and U1498 (N_1498,N_1423,N_1419);
or U1499 (N_1499,N_1417,N_1420);
or U1500 (N_1500,N_1497,N_1493);
and U1501 (N_1501,N_1484,N_1476);
or U1502 (N_1502,N_1468,N_1466);
xnor U1503 (N_1503,N_1460,N_1469);
xor U1504 (N_1504,N_1450,N_1459);
nor U1505 (N_1505,N_1463,N_1479);
and U1506 (N_1506,N_1451,N_1487);
nand U1507 (N_1507,N_1478,N_1494);
or U1508 (N_1508,N_1455,N_1495);
nor U1509 (N_1509,N_1470,N_1472);
nor U1510 (N_1510,N_1480,N_1488);
xor U1511 (N_1511,N_1461,N_1496);
or U1512 (N_1512,N_1498,N_1471);
and U1513 (N_1513,N_1481,N_1462);
xnor U1514 (N_1514,N_1458,N_1483);
nor U1515 (N_1515,N_1490,N_1457);
nor U1516 (N_1516,N_1492,N_1456);
nor U1517 (N_1517,N_1486,N_1489);
nand U1518 (N_1518,N_1465,N_1473);
or U1519 (N_1519,N_1452,N_1453);
nand U1520 (N_1520,N_1475,N_1485);
and U1521 (N_1521,N_1467,N_1491);
and U1522 (N_1522,N_1499,N_1482);
nand U1523 (N_1523,N_1454,N_1474);
nor U1524 (N_1524,N_1477,N_1464);
or U1525 (N_1525,N_1488,N_1475);
nor U1526 (N_1526,N_1457,N_1462);
xor U1527 (N_1527,N_1495,N_1484);
xnor U1528 (N_1528,N_1493,N_1470);
nand U1529 (N_1529,N_1482,N_1487);
or U1530 (N_1530,N_1474,N_1494);
nor U1531 (N_1531,N_1493,N_1480);
and U1532 (N_1532,N_1486,N_1460);
and U1533 (N_1533,N_1484,N_1488);
and U1534 (N_1534,N_1456,N_1474);
nand U1535 (N_1535,N_1475,N_1499);
nand U1536 (N_1536,N_1472,N_1494);
nand U1537 (N_1537,N_1456,N_1484);
xor U1538 (N_1538,N_1498,N_1451);
or U1539 (N_1539,N_1454,N_1486);
xnor U1540 (N_1540,N_1461,N_1473);
nand U1541 (N_1541,N_1455,N_1464);
or U1542 (N_1542,N_1451,N_1483);
nor U1543 (N_1543,N_1494,N_1465);
xor U1544 (N_1544,N_1455,N_1457);
xnor U1545 (N_1545,N_1461,N_1456);
nor U1546 (N_1546,N_1498,N_1462);
or U1547 (N_1547,N_1494,N_1475);
or U1548 (N_1548,N_1479,N_1496);
nand U1549 (N_1549,N_1487,N_1480);
xnor U1550 (N_1550,N_1505,N_1521);
nor U1551 (N_1551,N_1528,N_1503);
xor U1552 (N_1552,N_1501,N_1523);
nor U1553 (N_1553,N_1544,N_1540);
nor U1554 (N_1554,N_1507,N_1506);
or U1555 (N_1555,N_1511,N_1532);
xnor U1556 (N_1556,N_1546,N_1527);
nand U1557 (N_1557,N_1535,N_1549);
and U1558 (N_1558,N_1533,N_1512);
xnor U1559 (N_1559,N_1514,N_1500);
nand U1560 (N_1560,N_1502,N_1539);
nor U1561 (N_1561,N_1515,N_1545);
nand U1562 (N_1562,N_1548,N_1510);
or U1563 (N_1563,N_1524,N_1519);
nand U1564 (N_1564,N_1537,N_1538);
and U1565 (N_1565,N_1509,N_1518);
nor U1566 (N_1566,N_1534,N_1504);
nor U1567 (N_1567,N_1542,N_1529);
nand U1568 (N_1568,N_1522,N_1520);
xor U1569 (N_1569,N_1547,N_1517);
xor U1570 (N_1570,N_1508,N_1543);
or U1571 (N_1571,N_1526,N_1531);
nand U1572 (N_1572,N_1516,N_1525);
or U1573 (N_1573,N_1541,N_1530);
nor U1574 (N_1574,N_1536,N_1513);
and U1575 (N_1575,N_1548,N_1506);
nor U1576 (N_1576,N_1547,N_1524);
and U1577 (N_1577,N_1524,N_1512);
or U1578 (N_1578,N_1505,N_1525);
or U1579 (N_1579,N_1508,N_1523);
nor U1580 (N_1580,N_1506,N_1540);
nor U1581 (N_1581,N_1547,N_1512);
nor U1582 (N_1582,N_1524,N_1508);
xnor U1583 (N_1583,N_1527,N_1549);
or U1584 (N_1584,N_1517,N_1509);
or U1585 (N_1585,N_1532,N_1547);
nor U1586 (N_1586,N_1512,N_1546);
nor U1587 (N_1587,N_1542,N_1513);
nor U1588 (N_1588,N_1547,N_1529);
nand U1589 (N_1589,N_1514,N_1524);
nand U1590 (N_1590,N_1529,N_1506);
nand U1591 (N_1591,N_1522,N_1503);
and U1592 (N_1592,N_1531,N_1523);
xnor U1593 (N_1593,N_1544,N_1515);
xor U1594 (N_1594,N_1536,N_1515);
and U1595 (N_1595,N_1514,N_1507);
or U1596 (N_1596,N_1541,N_1547);
nand U1597 (N_1597,N_1502,N_1524);
or U1598 (N_1598,N_1517,N_1507);
or U1599 (N_1599,N_1530,N_1510);
nor U1600 (N_1600,N_1552,N_1570);
and U1601 (N_1601,N_1584,N_1591);
or U1602 (N_1602,N_1586,N_1581);
and U1603 (N_1603,N_1551,N_1589);
xnor U1604 (N_1604,N_1582,N_1573);
nor U1605 (N_1605,N_1594,N_1553);
nand U1606 (N_1606,N_1593,N_1554);
and U1607 (N_1607,N_1564,N_1588);
or U1608 (N_1608,N_1592,N_1558);
nor U1609 (N_1609,N_1568,N_1571);
xnor U1610 (N_1610,N_1550,N_1555);
nor U1611 (N_1611,N_1595,N_1579);
nor U1612 (N_1612,N_1572,N_1566);
xor U1613 (N_1613,N_1578,N_1587);
xnor U1614 (N_1614,N_1597,N_1590);
and U1615 (N_1615,N_1561,N_1575);
or U1616 (N_1616,N_1596,N_1577);
or U1617 (N_1617,N_1576,N_1556);
nand U1618 (N_1618,N_1583,N_1557);
xnor U1619 (N_1619,N_1574,N_1569);
and U1620 (N_1620,N_1580,N_1599);
nand U1621 (N_1621,N_1585,N_1565);
and U1622 (N_1622,N_1598,N_1559);
xor U1623 (N_1623,N_1562,N_1560);
nand U1624 (N_1624,N_1563,N_1567);
and U1625 (N_1625,N_1581,N_1599);
nand U1626 (N_1626,N_1577,N_1552);
and U1627 (N_1627,N_1594,N_1582);
nand U1628 (N_1628,N_1580,N_1594);
nand U1629 (N_1629,N_1572,N_1561);
nand U1630 (N_1630,N_1568,N_1579);
or U1631 (N_1631,N_1593,N_1562);
nand U1632 (N_1632,N_1553,N_1593);
nor U1633 (N_1633,N_1585,N_1593);
xnor U1634 (N_1634,N_1571,N_1578);
xor U1635 (N_1635,N_1598,N_1596);
nor U1636 (N_1636,N_1598,N_1587);
or U1637 (N_1637,N_1553,N_1582);
nand U1638 (N_1638,N_1558,N_1561);
xnor U1639 (N_1639,N_1583,N_1560);
or U1640 (N_1640,N_1572,N_1586);
nor U1641 (N_1641,N_1550,N_1568);
or U1642 (N_1642,N_1578,N_1594);
nand U1643 (N_1643,N_1559,N_1557);
xor U1644 (N_1644,N_1558,N_1554);
nand U1645 (N_1645,N_1552,N_1568);
xor U1646 (N_1646,N_1599,N_1588);
nand U1647 (N_1647,N_1574,N_1553);
xor U1648 (N_1648,N_1582,N_1567);
xor U1649 (N_1649,N_1570,N_1579);
nand U1650 (N_1650,N_1622,N_1620);
or U1651 (N_1651,N_1624,N_1649);
nor U1652 (N_1652,N_1616,N_1606);
nand U1653 (N_1653,N_1645,N_1633);
nand U1654 (N_1654,N_1621,N_1637);
xnor U1655 (N_1655,N_1605,N_1635);
xnor U1656 (N_1656,N_1601,N_1634);
nor U1657 (N_1657,N_1640,N_1630);
xor U1658 (N_1658,N_1647,N_1612);
or U1659 (N_1659,N_1648,N_1642);
and U1660 (N_1660,N_1614,N_1600);
or U1661 (N_1661,N_1636,N_1617);
and U1662 (N_1662,N_1628,N_1641);
nand U1663 (N_1663,N_1613,N_1644);
or U1664 (N_1664,N_1632,N_1643);
and U1665 (N_1665,N_1602,N_1646);
and U1666 (N_1666,N_1604,N_1629);
or U1667 (N_1667,N_1611,N_1609);
or U1668 (N_1668,N_1639,N_1603);
xnor U1669 (N_1669,N_1626,N_1619);
and U1670 (N_1670,N_1623,N_1638);
or U1671 (N_1671,N_1631,N_1618);
and U1672 (N_1672,N_1610,N_1607);
and U1673 (N_1673,N_1627,N_1625);
xnor U1674 (N_1674,N_1615,N_1608);
nand U1675 (N_1675,N_1646,N_1628);
nor U1676 (N_1676,N_1616,N_1622);
or U1677 (N_1677,N_1611,N_1649);
xor U1678 (N_1678,N_1647,N_1645);
xor U1679 (N_1679,N_1634,N_1628);
nand U1680 (N_1680,N_1632,N_1615);
nor U1681 (N_1681,N_1622,N_1610);
nor U1682 (N_1682,N_1626,N_1612);
or U1683 (N_1683,N_1607,N_1626);
and U1684 (N_1684,N_1619,N_1623);
nor U1685 (N_1685,N_1617,N_1609);
and U1686 (N_1686,N_1648,N_1617);
or U1687 (N_1687,N_1604,N_1623);
or U1688 (N_1688,N_1634,N_1613);
and U1689 (N_1689,N_1632,N_1623);
nor U1690 (N_1690,N_1614,N_1644);
and U1691 (N_1691,N_1636,N_1622);
or U1692 (N_1692,N_1638,N_1636);
xnor U1693 (N_1693,N_1619,N_1625);
nand U1694 (N_1694,N_1616,N_1633);
nor U1695 (N_1695,N_1629,N_1601);
nor U1696 (N_1696,N_1620,N_1606);
nor U1697 (N_1697,N_1636,N_1610);
or U1698 (N_1698,N_1604,N_1633);
and U1699 (N_1699,N_1631,N_1619);
nor U1700 (N_1700,N_1650,N_1684);
or U1701 (N_1701,N_1691,N_1694);
and U1702 (N_1702,N_1697,N_1695);
or U1703 (N_1703,N_1674,N_1652);
or U1704 (N_1704,N_1696,N_1688);
xor U1705 (N_1705,N_1672,N_1654);
nor U1706 (N_1706,N_1683,N_1670);
nor U1707 (N_1707,N_1653,N_1699);
nor U1708 (N_1708,N_1685,N_1689);
and U1709 (N_1709,N_1665,N_1678);
nand U1710 (N_1710,N_1667,N_1679);
nand U1711 (N_1711,N_1676,N_1659);
nor U1712 (N_1712,N_1651,N_1658);
xnor U1713 (N_1713,N_1680,N_1692);
nand U1714 (N_1714,N_1656,N_1661);
nor U1715 (N_1715,N_1698,N_1673);
xnor U1716 (N_1716,N_1666,N_1655);
or U1717 (N_1717,N_1664,N_1663);
and U1718 (N_1718,N_1669,N_1686);
nand U1719 (N_1719,N_1677,N_1687);
and U1720 (N_1720,N_1690,N_1668);
or U1721 (N_1721,N_1675,N_1662);
and U1722 (N_1722,N_1671,N_1682);
nor U1723 (N_1723,N_1681,N_1660);
or U1724 (N_1724,N_1657,N_1693);
nand U1725 (N_1725,N_1689,N_1684);
nor U1726 (N_1726,N_1659,N_1668);
and U1727 (N_1727,N_1654,N_1671);
nor U1728 (N_1728,N_1673,N_1691);
xnor U1729 (N_1729,N_1678,N_1651);
and U1730 (N_1730,N_1687,N_1658);
nor U1731 (N_1731,N_1697,N_1676);
nand U1732 (N_1732,N_1657,N_1659);
and U1733 (N_1733,N_1699,N_1679);
and U1734 (N_1734,N_1695,N_1658);
xnor U1735 (N_1735,N_1662,N_1670);
nand U1736 (N_1736,N_1666,N_1656);
and U1737 (N_1737,N_1678,N_1653);
or U1738 (N_1738,N_1699,N_1694);
and U1739 (N_1739,N_1667,N_1697);
nand U1740 (N_1740,N_1655,N_1676);
xor U1741 (N_1741,N_1670,N_1656);
xor U1742 (N_1742,N_1677,N_1691);
or U1743 (N_1743,N_1656,N_1677);
xor U1744 (N_1744,N_1677,N_1670);
or U1745 (N_1745,N_1690,N_1691);
and U1746 (N_1746,N_1692,N_1653);
xnor U1747 (N_1747,N_1654,N_1665);
and U1748 (N_1748,N_1670,N_1690);
or U1749 (N_1749,N_1659,N_1688);
xnor U1750 (N_1750,N_1709,N_1728);
xor U1751 (N_1751,N_1736,N_1702);
or U1752 (N_1752,N_1713,N_1744);
xor U1753 (N_1753,N_1717,N_1747);
nor U1754 (N_1754,N_1727,N_1730);
or U1755 (N_1755,N_1738,N_1743);
xor U1756 (N_1756,N_1714,N_1742);
nor U1757 (N_1757,N_1710,N_1731);
nor U1758 (N_1758,N_1748,N_1749);
and U1759 (N_1759,N_1716,N_1708);
or U1760 (N_1760,N_1739,N_1735);
nor U1761 (N_1761,N_1705,N_1706);
or U1762 (N_1762,N_1700,N_1704);
nor U1763 (N_1763,N_1723,N_1729);
nand U1764 (N_1764,N_1740,N_1722);
xnor U1765 (N_1765,N_1726,N_1719);
nand U1766 (N_1766,N_1725,N_1721);
or U1767 (N_1767,N_1745,N_1733);
xnor U1768 (N_1768,N_1732,N_1720);
nor U1769 (N_1769,N_1724,N_1715);
nor U1770 (N_1770,N_1711,N_1737);
or U1771 (N_1771,N_1707,N_1734);
nor U1772 (N_1772,N_1712,N_1701);
and U1773 (N_1773,N_1741,N_1746);
or U1774 (N_1774,N_1703,N_1718);
nand U1775 (N_1775,N_1747,N_1714);
or U1776 (N_1776,N_1717,N_1731);
nand U1777 (N_1777,N_1711,N_1743);
nand U1778 (N_1778,N_1719,N_1715);
and U1779 (N_1779,N_1741,N_1743);
and U1780 (N_1780,N_1702,N_1737);
and U1781 (N_1781,N_1728,N_1739);
nor U1782 (N_1782,N_1715,N_1705);
or U1783 (N_1783,N_1747,N_1701);
and U1784 (N_1784,N_1716,N_1702);
nand U1785 (N_1785,N_1717,N_1718);
xnor U1786 (N_1786,N_1722,N_1721);
xnor U1787 (N_1787,N_1740,N_1733);
xor U1788 (N_1788,N_1728,N_1722);
or U1789 (N_1789,N_1737,N_1744);
xor U1790 (N_1790,N_1731,N_1724);
and U1791 (N_1791,N_1723,N_1731);
nand U1792 (N_1792,N_1744,N_1707);
nand U1793 (N_1793,N_1729,N_1711);
nor U1794 (N_1794,N_1741,N_1733);
or U1795 (N_1795,N_1715,N_1711);
and U1796 (N_1796,N_1705,N_1730);
and U1797 (N_1797,N_1712,N_1726);
nor U1798 (N_1798,N_1740,N_1716);
nand U1799 (N_1799,N_1747,N_1713);
nor U1800 (N_1800,N_1772,N_1786);
or U1801 (N_1801,N_1769,N_1771);
nand U1802 (N_1802,N_1782,N_1775);
xor U1803 (N_1803,N_1780,N_1756);
xnor U1804 (N_1804,N_1778,N_1753);
nor U1805 (N_1805,N_1752,N_1776);
or U1806 (N_1806,N_1773,N_1759);
nor U1807 (N_1807,N_1792,N_1784);
xor U1808 (N_1808,N_1755,N_1754);
nand U1809 (N_1809,N_1788,N_1794);
nor U1810 (N_1810,N_1757,N_1789);
nand U1811 (N_1811,N_1777,N_1760);
and U1812 (N_1812,N_1766,N_1799);
xor U1813 (N_1813,N_1793,N_1796);
nand U1814 (N_1814,N_1750,N_1768);
nand U1815 (N_1815,N_1791,N_1781);
and U1816 (N_1816,N_1751,N_1795);
or U1817 (N_1817,N_1798,N_1762);
nor U1818 (N_1818,N_1774,N_1765);
xnor U1819 (N_1819,N_1764,N_1767);
and U1820 (N_1820,N_1790,N_1783);
nand U1821 (N_1821,N_1761,N_1770);
nor U1822 (N_1822,N_1787,N_1785);
xnor U1823 (N_1823,N_1763,N_1779);
or U1824 (N_1824,N_1758,N_1797);
and U1825 (N_1825,N_1792,N_1796);
nor U1826 (N_1826,N_1795,N_1761);
nand U1827 (N_1827,N_1795,N_1787);
nand U1828 (N_1828,N_1753,N_1795);
nor U1829 (N_1829,N_1776,N_1770);
nand U1830 (N_1830,N_1798,N_1774);
and U1831 (N_1831,N_1759,N_1767);
and U1832 (N_1832,N_1796,N_1764);
xnor U1833 (N_1833,N_1767,N_1792);
and U1834 (N_1834,N_1792,N_1777);
nand U1835 (N_1835,N_1767,N_1766);
or U1836 (N_1836,N_1781,N_1794);
and U1837 (N_1837,N_1791,N_1755);
or U1838 (N_1838,N_1792,N_1753);
nor U1839 (N_1839,N_1764,N_1782);
nor U1840 (N_1840,N_1783,N_1759);
and U1841 (N_1841,N_1796,N_1755);
nand U1842 (N_1842,N_1799,N_1774);
and U1843 (N_1843,N_1753,N_1793);
nor U1844 (N_1844,N_1798,N_1763);
nand U1845 (N_1845,N_1767,N_1798);
or U1846 (N_1846,N_1759,N_1755);
xor U1847 (N_1847,N_1784,N_1791);
and U1848 (N_1848,N_1782,N_1769);
xnor U1849 (N_1849,N_1767,N_1778);
nor U1850 (N_1850,N_1847,N_1818);
and U1851 (N_1851,N_1810,N_1844);
nand U1852 (N_1852,N_1802,N_1828);
and U1853 (N_1853,N_1820,N_1830);
nor U1854 (N_1854,N_1803,N_1839);
xor U1855 (N_1855,N_1817,N_1834);
nor U1856 (N_1856,N_1827,N_1842);
and U1857 (N_1857,N_1807,N_1809);
and U1858 (N_1858,N_1832,N_1814);
nor U1859 (N_1859,N_1816,N_1835);
or U1860 (N_1860,N_1806,N_1833);
or U1861 (N_1861,N_1819,N_1825);
nand U1862 (N_1862,N_1849,N_1804);
and U1863 (N_1863,N_1811,N_1848);
xnor U1864 (N_1864,N_1846,N_1837);
nand U1865 (N_1865,N_1826,N_1813);
nand U1866 (N_1866,N_1805,N_1823);
xor U1867 (N_1867,N_1840,N_1812);
nor U1868 (N_1868,N_1838,N_1808);
nor U1869 (N_1869,N_1829,N_1801);
xor U1870 (N_1870,N_1836,N_1800);
and U1871 (N_1871,N_1822,N_1815);
nor U1872 (N_1872,N_1824,N_1841);
nor U1873 (N_1873,N_1831,N_1845);
and U1874 (N_1874,N_1821,N_1843);
and U1875 (N_1875,N_1808,N_1809);
xor U1876 (N_1876,N_1845,N_1838);
nor U1877 (N_1877,N_1840,N_1830);
or U1878 (N_1878,N_1828,N_1848);
nor U1879 (N_1879,N_1802,N_1819);
and U1880 (N_1880,N_1829,N_1828);
nand U1881 (N_1881,N_1810,N_1840);
or U1882 (N_1882,N_1849,N_1845);
or U1883 (N_1883,N_1807,N_1831);
nor U1884 (N_1884,N_1834,N_1820);
and U1885 (N_1885,N_1838,N_1803);
nor U1886 (N_1886,N_1800,N_1803);
and U1887 (N_1887,N_1842,N_1814);
nor U1888 (N_1888,N_1800,N_1823);
or U1889 (N_1889,N_1836,N_1829);
and U1890 (N_1890,N_1816,N_1842);
nor U1891 (N_1891,N_1823,N_1837);
and U1892 (N_1892,N_1823,N_1808);
nor U1893 (N_1893,N_1844,N_1802);
nand U1894 (N_1894,N_1808,N_1806);
nand U1895 (N_1895,N_1811,N_1800);
nor U1896 (N_1896,N_1849,N_1807);
or U1897 (N_1897,N_1814,N_1818);
or U1898 (N_1898,N_1815,N_1828);
nor U1899 (N_1899,N_1824,N_1810);
xor U1900 (N_1900,N_1886,N_1852);
and U1901 (N_1901,N_1885,N_1867);
and U1902 (N_1902,N_1864,N_1887);
nor U1903 (N_1903,N_1858,N_1897);
nor U1904 (N_1904,N_1894,N_1851);
and U1905 (N_1905,N_1890,N_1884);
nand U1906 (N_1906,N_1881,N_1891);
and U1907 (N_1907,N_1869,N_1888);
xnor U1908 (N_1908,N_1883,N_1876);
or U1909 (N_1909,N_1878,N_1874);
nand U1910 (N_1910,N_1880,N_1859);
and U1911 (N_1911,N_1896,N_1892);
nand U1912 (N_1912,N_1871,N_1889);
and U1913 (N_1913,N_1877,N_1873);
xor U1914 (N_1914,N_1882,N_1865);
and U1915 (N_1915,N_1879,N_1854);
xnor U1916 (N_1916,N_1857,N_1850);
xor U1917 (N_1917,N_1856,N_1863);
or U1918 (N_1918,N_1862,N_1866);
and U1919 (N_1919,N_1899,N_1872);
nor U1920 (N_1920,N_1895,N_1893);
or U1921 (N_1921,N_1898,N_1853);
xnor U1922 (N_1922,N_1861,N_1860);
nor U1923 (N_1923,N_1855,N_1875);
nand U1924 (N_1924,N_1870,N_1868);
nor U1925 (N_1925,N_1874,N_1890);
xor U1926 (N_1926,N_1852,N_1884);
nand U1927 (N_1927,N_1878,N_1879);
xor U1928 (N_1928,N_1874,N_1876);
xnor U1929 (N_1929,N_1875,N_1874);
nor U1930 (N_1930,N_1899,N_1895);
or U1931 (N_1931,N_1857,N_1875);
or U1932 (N_1932,N_1871,N_1893);
or U1933 (N_1933,N_1893,N_1886);
xnor U1934 (N_1934,N_1860,N_1870);
nor U1935 (N_1935,N_1871,N_1855);
xnor U1936 (N_1936,N_1885,N_1887);
xnor U1937 (N_1937,N_1850,N_1899);
nand U1938 (N_1938,N_1880,N_1851);
xor U1939 (N_1939,N_1863,N_1875);
or U1940 (N_1940,N_1867,N_1880);
xor U1941 (N_1941,N_1860,N_1872);
nand U1942 (N_1942,N_1857,N_1856);
xnor U1943 (N_1943,N_1861,N_1868);
xnor U1944 (N_1944,N_1881,N_1894);
nor U1945 (N_1945,N_1873,N_1893);
nor U1946 (N_1946,N_1858,N_1870);
and U1947 (N_1947,N_1872,N_1861);
and U1948 (N_1948,N_1853,N_1852);
nand U1949 (N_1949,N_1854,N_1882);
xor U1950 (N_1950,N_1902,N_1924);
xnor U1951 (N_1951,N_1947,N_1918);
nand U1952 (N_1952,N_1932,N_1942);
and U1953 (N_1953,N_1938,N_1922);
nand U1954 (N_1954,N_1933,N_1945);
or U1955 (N_1955,N_1904,N_1939);
nor U1956 (N_1956,N_1909,N_1919);
and U1957 (N_1957,N_1920,N_1915);
nor U1958 (N_1958,N_1928,N_1903);
nand U1959 (N_1959,N_1906,N_1948);
and U1960 (N_1960,N_1917,N_1944);
or U1961 (N_1961,N_1936,N_1910);
or U1962 (N_1962,N_1911,N_1912);
xnor U1963 (N_1963,N_1930,N_1914);
xnor U1964 (N_1964,N_1923,N_1949);
and U1965 (N_1965,N_1937,N_1901);
xor U1966 (N_1966,N_1927,N_1941);
xor U1967 (N_1967,N_1926,N_1913);
xor U1968 (N_1968,N_1940,N_1905);
xnor U1969 (N_1969,N_1900,N_1935);
xor U1970 (N_1970,N_1929,N_1943);
xnor U1971 (N_1971,N_1916,N_1931);
nand U1972 (N_1972,N_1946,N_1907);
or U1973 (N_1973,N_1934,N_1921);
and U1974 (N_1974,N_1908,N_1925);
xnor U1975 (N_1975,N_1917,N_1925);
and U1976 (N_1976,N_1948,N_1942);
xnor U1977 (N_1977,N_1902,N_1947);
and U1978 (N_1978,N_1919,N_1924);
xor U1979 (N_1979,N_1900,N_1916);
and U1980 (N_1980,N_1909,N_1900);
xnor U1981 (N_1981,N_1945,N_1948);
nand U1982 (N_1982,N_1948,N_1924);
nor U1983 (N_1983,N_1946,N_1944);
xnor U1984 (N_1984,N_1927,N_1929);
xor U1985 (N_1985,N_1943,N_1903);
or U1986 (N_1986,N_1902,N_1939);
nand U1987 (N_1987,N_1945,N_1927);
xnor U1988 (N_1988,N_1924,N_1918);
or U1989 (N_1989,N_1906,N_1919);
or U1990 (N_1990,N_1940,N_1916);
and U1991 (N_1991,N_1935,N_1928);
and U1992 (N_1992,N_1909,N_1938);
nand U1993 (N_1993,N_1917,N_1928);
nor U1994 (N_1994,N_1909,N_1944);
and U1995 (N_1995,N_1941,N_1949);
xor U1996 (N_1996,N_1930,N_1900);
xnor U1997 (N_1997,N_1937,N_1924);
nand U1998 (N_1998,N_1940,N_1934);
nor U1999 (N_1999,N_1938,N_1921);
and U2000 (N_2000,N_1974,N_1956);
nand U2001 (N_2001,N_1959,N_1980);
xor U2002 (N_2002,N_1985,N_1972);
xnor U2003 (N_2003,N_1968,N_1984);
or U2004 (N_2004,N_1966,N_1994);
or U2005 (N_2005,N_1997,N_1996);
and U2006 (N_2006,N_1998,N_1955);
nor U2007 (N_2007,N_1951,N_1995);
and U2008 (N_2008,N_1975,N_1989);
xnor U2009 (N_2009,N_1961,N_1982);
or U2010 (N_2010,N_1962,N_1973);
and U2011 (N_2011,N_1960,N_1967);
nor U2012 (N_2012,N_1964,N_1993);
nand U2013 (N_2013,N_1970,N_1965);
nand U2014 (N_2014,N_1954,N_1990);
and U2015 (N_2015,N_1963,N_1957);
nand U2016 (N_2016,N_1981,N_1979);
or U2017 (N_2017,N_1950,N_1976);
or U2018 (N_2018,N_1958,N_1983);
nor U2019 (N_2019,N_1953,N_1999);
xnor U2020 (N_2020,N_1987,N_1988);
nor U2021 (N_2021,N_1992,N_1952);
nand U2022 (N_2022,N_1986,N_1991);
or U2023 (N_2023,N_1969,N_1977);
and U2024 (N_2024,N_1971,N_1978);
or U2025 (N_2025,N_1990,N_1995);
xnor U2026 (N_2026,N_1970,N_1962);
and U2027 (N_2027,N_1982,N_1959);
nor U2028 (N_2028,N_1995,N_1980);
xnor U2029 (N_2029,N_1982,N_1967);
and U2030 (N_2030,N_1959,N_1970);
or U2031 (N_2031,N_1965,N_1956);
and U2032 (N_2032,N_1958,N_1972);
nand U2033 (N_2033,N_1953,N_1980);
nor U2034 (N_2034,N_1965,N_1973);
xnor U2035 (N_2035,N_1959,N_1962);
or U2036 (N_2036,N_1952,N_1973);
xor U2037 (N_2037,N_1991,N_1980);
nand U2038 (N_2038,N_1978,N_1972);
xnor U2039 (N_2039,N_1965,N_1983);
nor U2040 (N_2040,N_1969,N_1976);
xnor U2041 (N_2041,N_1978,N_1999);
and U2042 (N_2042,N_1968,N_1966);
and U2043 (N_2043,N_1966,N_1972);
nand U2044 (N_2044,N_1988,N_1979);
xor U2045 (N_2045,N_1998,N_1950);
xnor U2046 (N_2046,N_1975,N_1964);
nand U2047 (N_2047,N_1963,N_1998);
xor U2048 (N_2048,N_1993,N_1957);
xor U2049 (N_2049,N_1981,N_1978);
xnor U2050 (N_2050,N_2018,N_2015);
or U2051 (N_2051,N_2030,N_2008);
nor U2052 (N_2052,N_2003,N_2046);
nand U2053 (N_2053,N_2031,N_2029);
nand U2054 (N_2054,N_2026,N_2043);
xnor U2055 (N_2055,N_2034,N_2012);
xnor U2056 (N_2056,N_2011,N_2006);
nor U2057 (N_2057,N_2014,N_2004);
xor U2058 (N_2058,N_2047,N_2013);
xnor U2059 (N_2059,N_2045,N_2020);
or U2060 (N_2060,N_2021,N_2028);
or U2061 (N_2061,N_2019,N_2037);
or U2062 (N_2062,N_2039,N_2048);
and U2063 (N_2063,N_2001,N_2044);
nand U2064 (N_2064,N_2035,N_2016);
nor U2065 (N_2065,N_2017,N_2000);
nor U2066 (N_2066,N_2027,N_2005);
and U2067 (N_2067,N_2007,N_2024);
or U2068 (N_2068,N_2041,N_2049);
nor U2069 (N_2069,N_2033,N_2038);
and U2070 (N_2070,N_2009,N_2010);
or U2071 (N_2071,N_2036,N_2042);
nand U2072 (N_2072,N_2032,N_2022);
xnor U2073 (N_2073,N_2002,N_2040);
or U2074 (N_2074,N_2023,N_2025);
or U2075 (N_2075,N_2034,N_2038);
nand U2076 (N_2076,N_2022,N_2049);
nor U2077 (N_2077,N_2048,N_2028);
or U2078 (N_2078,N_2020,N_2032);
nand U2079 (N_2079,N_2021,N_2008);
nand U2080 (N_2080,N_2029,N_2016);
and U2081 (N_2081,N_2026,N_2000);
nor U2082 (N_2082,N_2037,N_2002);
nand U2083 (N_2083,N_2016,N_2038);
nor U2084 (N_2084,N_2002,N_2000);
or U2085 (N_2085,N_2020,N_2019);
and U2086 (N_2086,N_2034,N_2049);
nor U2087 (N_2087,N_2042,N_2025);
nor U2088 (N_2088,N_2016,N_2009);
and U2089 (N_2089,N_2007,N_2044);
or U2090 (N_2090,N_2022,N_2031);
or U2091 (N_2091,N_2040,N_2048);
xnor U2092 (N_2092,N_2047,N_2016);
nand U2093 (N_2093,N_2011,N_2048);
and U2094 (N_2094,N_2026,N_2032);
or U2095 (N_2095,N_2002,N_2024);
nor U2096 (N_2096,N_2005,N_2007);
nor U2097 (N_2097,N_2009,N_2006);
and U2098 (N_2098,N_2039,N_2025);
or U2099 (N_2099,N_2015,N_2027);
nor U2100 (N_2100,N_2053,N_2068);
xor U2101 (N_2101,N_2071,N_2081);
nand U2102 (N_2102,N_2064,N_2054);
xor U2103 (N_2103,N_2097,N_2087);
nand U2104 (N_2104,N_2060,N_2072);
xnor U2105 (N_2105,N_2063,N_2069);
nor U2106 (N_2106,N_2088,N_2078);
and U2107 (N_2107,N_2075,N_2086);
or U2108 (N_2108,N_2089,N_2061);
and U2109 (N_2109,N_2091,N_2082);
xor U2110 (N_2110,N_2058,N_2074);
xnor U2111 (N_2111,N_2084,N_2055);
or U2112 (N_2112,N_2057,N_2093);
nand U2113 (N_2113,N_2066,N_2090);
nand U2114 (N_2114,N_2073,N_2095);
nor U2115 (N_2115,N_2077,N_2079);
nand U2116 (N_2116,N_2056,N_2070);
and U2117 (N_2117,N_2059,N_2052);
nor U2118 (N_2118,N_2085,N_2099);
and U2119 (N_2119,N_2050,N_2080);
or U2120 (N_2120,N_2076,N_2092);
or U2121 (N_2121,N_2094,N_2083);
xor U2122 (N_2122,N_2098,N_2065);
and U2123 (N_2123,N_2062,N_2051);
xnor U2124 (N_2124,N_2067,N_2096);
nand U2125 (N_2125,N_2067,N_2076);
and U2126 (N_2126,N_2064,N_2059);
and U2127 (N_2127,N_2076,N_2084);
or U2128 (N_2128,N_2070,N_2074);
xor U2129 (N_2129,N_2066,N_2088);
or U2130 (N_2130,N_2075,N_2051);
and U2131 (N_2131,N_2064,N_2092);
or U2132 (N_2132,N_2097,N_2066);
or U2133 (N_2133,N_2065,N_2077);
nand U2134 (N_2134,N_2068,N_2093);
nand U2135 (N_2135,N_2050,N_2054);
xnor U2136 (N_2136,N_2051,N_2053);
and U2137 (N_2137,N_2064,N_2052);
or U2138 (N_2138,N_2078,N_2053);
and U2139 (N_2139,N_2077,N_2059);
nand U2140 (N_2140,N_2054,N_2061);
nand U2141 (N_2141,N_2087,N_2093);
and U2142 (N_2142,N_2067,N_2084);
or U2143 (N_2143,N_2060,N_2052);
nand U2144 (N_2144,N_2059,N_2092);
nor U2145 (N_2145,N_2097,N_2053);
or U2146 (N_2146,N_2064,N_2058);
nand U2147 (N_2147,N_2092,N_2055);
nor U2148 (N_2148,N_2066,N_2065);
nand U2149 (N_2149,N_2089,N_2079);
and U2150 (N_2150,N_2118,N_2123);
nor U2151 (N_2151,N_2104,N_2106);
and U2152 (N_2152,N_2140,N_2117);
or U2153 (N_2153,N_2107,N_2127);
or U2154 (N_2154,N_2124,N_2128);
or U2155 (N_2155,N_2136,N_2135);
nand U2156 (N_2156,N_2125,N_2116);
and U2157 (N_2157,N_2105,N_2148);
nand U2158 (N_2158,N_2130,N_2132);
and U2159 (N_2159,N_2138,N_2131);
xnor U2160 (N_2160,N_2146,N_2114);
or U2161 (N_2161,N_2108,N_2126);
or U2162 (N_2162,N_2122,N_2101);
nor U2163 (N_2163,N_2149,N_2133);
xor U2164 (N_2164,N_2100,N_2139);
nor U2165 (N_2165,N_2113,N_2147);
or U2166 (N_2166,N_2119,N_2142);
and U2167 (N_2167,N_2102,N_2120);
xor U2168 (N_2168,N_2134,N_2111);
xor U2169 (N_2169,N_2144,N_2129);
and U2170 (N_2170,N_2110,N_2103);
or U2171 (N_2171,N_2112,N_2137);
and U2172 (N_2172,N_2145,N_2143);
and U2173 (N_2173,N_2141,N_2109);
and U2174 (N_2174,N_2115,N_2121);
or U2175 (N_2175,N_2127,N_2109);
nand U2176 (N_2176,N_2131,N_2121);
xor U2177 (N_2177,N_2119,N_2141);
and U2178 (N_2178,N_2136,N_2124);
and U2179 (N_2179,N_2145,N_2108);
xnor U2180 (N_2180,N_2108,N_2102);
nand U2181 (N_2181,N_2127,N_2108);
nand U2182 (N_2182,N_2128,N_2104);
nand U2183 (N_2183,N_2116,N_2142);
nand U2184 (N_2184,N_2144,N_2132);
nand U2185 (N_2185,N_2135,N_2149);
nand U2186 (N_2186,N_2142,N_2126);
nand U2187 (N_2187,N_2109,N_2137);
nor U2188 (N_2188,N_2108,N_2105);
and U2189 (N_2189,N_2124,N_2142);
nand U2190 (N_2190,N_2120,N_2133);
and U2191 (N_2191,N_2104,N_2118);
nand U2192 (N_2192,N_2133,N_2128);
xnor U2193 (N_2193,N_2115,N_2102);
and U2194 (N_2194,N_2106,N_2107);
nand U2195 (N_2195,N_2146,N_2123);
or U2196 (N_2196,N_2142,N_2114);
xor U2197 (N_2197,N_2117,N_2102);
xnor U2198 (N_2198,N_2100,N_2104);
nand U2199 (N_2199,N_2147,N_2121);
or U2200 (N_2200,N_2198,N_2157);
nand U2201 (N_2201,N_2152,N_2195);
nor U2202 (N_2202,N_2174,N_2169);
nor U2203 (N_2203,N_2189,N_2184);
or U2204 (N_2204,N_2150,N_2182);
xor U2205 (N_2205,N_2190,N_2160);
or U2206 (N_2206,N_2159,N_2197);
and U2207 (N_2207,N_2181,N_2199);
nor U2208 (N_2208,N_2186,N_2171);
nor U2209 (N_2209,N_2155,N_2168);
nor U2210 (N_2210,N_2187,N_2167);
or U2211 (N_2211,N_2192,N_2153);
nor U2212 (N_2212,N_2177,N_2178);
and U2213 (N_2213,N_2172,N_2163);
nand U2214 (N_2214,N_2196,N_2170);
or U2215 (N_2215,N_2180,N_2154);
xnor U2216 (N_2216,N_2188,N_2191);
or U2217 (N_2217,N_2194,N_2166);
xor U2218 (N_2218,N_2175,N_2156);
nand U2219 (N_2219,N_2164,N_2185);
xor U2220 (N_2220,N_2151,N_2179);
or U2221 (N_2221,N_2193,N_2176);
nor U2222 (N_2222,N_2165,N_2158);
or U2223 (N_2223,N_2161,N_2183);
nor U2224 (N_2224,N_2173,N_2162);
and U2225 (N_2225,N_2160,N_2199);
and U2226 (N_2226,N_2180,N_2173);
nand U2227 (N_2227,N_2154,N_2187);
nor U2228 (N_2228,N_2187,N_2175);
xnor U2229 (N_2229,N_2185,N_2157);
and U2230 (N_2230,N_2172,N_2184);
or U2231 (N_2231,N_2181,N_2170);
or U2232 (N_2232,N_2154,N_2175);
nand U2233 (N_2233,N_2163,N_2174);
or U2234 (N_2234,N_2182,N_2166);
nand U2235 (N_2235,N_2192,N_2198);
or U2236 (N_2236,N_2198,N_2193);
and U2237 (N_2237,N_2157,N_2197);
xor U2238 (N_2238,N_2180,N_2170);
or U2239 (N_2239,N_2186,N_2169);
nor U2240 (N_2240,N_2170,N_2166);
and U2241 (N_2241,N_2162,N_2158);
nor U2242 (N_2242,N_2154,N_2194);
nor U2243 (N_2243,N_2152,N_2155);
or U2244 (N_2244,N_2183,N_2152);
xnor U2245 (N_2245,N_2171,N_2165);
nor U2246 (N_2246,N_2181,N_2198);
nor U2247 (N_2247,N_2155,N_2166);
or U2248 (N_2248,N_2174,N_2191);
nand U2249 (N_2249,N_2153,N_2191);
or U2250 (N_2250,N_2235,N_2219);
xnor U2251 (N_2251,N_2230,N_2209);
xor U2252 (N_2252,N_2215,N_2222);
nand U2253 (N_2253,N_2240,N_2217);
and U2254 (N_2254,N_2244,N_2206);
nor U2255 (N_2255,N_2205,N_2227);
and U2256 (N_2256,N_2243,N_2247);
nand U2257 (N_2257,N_2238,N_2220);
xor U2258 (N_2258,N_2200,N_2225);
or U2259 (N_2259,N_2213,N_2237);
or U2260 (N_2260,N_2211,N_2229);
nand U2261 (N_2261,N_2236,N_2226);
or U2262 (N_2262,N_2216,N_2214);
and U2263 (N_2263,N_2248,N_2221);
or U2264 (N_2264,N_2241,N_2234);
nor U2265 (N_2265,N_2232,N_2246);
nand U2266 (N_2266,N_2212,N_2201);
nand U2267 (N_2267,N_2228,N_2239);
nor U2268 (N_2268,N_2207,N_2203);
and U2269 (N_2269,N_2208,N_2242);
and U2270 (N_2270,N_2249,N_2224);
nor U2271 (N_2271,N_2245,N_2218);
and U2272 (N_2272,N_2210,N_2231);
and U2273 (N_2273,N_2233,N_2223);
xor U2274 (N_2274,N_2204,N_2202);
and U2275 (N_2275,N_2232,N_2209);
nor U2276 (N_2276,N_2224,N_2235);
xor U2277 (N_2277,N_2212,N_2244);
nor U2278 (N_2278,N_2231,N_2208);
and U2279 (N_2279,N_2225,N_2220);
or U2280 (N_2280,N_2201,N_2200);
nor U2281 (N_2281,N_2201,N_2220);
and U2282 (N_2282,N_2242,N_2220);
and U2283 (N_2283,N_2249,N_2218);
nor U2284 (N_2284,N_2212,N_2237);
xor U2285 (N_2285,N_2217,N_2212);
nor U2286 (N_2286,N_2230,N_2215);
and U2287 (N_2287,N_2222,N_2221);
xor U2288 (N_2288,N_2221,N_2210);
and U2289 (N_2289,N_2246,N_2234);
nor U2290 (N_2290,N_2244,N_2203);
and U2291 (N_2291,N_2216,N_2240);
nor U2292 (N_2292,N_2231,N_2207);
or U2293 (N_2293,N_2248,N_2234);
xor U2294 (N_2294,N_2239,N_2229);
and U2295 (N_2295,N_2239,N_2223);
or U2296 (N_2296,N_2220,N_2207);
nor U2297 (N_2297,N_2201,N_2245);
and U2298 (N_2298,N_2233,N_2244);
nand U2299 (N_2299,N_2233,N_2241);
nor U2300 (N_2300,N_2264,N_2255);
and U2301 (N_2301,N_2290,N_2288);
nand U2302 (N_2302,N_2254,N_2287);
or U2303 (N_2303,N_2286,N_2279);
and U2304 (N_2304,N_2268,N_2269);
and U2305 (N_2305,N_2270,N_2257);
and U2306 (N_2306,N_2267,N_2261);
nor U2307 (N_2307,N_2262,N_2251);
xor U2308 (N_2308,N_2297,N_2276);
or U2309 (N_2309,N_2273,N_2274);
xnor U2310 (N_2310,N_2252,N_2265);
xor U2311 (N_2311,N_2284,N_2258);
nand U2312 (N_2312,N_2296,N_2282);
and U2313 (N_2313,N_2281,N_2263);
xnor U2314 (N_2314,N_2289,N_2278);
or U2315 (N_2315,N_2298,N_2294);
nor U2316 (N_2316,N_2260,N_2271);
xnor U2317 (N_2317,N_2299,N_2295);
or U2318 (N_2318,N_2250,N_2283);
and U2319 (N_2319,N_2293,N_2272);
or U2320 (N_2320,N_2275,N_2253);
and U2321 (N_2321,N_2266,N_2277);
and U2322 (N_2322,N_2285,N_2292);
nand U2323 (N_2323,N_2291,N_2280);
nand U2324 (N_2324,N_2259,N_2256);
xor U2325 (N_2325,N_2280,N_2250);
or U2326 (N_2326,N_2258,N_2278);
nand U2327 (N_2327,N_2296,N_2276);
or U2328 (N_2328,N_2256,N_2295);
xor U2329 (N_2329,N_2277,N_2296);
nor U2330 (N_2330,N_2251,N_2288);
and U2331 (N_2331,N_2258,N_2267);
nor U2332 (N_2332,N_2290,N_2252);
xnor U2333 (N_2333,N_2280,N_2251);
or U2334 (N_2334,N_2289,N_2275);
xnor U2335 (N_2335,N_2292,N_2271);
xor U2336 (N_2336,N_2255,N_2282);
and U2337 (N_2337,N_2260,N_2255);
and U2338 (N_2338,N_2275,N_2250);
xor U2339 (N_2339,N_2295,N_2289);
and U2340 (N_2340,N_2258,N_2271);
nor U2341 (N_2341,N_2258,N_2257);
nand U2342 (N_2342,N_2265,N_2261);
xor U2343 (N_2343,N_2288,N_2268);
nand U2344 (N_2344,N_2280,N_2261);
xnor U2345 (N_2345,N_2295,N_2262);
nand U2346 (N_2346,N_2284,N_2297);
nand U2347 (N_2347,N_2279,N_2253);
and U2348 (N_2348,N_2257,N_2283);
nand U2349 (N_2349,N_2271,N_2253);
and U2350 (N_2350,N_2347,N_2306);
xnor U2351 (N_2351,N_2312,N_2330);
nand U2352 (N_2352,N_2326,N_2303);
xnor U2353 (N_2353,N_2344,N_2333);
xor U2354 (N_2354,N_2346,N_2323);
nor U2355 (N_2355,N_2318,N_2329);
xor U2356 (N_2356,N_2310,N_2337);
nand U2357 (N_2357,N_2336,N_2327);
nand U2358 (N_2358,N_2335,N_2322);
or U2359 (N_2359,N_2313,N_2301);
nor U2360 (N_2360,N_2345,N_2307);
nor U2361 (N_2361,N_2311,N_2339);
nor U2362 (N_2362,N_2300,N_2308);
nor U2363 (N_2363,N_2325,N_2338);
nor U2364 (N_2364,N_2348,N_2316);
nand U2365 (N_2365,N_2331,N_2317);
nand U2366 (N_2366,N_2349,N_2334);
and U2367 (N_2367,N_2342,N_2320);
and U2368 (N_2368,N_2328,N_2309);
nor U2369 (N_2369,N_2314,N_2321);
nand U2370 (N_2370,N_2305,N_2302);
xor U2371 (N_2371,N_2315,N_2332);
nand U2372 (N_2372,N_2304,N_2319);
and U2373 (N_2373,N_2340,N_2324);
and U2374 (N_2374,N_2343,N_2341);
xor U2375 (N_2375,N_2322,N_2345);
or U2376 (N_2376,N_2348,N_2318);
nor U2377 (N_2377,N_2305,N_2308);
xor U2378 (N_2378,N_2317,N_2302);
xnor U2379 (N_2379,N_2342,N_2307);
nor U2380 (N_2380,N_2309,N_2333);
or U2381 (N_2381,N_2327,N_2345);
nor U2382 (N_2382,N_2342,N_2341);
nand U2383 (N_2383,N_2325,N_2349);
or U2384 (N_2384,N_2330,N_2348);
and U2385 (N_2385,N_2309,N_2342);
xnor U2386 (N_2386,N_2300,N_2327);
and U2387 (N_2387,N_2307,N_2325);
nor U2388 (N_2388,N_2326,N_2330);
nor U2389 (N_2389,N_2304,N_2329);
nor U2390 (N_2390,N_2311,N_2337);
or U2391 (N_2391,N_2316,N_2337);
and U2392 (N_2392,N_2315,N_2310);
xnor U2393 (N_2393,N_2337,N_2341);
and U2394 (N_2394,N_2305,N_2316);
and U2395 (N_2395,N_2307,N_2343);
or U2396 (N_2396,N_2323,N_2317);
xor U2397 (N_2397,N_2320,N_2343);
and U2398 (N_2398,N_2336,N_2314);
nor U2399 (N_2399,N_2307,N_2317);
and U2400 (N_2400,N_2367,N_2386);
xnor U2401 (N_2401,N_2383,N_2380);
or U2402 (N_2402,N_2397,N_2352);
and U2403 (N_2403,N_2377,N_2385);
and U2404 (N_2404,N_2372,N_2362);
xor U2405 (N_2405,N_2370,N_2360);
nand U2406 (N_2406,N_2361,N_2356);
nand U2407 (N_2407,N_2388,N_2378);
nand U2408 (N_2408,N_2376,N_2399);
xor U2409 (N_2409,N_2384,N_2358);
nand U2410 (N_2410,N_2364,N_2351);
nand U2411 (N_2411,N_2390,N_2373);
or U2412 (N_2412,N_2350,N_2357);
nor U2413 (N_2413,N_2374,N_2395);
and U2414 (N_2414,N_2387,N_2363);
nor U2415 (N_2415,N_2359,N_2393);
nand U2416 (N_2416,N_2368,N_2392);
xnor U2417 (N_2417,N_2365,N_2354);
nor U2418 (N_2418,N_2382,N_2355);
xnor U2419 (N_2419,N_2371,N_2389);
or U2420 (N_2420,N_2375,N_2379);
nand U2421 (N_2421,N_2391,N_2394);
and U2422 (N_2422,N_2398,N_2381);
and U2423 (N_2423,N_2366,N_2396);
xor U2424 (N_2424,N_2369,N_2353);
and U2425 (N_2425,N_2391,N_2378);
nor U2426 (N_2426,N_2378,N_2356);
and U2427 (N_2427,N_2379,N_2352);
nor U2428 (N_2428,N_2388,N_2364);
or U2429 (N_2429,N_2396,N_2376);
xor U2430 (N_2430,N_2371,N_2383);
nand U2431 (N_2431,N_2387,N_2367);
nor U2432 (N_2432,N_2390,N_2356);
nand U2433 (N_2433,N_2365,N_2391);
and U2434 (N_2434,N_2367,N_2374);
and U2435 (N_2435,N_2390,N_2395);
nor U2436 (N_2436,N_2396,N_2388);
and U2437 (N_2437,N_2396,N_2373);
nor U2438 (N_2438,N_2386,N_2359);
nor U2439 (N_2439,N_2392,N_2352);
or U2440 (N_2440,N_2363,N_2383);
nor U2441 (N_2441,N_2351,N_2357);
xnor U2442 (N_2442,N_2382,N_2392);
nand U2443 (N_2443,N_2358,N_2392);
and U2444 (N_2444,N_2378,N_2371);
nand U2445 (N_2445,N_2397,N_2398);
nand U2446 (N_2446,N_2393,N_2385);
and U2447 (N_2447,N_2385,N_2361);
or U2448 (N_2448,N_2398,N_2369);
or U2449 (N_2449,N_2357,N_2384);
and U2450 (N_2450,N_2408,N_2405);
or U2451 (N_2451,N_2443,N_2404);
or U2452 (N_2452,N_2400,N_2435);
nand U2453 (N_2453,N_2433,N_2426);
nor U2454 (N_2454,N_2428,N_2422);
and U2455 (N_2455,N_2448,N_2427);
nand U2456 (N_2456,N_2441,N_2401);
or U2457 (N_2457,N_2406,N_2439);
nand U2458 (N_2458,N_2403,N_2434);
nor U2459 (N_2459,N_2449,N_2430);
nor U2460 (N_2460,N_2423,N_2416);
nor U2461 (N_2461,N_2402,N_2420);
and U2462 (N_2462,N_2431,N_2429);
nand U2463 (N_2463,N_2419,N_2444);
nor U2464 (N_2464,N_2438,N_2414);
nor U2465 (N_2465,N_2413,N_2417);
nand U2466 (N_2466,N_2424,N_2436);
and U2467 (N_2467,N_2418,N_2415);
and U2468 (N_2468,N_2447,N_2407);
nor U2469 (N_2469,N_2409,N_2446);
xor U2470 (N_2470,N_2421,N_2437);
or U2471 (N_2471,N_2425,N_2432);
or U2472 (N_2472,N_2442,N_2411);
xor U2473 (N_2473,N_2445,N_2412);
nand U2474 (N_2474,N_2410,N_2440);
and U2475 (N_2475,N_2406,N_2436);
nor U2476 (N_2476,N_2446,N_2400);
nor U2477 (N_2477,N_2406,N_2430);
or U2478 (N_2478,N_2436,N_2430);
nor U2479 (N_2479,N_2447,N_2429);
or U2480 (N_2480,N_2426,N_2411);
nor U2481 (N_2481,N_2440,N_2447);
nand U2482 (N_2482,N_2402,N_2447);
and U2483 (N_2483,N_2438,N_2421);
or U2484 (N_2484,N_2446,N_2429);
nand U2485 (N_2485,N_2432,N_2408);
nor U2486 (N_2486,N_2429,N_2445);
nor U2487 (N_2487,N_2407,N_2406);
nand U2488 (N_2488,N_2416,N_2421);
and U2489 (N_2489,N_2438,N_2445);
nand U2490 (N_2490,N_2444,N_2449);
and U2491 (N_2491,N_2429,N_2427);
and U2492 (N_2492,N_2442,N_2432);
nor U2493 (N_2493,N_2447,N_2433);
or U2494 (N_2494,N_2412,N_2421);
xor U2495 (N_2495,N_2410,N_2419);
and U2496 (N_2496,N_2404,N_2444);
nor U2497 (N_2497,N_2403,N_2425);
nand U2498 (N_2498,N_2425,N_2433);
and U2499 (N_2499,N_2403,N_2444);
and U2500 (N_2500,N_2450,N_2464);
or U2501 (N_2501,N_2490,N_2482);
or U2502 (N_2502,N_2459,N_2476);
nor U2503 (N_2503,N_2455,N_2496);
or U2504 (N_2504,N_2492,N_2454);
xor U2505 (N_2505,N_2456,N_2453);
nand U2506 (N_2506,N_2480,N_2462);
or U2507 (N_2507,N_2484,N_2493);
or U2508 (N_2508,N_2461,N_2474);
and U2509 (N_2509,N_2473,N_2460);
or U2510 (N_2510,N_2471,N_2488);
xnor U2511 (N_2511,N_2497,N_2498);
nor U2512 (N_2512,N_2494,N_2478);
and U2513 (N_2513,N_2466,N_2475);
and U2514 (N_2514,N_2465,N_2452);
nor U2515 (N_2515,N_2463,N_2479);
nand U2516 (N_2516,N_2495,N_2489);
nor U2517 (N_2517,N_2458,N_2483);
nor U2518 (N_2518,N_2499,N_2468);
and U2519 (N_2519,N_2477,N_2457);
xnor U2520 (N_2520,N_2481,N_2472);
and U2521 (N_2521,N_2469,N_2470);
and U2522 (N_2522,N_2451,N_2486);
or U2523 (N_2523,N_2485,N_2487);
xor U2524 (N_2524,N_2467,N_2491);
and U2525 (N_2525,N_2488,N_2480);
and U2526 (N_2526,N_2488,N_2453);
xnor U2527 (N_2527,N_2478,N_2472);
nor U2528 (N_2528,N_2485,N_2499);
xor U2529 (N_2529,N_2470,N_2475);
nand U2530 (N_2530,N_2467,N_2483);
or U2531 (N_2531,N_2461,N_2476);
xnor U2532 (N_2532,N_2483,N_2454);
nor U2533 (N_2533,N_2456,N_2458);
and U2534 (N_2534,N_2454,N_2482);
xnor U2535 (N_2535,N_2465,N_2467);
xnor U2536 (N_2536,N_2460,N_2475);
and U2537 (N_2537,N_2469,N_2466);
or U2538 (N_2538,N_2494,N_2499);
nand U2539 (N_2539,N_2454,N_2488);
nand U2540 (N_2540,N_2488,N_2474);
nand U2541 (N_2541,N_2470,N_2457);
nor U2542 (N_2542,N_2473,N_2498);
nand U2543 (N_2543,N_2454,N_2486);
or U2544 (N_2544,N_2478,N_2453);
nor U2545 (N_2545,N_2466,N_2487);
and U2546 (N_2546,N_2478,N_2498);
nand U2547 (N_2547,N_2492,N_2476);
nor U2548 (N_2548,N_2451,N_2475);
nand U2549 (N_2549,N_2481,N_2454);
nor U2550 (N_2550,N_2517,N_2534);
xnor U2551 (N_2551,N_2508,N_2505);
and U2552 (N_2552,N_2548,N_2513);
nor U2553 (N_2553,N_2542,N_2515);
nand U2554 (N_2554,N_2546,N_2514);
xnor U2555 (N_2555,N_2527,N_2500);
and U2556 (N_2556,N_2511,N_2520);
or U2557 (N_2557,N_2536,N_2545);
nand U2558 (N_2558,N_2543,N_2549);
nand U2559 (N_2559,N_2535,N_2537);
nor U2560 (N_2560,N_2533,N_2510);
xnor U2561 (N_2561,N_2529,N_2522);
or U2562 (N_2562,N_2501,N_2538);
nand U2563 (N_2563,N_2512,N_2528);
nor U2564 (N_2564,N_2507,N_2504);
xor U2565 (N_2565,N_2503,N_2516);
nand U2566 (N_2566,N_2525,N_2526);
and U2567 (N_2567,N_2541,N_2540);
nand U2568 (N_2568,N_2531,N_2519);
and U2569 (N_2569,N_2544,N_2539);
xnor U2570 (N_2570,N_2518,N_2502);
nand U2571 (N_2571,N_2523,N_2521);
xnor U2572 (N_2572,N_2524,N_2506);
and U2573 (N_2573,N_2532,N_2547);
or U2574 (N_2574,N_2509,N_2530);
nor U2575 (N_2575,N_2510,N_2537);
nand U2576 (N_2576,N_2500,N_2531);
and U2577 (N_2577,N_2520,N_2530);
nand U2578 (N_2578,N_2549,N_2502);
and U2579 (N_2579,N_2519,N_2544);
xor U2580 (N_2580,N_2503,N_2513);
nand U2581 (N_2581,N_2517,N_2527);
nand U2582 (N_2582,N_2521,N_2507);
or U2583 (N_2583,N_2533,N_2521);
nand U2584 (N_2584,N_2512,N_2500);
nor U2585 (N_2585,N_2512,N_2510);
and U2586 (N_2586,N_2529,N_2515);
nor U2587 (N_2587,N_2525,N_2541);
xor U2588 (N_2588,N_2547,N_2539);
and U2589 (N_2589,N_2543,N_2500);
xor U2590 (N_2590,N_2544,N_2521);
or U2591 (N_2591,N_2521,N_2548);
nand U2592 (N_2592,N_2545,N_2502);
xor U2593 (N_2593,N_2511,N_2547);
and U2594 (N_2594,N_2538,N_2548);
nand U2595 (N_2595,N_2514,N_2504);
nand U2596 (N_2596,N_2513,N_2502);
nand U2597 (N_2597,N_2538,N_2539);
and U2598 (N_2598,N_2547,N_2540);
and U2599 (N_2599,N_2536,N_2517);
xor U2600 (N_2600,N_2576,N_2574);
or U2601 (N_2601,N_2586,N_2570);
xor U2602 (N_2602,N_2562,N_2557);
or U2603 (N_2603,N_2566,N_2560);
xor U2604 (N_2604,N_2588,N_2572);
nor U2605 (N_2605,N_2550,N_2573);
xor U2606 (N_2606,N_2592,N_2577);
or U2607 (N_2607,N_2590,N_2551);
or U2608 (N_2608,N_2571,N_2591);
or U2609 (N_2609,N_2568,N_2594);
xor U2610 (N_2610,N_2569,N_2564);
or U2611 (N_2611,N_2575,N_2565);
nand U2612 (N_2612,N_2558,N_2579);
xor U2613 (N_2613,N_2597,N_2582);
and U2614 (N_2614,N_2555,N_2599);
and U2615 (N_2615,N_2559,N_2552);
or U2616 (N_2616,N_2583,N_2584);
and U2617 (N_2617,N_2595,N_2598);
xnor U2618 (N_2618,N_2578,N_2593);
xnor U2619 (N_2619,N_2553,N_2556);
nor U2620 (N_2620,N_2580,N_2589);
xor U2621 (N_2621,N_2563,N_2587);
or U2622 (N_2622,N_2561,N_2585);
or U2623 (N_2623,N_2581,N_2596);
nor U2624 (N_2624,N_2554,N_2567);
nand U2625 (N_2625,N_2564,N_2563);
and U2626 (N_2626,N_2551,N_2571);
nand U2627 (N_2627,N_2573,N_2551);
xnor U2628 (N_2628,N_2579,N_2575);
or U2629 (N_2629,N_2555,N_2566);
or U2630 (N_2630,N_2564,N_2580);
and U2631 (N_2631,N_2568,N_2566);
and U2632 (N_2632,N_2592,N_2586);
and U2633 (N_2633,N_2580,N_2578);
or U2634 (N_2634,N_2555,N_2595);
nor U2635 (N_2635,N_2573,N_2565);
nor U2636 (N_2636,N_2567,N_2560);
or U2637 (N_2637,N_2570,N_2587);
and U2638 (N_2638,N_2565,N_2596);
nor U2639 (N_2639,N_2561,N_2587);
xor U2640 (N_2640,N_2584,N_2595);
nand U2641 (N_2641,N_2567,N_2563);
and U2642 (N_2642,N_2571,N_2569);
nand U2643 (N_2643,N_2557,N_2596);
nor U2644 (N_2644,N_2566,N_2565);
and U2645 (N_2645,N_2568,N_2595);
xnor U2646 (N_2646,N_2598,N_2560);
and U2647 (N_2647,N_2574,N_2594);
and U2648 (N_2648,N_2585,N_2587);
nor U2649 (N_2649,N_2594,N_2584);
or U2650 (N_2650,N_2649,N_2628);
or U2651 (N_2651,N_2634,N_2641);
or U2652 (N_2652,N_2601,N_2622);
xor U2653 (N_2653,N_2640,N_2636);
or U2654 (N_2654,N_2603,N_2630);
or U2655 (N_2655,N_2619,N_2617);
and U2656 (N_2656,N_2608,N_2607);
or U2657 (N_2657,N_2631,N_2637);
or U2658 (N_2658,N_2609,N_2638);
xnor U2659 (N_2659,N_2633,N_2611);
and U2660 (N_2660,N_2606,N_2627);
or U2661 (N_2661,N_2621,N_2610);
and U2662 (N_2662,N_2602,N_2626);
or U2663 (N_2663,N_2604,N_2614);
nand U2664 (N_2664,N_2623,N_2629);
nand U2665 (N_2665,N_2645,N_2639);
or U2666 (N_2666,N_2620,N_2632);
or U2667 (N_2667,N_2635,N_2642);
xor U2668 (N_2668,N_2647,N_2643);
xnor U2669 (N_2669,N_2615,N_2644);
xnor U2670 (N_2670,N_2618,N_2616);
xnor U2671 (N_2671,N_2625,N_2600);
nor U2672 (N_2672,N_2612,N_2624);
nor U2673 (N_2673,N_2646,N_2605);
nor U2674 (N_2674,N_2648,N_2613);
and U2675 (N_2675,N_2606,N_2600);
or U2676 (N_2676,N_2612,N_2607);
xor U2677 (N_2677,N_2645,N_2617);
and U2678 (N_2678,N_2613,N_2629);
nand U2679 (N_2679,N_2603,N_2633);
xor U2680 (N_2680,N_2642,N_2640);
or U2681 (N_2681,N_2617,N_2638);
and U2682 (N_2682,N_2623,N_2614);
nand U2683 (N_2683,N_2640,N_2613);
and U2684 (N_2684,N_2633,N_2614);
nor U2685 (N_2685,N_2631,N_2636);
nand U2686 (N_2686,N_2612,N_2645);
and U2687 (N_2687,N_2644,N_2600);
xor U2688 (N_2688,N_2634,N_2627);
xnor U2689 (N_2689,N_2612,N_2631);
nand U2690 (N_2690,N_2615,N_2622);
or U2691 (N_2691,N_2642,N_2630);
and U2692 (N_2692,N_2648,N_2616);
or U2693 (N_2693,N_2644,N_2645);
or U2694 (N_2694,N_2635,N_2600);
or U2695 (N_2695,N_2635,N_2612);
and U2696 (N_2696,N_2629,N_2618);
or U2697 (N_2697,N_2648,N_2621);
or U2698 (N_2698,N_2611,N_2637);
nor U2699 (N_2699,N_2607,N_2643);
nor U2700 (N_2700,N_2688,N_2655);
xnor U2701 (N_2701,N_2694,N_2691);
nand U2702 (N_2702,N_2651,N_2667);
or U2703 (N_2703,N_2693,N_2689);
nand U2704 (N_2704,N_2696,N_2650);
nand U2705 (N_2705,N_2660,N_2673);
nor U2706 (N_2706,N_2664,N_2685);
and U2707 (N_2707,N_2678,N_2668);
and U2708 (N_2708,N_2695,N_2681);
and U2709 (N_2709,N_2699,N_2676);
nand U2710 (N_2710,N_2677,N_2687);
xor U2711 (N_2711,N_2690,N_2663);
or U2712 (N_2712,N_2659,N_2697);
or U2713 (N_2713,N_2698,N_2675);
or U2714 (N_2714,N_2652,N_2665);
nand U2715 (N_2715,N_2662,N_2672);
and U2716 (N_2716,N_2666,N_2686);
or U2717 (N_2717,N_2679,N_2684);
and U2718 (N_2718,N_2669,N_2692);
nand U2719 (N_2719,N_2682,N_2657);
nor U2720 (N_2720,N_2661,N_2670);
and U2721 (N_2721,N_2680,N_2654);
or U2722 (N_2722,N_2658,N_2671);
nor U2723 (N_2723,N_2653,N_2656);
nand U2724 (N_2724,N_2683,N_2674);
and U2725 (N_2725,N_2667,N_2673);
nor U2726 (N_2726,N_2662,N_2661);
and U2727 (N_2727,N_2667,N_2685);
nor U2728 (N_2728,N_2651,N_2683);
or U2729 (N_2729,N_2690,N_2692);
xnor U2730 (N_2730,N_2651,N_2681);
and U2731 (N_2731,N_2679,N_2652);
and U2732 (N_2732,N_2663,N_2692);
nor U2733 (N_2733,N_2690,N_2655);
nand U2734 (N_2734,N_2650,N_2658);
nor U2735 (N_2735,N_2699,N_2671);
nand U2736 (N_2736,N_2672,N_2686);
nand U2737 (N_2737,N_2691,N_2665);
or U2738 (N_2738,N_2651,N_2693);
nand U2739 (N_2739,N_2698,N_2677);
nor U2740 (N_2740,N_2651,N_2695);
and U2741 (N_2741,N_2670,N_2681);
and U2742 (N_2742,N_2689,N_2663);
and U2743 (N_2743,N_2675,N_2659);
or U2744 (N_2744,N_2670,N_2680);
xnor U2745 (N_2745,N_2677,N_2665);
nand U2746 (N_2746,N_2697,N_2684);
xnor U2747 (N_2747,N_2697,N_2670);
xnor U2748 (N_2748,N_2694,N_2654);
nor U2749 (N_2749,N_2694,N_2693);
xor U2750 (N_2750,N_2708,N_2739);
and U2751 (N_2751,N_2736,N_2702);
nand U2752 (N_2752,N_2720,N_2724);
xnor U2753 (N_2753,N_2743,N_2718);
nand U2754 (N_2754,N_2716,N_2712);
xnor U2755 (N_2755,N_2740,N_2734);
or U2756 (N_2756,N_2721,N_2749);
xnor U2757 (N_2757,N_2713,N_2730);
nand U2758 (N_2758,N_2703,N_2711);
and U2759 (N_2759,N_2729,N_2727);
nand U2760 (N_2760,N_2714,N_2735);
or U2761 (N_2761,N_2726,N_2733);
and U2762 (N_2762,N_2748,N_2705);
xnor U2763 (N_2763,N_2744,N_2737);
xor U2764 (N_2764,N_2728,N_2745);
nand U2765 (N_2765,N_2731,N_2710);
or U2766 (N_2766,N_2715,N_2723);
and U2767 (N_2767,N_2700,N_2725);
and U2768 (N_2768,N_2738,N_2741);
nor U2769 (N_2769,N_2709,N_2701);
or U2770 (N_2770,N_2722,N_2717);
xnor U2771 (N_2771,N_2719,N_2747);
and U2772 (N_2772,N_2732,N_2707);
xor U2773 (N_2773,N_2704,N_2706);
nor U2774 (N_2774,N_2742,N_2746);
nor U2775 (N_2775,N_2739,N_2744);
nor U2776 (N_2776,N_2726,N_2713);
and U2777 (N_2777,N_2739,N_2748);
xnor U2778 (N_2778,N_2743,N_2719);
and U2779 (N_2779,N_2709,N_2730);
xor U2780 (N_2780,N_2717,N_2701);
nand U2781 (N_2781,N_2730,N_2725);
nand U2782 (N_2782,N_2736,N_2720);
or U2783 (N_2783,N_2732,N_2704);
nor U2784 (N_2784,N_2702,N_2737);
xor U2785 (N_2785,N_2709,N_2728);
nor U2786 (N_2786,N_2708,N_2720);
nor U2787 (N_2787,N_2727,N_2740);
nand U2788 (N_2788,N_2708,N_2722);
nor U2789 (N_2789,N_2701,N_2702);
nor U2790 (N_2790,N_2742,N_2704);
nand U2791 (N_2791,N_2702,N_2705);
xnor U2792 (N_2792,N_2723,N_2720);
nor U2793 (N_2793,N_2714,N_2726);
xor U2794 (N_2794,N_2700,N_2721);
and U2795 (N_2795,N_2702,N_2745);
and U2796 (N_2796,N_2724,N_2739);
xor U2797 (N_2797,N_2739,N_2731);
or U2798 (N_2798,N_2734,N_2723);
and U2799 (N_2799,N_2718,N_2747);
nor U2800 (N_2800,N_2797,N_2766);
xor U2801 (N_2801,N_2762,N_2784);
and U2802 (N_2802,N_2796,N_2793);
xor U2803 (N_2803,N_2755,N_2776);
or U2804 (N_2804,N_2798,N_2787);
xnor U2805 (N_2805,N_2783,N_2778);
xnor U2806 (N_2806,N_2770,N_2779);
nand U2807 (N_2807,N_2794,N_2788);
nor U2808 (N_2808,N_2790,N_2756);
xor U2809 (N_2809,N_2752,N_2795);
nand U2810 (N_2810,N_2773,N_2754);
or U2811 (N_2811,N_2763,N_2758);
nor U2812 (N_2812,N_2774,N_2780);
xnor U2813 (N_2813,N_2789,N_2791);
and U2814 (N_2814,N_2759,N_2753);
nand U2815 (N_2815,N_2750,N_2751);
nand U2816 (N_2816,N_2757,N_2760);
or U2817 (N_2817,N_2769,N_2799);
nor U2818 (N_2818,N_2764,N_2761);
xnor U2819 (N_2819,N_2767,N_2782);
nand U2820 (N_2820,N_2765,N_2771);
or U2821 (N_2821,N_2777,N_2792);
xnor U2822 (N_2822,N_2775,N_2768);
nor U2823 (N_2823,N_2785,N_2786);
xor U2824 (N_2824,N_2781,N_2772);
or U2825 (N_2825,N_2753,N_2763);
xnor U2826 (N_2826,N_2761,N_2784);
nor U2827 (N_2827,N_2788,N_2785);
or U2828 (N_2828,N_2754,N_2784);
nor U2829 (N_2829,N_2776,N_2757);
nor U2830 (N_2830,N_2756,N_2796);
nand U2831 (N_2831,N_2775,N_2750);
or U2832 (N_2832,N_2786,N_2794);
nand U2833 (N_2833,N_2799,N_2756);
nor U2834 (N_2834,N_2758,N_2768);
nand U2835 (N_2835,N_2797,N_2769);
nor U2836 (N_2836,N_2757,N_2755);
xor U2837 (N_2837,N_2785,N_2765);
xnor U2838 (N_2838,N_2763,N_2780);
and U2839 (N_2839,N_2752,N_2764);
xor U2840 (N_2840,N_2795,N_2783);
and U2841 (N_2841,N_2765,N_2783);
xor U2842 (N_2842,N_2779,N_2766);
xnor U2843 (N_2843,N_2786,N_2751);
nand U2844 (N_2844,N_2752,N_2757);
or U2845 (N_2845,N_2792,N_2750);
nor U2846 (N_2846,N_2767,N_2757);
nand U2847 (N_2847,N_2774,N_2755);
nand U2848 (N_2848,N_2756,N_2792);
and U2849 (N_2849,N_2768,N_2770);
and U2850 (N_2850,N_2831,N_2842);
and U2851 (N_2851,N_2833,N_2813);
xnor U2852 (N_2852,N_2809,N_2834);
nor U2853 (N_2853,N_2816,N_2822);
nor U2854 (N_2854,N_2812,N_2808);
and U2855 (N_2855,N_2837,N_2814);
nand U2856 (N_2856,N_2828,N_2835);
or U2857 (N_2857,N_2817,N_2838);
nor U2858 (N_2858,N_2801,N_2830);
nor U2859 (N_2859,N_2823,N_2843);
nor U2860 (N_2860,N_2846,N_2802);
nor U2861 (N_2861,N_2847,N_2849);
or U2862 (N_2862,N_2811,N_2824);
nand U2863 (N_2863,N_2803,N_2804);
nor U2864 (N_2864,N_2832,N_2848);
and U2865 (N_2865,N_2826,N_2821);
xnor U2866 (N_2866,N_2839,N_2820);
and U2867 (N_2867,N_2841,N_2807);
nor U2868 (N_2868,N_2806,N_2819);
and U2869 (N_2869,N_2845,N_2805);
and U2870 (N_2870,N_2840,N_2836);
and U2871 (N_2871,N_2825,N_2800);
and U2872 (N_2872,N_2829,N_2810);
nand U2873 (N_2873,N_2827,N_2844);
and U2874 (N_2874,N_2815,N_2818);
or U2875 (N_2875,N_2813,N_2838);
nor U2876 (N_2876,N_2833,N_2825);
xnor U2877 (N_2877,N_2841,N_2810);
nand U2878 (N_2878,N_2801,N_2815);
xnor U2879 (N_2879,N_2846,N_2801);
nand U2880 (N_2880,N_2814,N_2832);
xnor U2881 (N_2881,N_2814,N_2803);
and U2882 (N_2882,N_2847,N_2803);
and U2883 (N_2883,N_2825,N_2841);
nor U2884 (N_2884,N_2849,N_2826);
nand U2885 (N_2885,N_2833,N_2803);
or U2886 (N_2886,N_2807,N_2806);
and U2887 (N_2887,N_2848,N_2829);
or U2888 (N_2888,N_2809,N_2839);
or U2889 (N_2889,N_2849,N_2835);
and U2890 (N_2890,N_2812,N_2818);
nor U2891 (N_2891,N_2804,N_2839);
or U2892 (N_2892,N_2808,N_2821);
nand U2893 (N_2893,N_2805,N_2816);
nand U2894 (N_2894,N_2832,N_2833);
and U2895 (N_2895,N_2836,N_2830);
and U2896 (N_2896,N_2835,N_2831);
and U2897 (N_2897,N_2801,N_2844);
nor U2898 (N_2898,N_2806,N_2817);
or U2899 (N_2899,N_2834,N_2817);
nor U2900 (N_2900,N_2882,N_2895);
or U2901 (N_2901,N_2857,N_2890);
nor U2902 (N_2902,N_2897,N_2883);
xnor U2903 (N_2903,N_2861,N_2887);
and U2904 (N_2904,N_2863,N_2893);
or U2905 (N_2905,N_2872,N_2871);
nand U2906 (N_2906,N_2858,N_2892);
xnor U2907 (N_2907,N_2888,N_2851);
xnor U2908 (N_2908,N_2884,N_2870);
and U2909 (N_2909,N_2880,N_2852);
xor U2910 (N_2910,N_2874,N_2868);
nand U2911 (N_2911,N_2864,N_2876);
xnor U2912 (N_2912,N_2860,N_2854);
xnor U2913 (N_2913,N_2862,N_2875);
xor U2914 (N_2914,N_2896,N_2885);
and U2915 (N_2915,N_2886,N_2856);
or U2916 (N_2916,N_2873,N_2898);
and U2917 (N_2917,N_2878,N_2881);
or U2918 (N_2918,N_2891,N_2855);
or U2919 (N_2919,N_2879,N_2866);
and U2920 (N_2920,N_2865,N_2894);
xnor U2921 (N_2921,N_2853,N_2859);
xor U2922 (N_2922,N_2850,N_2899);
or U2923 (N_2923,N_2869,N_2867);
nand U2924 (N_2924,N_2877,N_2889);
xnor U2925 (N_2925,N_2874,N_2857);
and U2926 (N_2926,N_2858,N_2856);
nand U2927 (N_2927,N_2885,N_2877);
or U2928 (N_2928,N_2860,N_2868);
and U2929 (N_2929,N_2863,N_2898);
and U2930 (N_2930,N_2861,N_2883);
xnor U2931 (N_2931,N_2893,N_2870);
nor U2932 (N_2932,N_2868,N_2857);
nor U2933 (N_2933,N_2897,N_2891);
nand U2934 (N_2934,N_2870,N_2888);
or U2935 (N_2935,N_2873,N_2856);
nand U2936 (N_2936,N_2889,N_2899);
and U2937 (N_2937,N_2863,N_2864);
or U2938 (N_2938,N_2879,N_2882);
xnor U2939 (N_2939,N_2887,N_2894);
nand U2940 (N_2940,N_2856,N_2894);
or U2941 (N_2941,N_2859,N_2897);
and U2942 (N_2942,N_2863,N_2862);
nor U2943 (N_2943,N_2857,N_2862);
nor U2944 (N_2944,N_2865,N_2863);
xor U2945 (N_2945,N_2888,N_2866);
and U2946 (N_2946,N_2861,N_2870);
nor U2947 (N_2947,N_2886,N_2897);
and U2948 (N_2948,N_2888,N_2875);
nor U2949 (N_2949,N_2856,N_2890);
nor U2950 (N_2950,N_2916,N_2911);
nor U2951 (N_2951,N_2929,N_2933);
nand U2952 (N_2952,N_2936,N_2940);
nor U2953 (N_2953,N_2921,N_2946);
or U2954 (N_2954,N_2923,N_2919);
xor U2955 (N_2955,N_2948,N_2926);
nand U2956 (N_2956,N_2942,N_2941);
nor U2957 (N_2957,N_2931,N_2901);
nand U2958 (N_2958,N_2938,N_2932);
nor U2959 (N_2959,N_2918,N_2900);
nor U2960 (N_2960,N_2943,N_2922);
and U2961 (N_2961,N_2908,N_2904);
nor U2962 (N_2962,N_2925,N_2905);
nor U2963 (N_2963,N_2947,N_2920);
nand U2964 (N_2964,N_2906,N_2934);
or U2965 (N_2965,N_2910,N_2928);
nor U2966 (N_2966,N_2903,N_2909);
or U2967 (N_2967,N_2902,N_2949);
nor U2968 (N_2968,N_2937,N_2917);
xnor U2969 (N_2969,N_2924,N_2914);
nor U2970 (N_2970,N_2944,N_2913);
and U2971 (N_2971,N_2915,N_2927);
nand U2972 (N_2972,N_2907,N_2912);
nand U2973 (N_2973,N_2935,N_2930);
or U2974 (N_2974,N_2939,N_2945);
nor U2975 (N_2975,N_2926,N_2924);
nor U2976 (N_2976,N_2941,N_2920);
xnor U2977 (N_2977,N_2947,N_2929);
xor U2978 (N_2978,N_2928,N_2902);
nor U2979 (N_2979,N_2906,N_2940);
nand U2980 (N_2980,N_2905,N_2938);
xnor U2981 (N_2981,N_2923,N_2941);
or U2982 (N_2982,N_2941,N_2931);
nor U2983 (N_2983,N_2928,N_2946);
and U2984 (N_2984,N_2931,N_2922);
xnor U2985 (N_2985,N_2946,N_2901);
xor U2986 (N_2986,N_2936,N_2948);
and U2987 (N_2987,N_2919,N_2909);
nor U2988 (N_2988,N_2948,N_2942);
nor U2989 (N_2989,N_2908,N_2937);
nand U2990 (N_2990,N_2903,N_2938);
and U2991 (N_2991,N_2904,N_2914);
xnor U2992 (N_2992,N_2945,N_2938);
nand U2993 (N_2993,N_2932,N_2927);
nor U2994 (N_2994,N_2911,N_2949);
nand U2995 (N_2995,N_2916,N_2917);
or U2996 (N_2996,N_2904,N_2939);
nor U2997 (N_2997,N_2946,N_2906);
and U2998 (N_2998,N_2943,N_2900);
nand U2999 (N_2999,N_2919,N_2927);
xnor UO_0 (O_0,N_2996,N_2960);
xor UO_1 (O_1,N_2988,N_2974);
or UO_2 (O_2,N_2993,N_2992);
xor UO_3 (O_3,N_2965,N_2971);
or UO_4 (O_4,N_2990,N_2977);
nor UO_5 (O_5,N_2950,N_2966);
xor UO_6 (O_6,N_2964,N_2987);
nor UO_7 (O_7,N_2978,N_2963);
or UO_8 (O_8,N_2957,N_2983);
nor UO_9 (O_9,N_2967,N_2961);
nor UO_10 (O_10,N_2998,N_2997);
nor UO_11 (O_11,N_2972,N_2975);
and UO_12 (O_12,N_2968,N_2958);
or UO_13 (O_13,N_2991,N_2969);
nand UO_14 (O_14,N_2986,N_2973);
nand UO_15 (O_15,N_2970,N_2979);
nand UO_16 (O_16,N_2953,N_2984);
or UO_17 (O_17,N_2995,N_2952);
or UO_18 (O_18,N_2981,N_2985);
nand UO_19 (O_19,N_2955,N_2999);
nor UO_20 (O_20,N_2951,N_2954);
nand UO_21 (O_21,N_2989,N_2980);
and UO_22 (O_22,N_2994,N_2962);
xor UO_23 (O_23,N_2956,N_2982);
or UO_24 (O_24,N_2976,N_2959);
and UO_25 (O_25,N_2988,N_2971);
nand UO_26 (O_26,N_2956,N_2969);
xnor UO_27 (O_27,N_2984,N_2965);
and UO_28 (O_28,N_2973,N_2965);
or UO_29 (O_29,N_2957,N_2979);
nor UO_30 (O_30,N_2950,N_2975);
and UO_31 (O_31,N_2964,N_2995);
nand UO_32 (O_32,N_2968,N_2964);
xor UO_33 (O_33,N_2957,N_2954);
or UO_34 (O_34,N_2990,N_2981);
or UO_35 (O_35,N_2951,N_2977);
nor UO_36 (O_36,N_2970,N_2951);
nand UO_37 (O_37,N_2970,N_2988);
xor UO_38 (O_38,N_2980,N_2963);
nor UO_39 (O_39,N_2965,N_2983);
nand UO_40 (O_40,N_2972,N_2998);
nor UO_41 (O_41,N_2987,N_2979);
and UO_42 (O_42,N_2950,N_2972);
nand UO_43 (O_43,N_2966,N_2967);
nand UO_44 (O_44,N_2966,N_2988);
nor UO_45 (O_45,N_2984,N_2967);
and UO_46 (O_46,N_2976,N_2986);
nor UO_47 (O_47,N_2985,N_2998);
nand UO_48 (O_48,N_2994,N_2950);
and UO_49 (O_49,N_2977,N_2982);
nor UO_50 (O_50,N_2973,N_2987);
and UO_51 (O_51,N_2987,N_2965);
and UO_52 (O_52,N_2966,N_2983);
nor UO_53 (O_53,N_2986,N_2967);
nor UO_54 (O_54,N_2972,N_2982);
or UO_55 (O_55,N_2993,N_2978);
or UO_56 (O_56,N_2970,N_2972);
nand UO_57 (O_57,N_2975,N_2953);
xor UO_58 (O_58,N_2976,N_2970);
nor UO_59 (O_59,N_2960,N_2986);
nor UO_60 (O_60,N_2955,N_2971);
nand UO_61 (O_61,N_2983,N_2961);
nor UO_62 (O_62,N_2956,N_2998);
and UO_63 (O_63,N_2958,N_2982);
nand UO_64 (O_64,N_2953,N_2971);
nor UO_65 (O_65,N_2959,N_2999);
nand UO_66 (O_66,N_2960,N_2992);
nor UO_67 (O_67,N_2972,N_2957);
and UO_68 (O_68,N_2976,N_2987);
nand UO_69 (O_69,N_2976,N_2958);
and UO_70 (O_70,N_2988,N_2990);
nand UO_71 (O_71,N_2981,N_2957);
nand UO_72 (O_72,N_2960,N_2962);
xor UO_73 (O_73,N_2979,N_2980);
or UO_74 (O_74,N_2968,N_2980);
nor UO_75 (O_75,N_2995,N_2986);
xnor UO_76 (O_76,N_2989,N_2997);
nand UO_77 (O_77,N_2960,N_2989);
nand UO_78 (O_78,N_2980,N_2996);
and UO_79 (O_79,N_2966,N_2965);
and UO_80 (O_80,N_2967,N_2975);
or UO_81 (O_81,N_2997,N_2966);
or UO_82 (O_82,N_2993,N_2953);
xor UO_83 (O_83,N_2960,N_2961);
or UO_84 (O_84,N_2966,N_2985);
nor UO_85 (O_85,N_2990,N_2965);
or UO_86 (O_86,N_2972,N_2973);
and UO_87 (O_87,N_2984,N_2968);
nand UO_88 (O_88,N_2999,N_2964);
and UO_89 (O_89,N_2976,N_2952);
xor UO_90 (O_90,N_2988,N_2987);
and UO_91 (O_91,N_2968,N_2983);
nor UO_92 (O_92,N_2957,N_2989);
nand UO_93 (O_93,N_2973,N_2958);
and UO_94 (O_94,N_2966,N_2993);
and UO_95 (O_95,N_2963,N_2964);
and UO_96 (O_96,N_2957,N_2980);
nand UO_97 (O_97,N_2999,N_2975);
xor UO_98 (O_98,N_2973,N_2952);
xnor UO_99 (O_99,N_2965,N_2996);
xnor UO_100 (O_100,N_2971,N_2991);
nor UO_101 (O_101,N_2988,N_2995);
or UO_102 (O_102,N_2973,N_2992);
nor UO_103 (O_103,N_2950,N_2970);
and UO_104 (O_104,N_2964,N_2991);
or UO_105 (O_105,N_2995,N_2960);
and UO_106 (O_106,N_2980,N_2978);
and UO_107 (O_107,N_2989,N_2953);
and UO_108 (O_108,N_2982,N_2957);
and UO_109 (O_109,N_2981,N_2997);
or UO_110 (O_110,N_2965,N_2963);
or UO_111 (O_111,N_2971,N_2996);
nor UO_112 (O_112,N_2967,N_2969);
and UO_113 (O_113,N_2972,N_2997);
nand UO_114 (O_114,N_2964,N_2988);
nor UO_115 (O_115,N_2970,N_2978);
nand UO_116 (O_116,N_2952,N_2984);
and UO_117 (O_117,N_2962,N_2973);
or UO_118 (O_118,N_2979,N_2996);
nand UO_119 (O_119,N_2987,N_2984);
nand UO_120 (O_120,N_2979,N_2964);
xor UO_121 (O_121,N_2971,N_2983);
and UO_122 (O_122,N_2962,N_2952);
nor UO_123 (O_123,N_2997,N_2959);
and UO_124 (O_124,N_2995,N_2968);
nor UO_125 (O_125,N_2981,N_2970);
xor UO_126 (O_126,N_2963,N_2987);
or UO_127 (O_127,N_2969,N_2963);
and UO_128 (O_128,N_2994,N_2986);
nand UO_129 (O_129,N_2962,N_2963);
nand UO_130 (O_130,N_2977,N_2964);
nand UO_131 (O_131,N_2961,N_2959);
nand UO_132 (O_132,N_2982,N_2976);
nand UO_133 (O_133,N_2953,N_2954);
and UO_134 (O_134,N_2959,N_2985);
nand UO_135 (O_135,N_2990,N_2951);
or UO_136 (O_136,N_2973,N_2977);
xor UO_137 (O_137,N_2961,N_2974);
or UO_138 (O_138,N_2977,N_2968);
nand UO_139 (O_139,N_2969,N_2966);
or UO_140 (O_140,N_2962,N_2954);
or UO_141 (O_141,N_2956,N_2965);
or UO_142 (O_142,N_2999,N_2987);
or UO_143 (O_143,N_2959,N_2956);
or UO_144 (O_144,N_2998,N_2983);
and UO_145 (O_145,N_2970,N_2995);
nand UO_146 (O_146,N_2954,N_2983);
xnor UO_147 (O_147,N_2971,N_2963);
nand UO_148 (O_148,N_2977,N_2963);
nand UO_149 (O_149,N_2999,N_2958);
xor UO_150 (O_150,N_2984,N_2982);
nand UO_151 (O_151,N_2982,N_2988);
nor UO_152 (O_152,N_2994,N_2980);
or UO_153 (O_153,N_2956,N_2957);
xor UO_154 (O_154,N_2961,N_2980);
or UO_155 (O_155,N_2960,N_2965);
and UO_156 (O_156,N_2975,N_2987);
or UO_157 (O_157,N_2963,N_2990);
nand UO_158 (O_158,N_2955,N_2962);
or UO_159 (O_159,N_2970,N_2993);
nand UO_160 (O_160,N_2955,N_2952);
nor UO_161 (O_161,N_2984,N_2956);
or UO_162 (O_162,N_2976,N_2974);
and UO_163 (O_163,N_2957,N_2975);
and UO_164 (O_164,N_2956,N_2997);
or UO_165 (O_165,N_2968,N_2969);
xor UO_166 (O_166,N_2984,N_2988);
nor UO_167 (O_167,N_2998,N_2964);
and UO_168 (O_168,N_2990,N_2966);
and UO_169 (O_169,N_2998,N_2959);
nor UO_170 (O_170,N_2972,N_2988);
nor UO_171 (O_171,N_2976,N_2962);
nor UO_172 (O_172,N_2995,N_2953);
nor UO_173 (O_173,N_2957,N_2998);
xor UO_174 (O_174,N_2974,N_2979);
and UO_175 (O_175,N_2977,N_2989);
nand UO_176 (O_176,N_2952,N_2980);
nor UO_177 (O_177,N_2973,N_2985);
xnor UO_178 (O_178,N_2972,N_2995);
nand UO_179 (O_179,N_2990,N_2961);
nand UO_180 (O_180,N_2971,N_2993);
and UO_181 (O_181,N_2997,N_2975);
and UO_182 (O_182,N_2979,N_2966);
and UO_183 (O_183,N_2994,N_2997);
or UO_184 (O_184,N_2990,N_2958);
or UO_185 (O_185,N_2971,N_2970);
nand UO_186 (O_186,N_2979,N_2999);
or UO_187 (O_187,N_2982,N_2987);
nand UO_188 (O_188,N_2979,N_2955);
nand UO_189 (O_189,N_2986,N_2961);
nor UO_190 (O_190,N_2970,N_2977);
and UO_191 (O_191,N_2971,N_2966);
nand UO_192 (O_192,N_2995,N_2950);
xnor UO_193 (O_193,N_2984,N_2986);
nand UO_194 (O_194,N_2966,N_2992);
nand UO_195 (O_195,N_2972,N_2968);
xnor UO_196 (O_196,N_2967,N_2991);
or UO_197 (O_197,N_2998,N_2960);
xnor UO_198 (O_198,N_2955,N_2975);
xnor UO_199 (O_199,N_2980,N_2992);
nor UO_200 (O_200,N_2984,N_2991);
nor UO_201 (O_201,N_2970,N_2968);
and UO_202 (O_202,N_2965,N_2999);
nor UO_203 (O_203,N_2994,N_2965);
or UO_204 (O_204,N_2977,N_2967);
and UO_205 (O_205,N_2954,N_2991);
and UO_206 (O_206,N_2958,N_2956);
or UO_207 (O_207,N_2969,N_2985);
xnor UO_208 (O_208,N_2968,N_2979);
nor UO_209 (O_209,N_2983,N_2967);
xnor UO_210 (O_210,N_2979,N_2977);
nand UO_211 (O_211,N_2993,N_2951);
and UO_212 (O_212,N_2996,N_2974);
nor UO_213 (O_213,N_2959,N_2968);
nor UO_214 (O_214,N_2966,N_2975);
nand UO_215 (O_215,N_2980,N_2970);
and UO_216 (O_216,N_2981,N_2951);
and UO_217 (O_217,N_2961,N_2968);
xor UO_218 (O_218,N_2959,N_2951);
nor UO_219 (O_219,N_2951,N_2976);
nand UO_220 (O_220,N_2956,N_2953);
xor UO_221 (O_221,N_2961,N_2965);
and UO_222 (O_222,N_2985,N_2992);
nand UO_223 (O_223,N_2981,N_2968);
nor UO_224 (O_224,N_2992,N_2964);
nand UO_225 (O_225,N_2963,N_2994);
nand UO_226 (O_226,N_2989,N_2987);
nor UO_227 (O_227,N_2967,N_2952);
and UO_228 (O_228,N_2973,N_2969);
nand UO_229 (O_229,N_2958,N_2989);
or UO_230 (O_230,N_2964,N_2996);
xnor UO_231 (O_231,N_2986,N_2978);
and UO_232 (O_232,N_2950,N_2957);
xnor UO_233 (O_233,N_2999,N_2988);
xor UO_234 (O_234,N_2967,N_2950);
nand UO_235 (O_235,N_2987,N_2983);
or UO_236 (O_236,N_2996,N_2983);
nor UO_237 (O_237,N_2986,N_2982);
xnor UO_238 (O_238,N_2960,N_2984);
nor UO_239 (O_239,N_2957,N_2990);
xnor UO_240 (O_240,N_2954,N_2963);
xnor UO_241 (O_241,N_2965,N_2989);
nand UO_242 (O_242,N_2976,N_2971);
and UO_243 (O_243,N_2959,N_2986);
nand UO_244 (O_244,N_2995,N_2979);
or UO_245 (O_245,N_2955,N_2992);
and UO_246 (O_246,N_2951,N_2997);
nand UO_247 (O_247,N_2965,N_2955);
nand UO_248 (O_248,N_2973,N_2976);
or UO_249 (O_249,N_2974,N_2987);
nand UO_250 (O_250,N_2974,N_2959);
and UO_251 (O_251,N_2995,N_2999);
xor UO_252 (O_252,N_2950,N_2955);
and UO_253 (O_253,N_2991,N_2975);
nand UO_254 (O_254,N_2952,N_2961);
nand UO_255 (O_255,N_2998,N_2978);
nand UO_256 (O_256,N_2987,N_2997);
xnor UO_257 (O_257,N_2972,N_2959);
nand UO_258 (O_258,N_2960,N_2959);
nor UO_259 (O_259,N_2970,N_2986);
xnor UO_260 (O_260,N_2990,N_2975);
nand UO_261 (O_261,N_2981,N_2965);
or UO_262 (O_262,N_2953,N_2998);
xor UO_263 (O_263,N_2984,N_2973);
nor UO_264 (O_264,N_2973,N_2953);
nor UO_265 (O_265,N_2951,N_2987);
and UO_266 (O_266,N_2987,N_2977);
nand UO_267 (O_267,N_2971,N_2972);
or UO_268 (O_268,N_2969,N_2959);
nor UO_269 (O_269,N_2996,N_2950);
nor UO_270 (O_270,N_2994,N_2977);
or UO_271 (O_271,N_2984,N_2970);
or UO_272 (O_272,N_2967,N_2972);
nor UO_273 (O_273,N_2977,N_2993);
xor UO_274 (O_274,N_2973,N_2975);
xnor UO_275 (O_275,N_2958,N_2963);
nor UO_276 (O_276,N_2997,N_2961);
xnor UO_277 (O_277,N_2970,N_2956);
nand UO_278 (O_278,N_2971,N_2974);
nand UO_279 (O_279,N_2965,N_2995);
nand UO_280 (O_280,N_2978,N_2950);
nand UO_281 (O_281,N_2950,N_2980);
and UO_282 (O_282,N_2975,N_2962);
or UO_283 (O_283,N_2997,N_2990);
xnor UO_284 (O_284,N_2998,N_2999);
xor UO_285 (O_285,N_2993,N_2984);
or UO_286 (O_286,N_2958,N_2964);
nand UO_287 (O_287,N_2955,N_2997);
nor UO_288 (O_288,N_2954,N_2995);
or UO_289 (O_289,N_2962,N_2999);
nand UO_290 (O_290,N_2970,N_2983);
nor UO_291 (O_291,N_2990,N_2964);
and UO_292 (O_292,N_2952,N_2994);
nor UO_293 (O_293,N_2996,N_2958);
and UO_294 (O_294,N_2978,N_2965);
xor UO_295 (O_295,N_2971,N_2957);
nand UO_296 (O_296,N_2988,N_2973);
and UO_297 (O_297,N_2965,N_2950);
or UO_298 (O_298,N_2986,N_2992);
nor UO_299 (O_299,N_2986,N_2979);
and UO_300 (O_300,N_2967,N_2956);
xnor UO_301 (O_301,N_2991,N_2961);
nor UO_302 (O_302,N_2967,N_2979);
and UO_303 (O_303,N_2964,N_2972);
or UO_304 (O_304,N_2973,N_2982);
or UO_305 (O_305,N_2955,N_2968);
nor UO_306 (O_306,N_2969,N_2954);
xor UO_307 (O_307,N_2998,N_2951);
or UO_308 (O_308,N_2998,N_2955);
nand UO_309 (O_309,N_2980,N_2960);
nand UO_310 (O_310,N_2961,N_2989);
nor UO_311 (O_311,N_2998,N_2967);
and UO_312 (O_312,N_2984,N_2955);
or UO_313 (O_313,N_2995,N_2981);
nor UO_314 (O_314,N_2984,N_2997);
xor UO_315 (O_315,N_2991,N_2973);
nor UO_316 (O_316,N_2984,N_2985);
nand UO_317 (O_317,N_2992,N_2953);
nor UO_318 (O_318,N_2988,N_2968);
or UO_319 (O_319,N_2997,N_2967);
and UO_320 (O_320,N_2959,N_2979);
xnor UO_321 (O_321,N_2955,N_2980);
and UO_322 (O_322,N_2957,N_2973);
nand UO_323 (O_323,N_2956,N_2968);
and UO_324 (O_324,N_2978,N_2996);
xor UO_325 (O_325,N_2958,N_2991);
xnor UO_326 (O_326,N_2950,N_2997);
and UO_327 (O_327,N_2975,N_2976);
nand UO_328 (O_328,N_2956,N_2992);
nand UO_329 (O_329,N_2950,N_2969);
or UO_330 (O_330,N_2966,N_2976);
nor UO_331 (O_331,N_2988,N_2986);
and UO_332 (O_332,N_2966,N_2958);
xnor UO_333 (O_333,N_2979,N_2983);
nor UO_334 (O_334,N_2956,N_2952);
and UO_335 (O_335,N_2993,N_2969);
nor UO_336 (O_336,N_2969,N_2953);
nand UO_337 (O_337,N_2979,N_2984);
nand UO_338 (O_338,N_2975,N_2959);
or UO_339 (O_339,N_2961,N_2987);
and UO_340 (O_340,N_2991,N_2950);
nor UO_341 (O_341,N_2957,N_2997);
nand UO_342 (O_342,N_2974,N_2980);
xnor UO_343 (O_343,N_2974,N_2986);
or UO_344 (O_344,N_2963,N_2999);
nor UO_345 (O_345,N_2962,N_2982);
xor UO_346 (O_346,N_2955,N_2961);
xnor UO_347 (O_347,N_2986,N_2966);
nand UO_348 (O_348,N_2969,N_2999);
nor UO_349 (O_349,N_2974,N_2990);
xor UO_350 (O_350,N_2957,N_2958);
nand UO_351 (O_351,N_2957,N_2967);
nand UO_352 (O_352,N_2963,N_2951);
and UO_353 (O_353,N_2951,N_2996);
xor UO_354 (O_354,N_2977,N_2985);
nand UO_355 (O_355,N_2953,N_2991);
or UO_356 (O_356,N_2993,N_2961);
nor UO_357 (O_357,N_2980,N_2975);
or UO_358 (O_358,N_2985,N_2956);
xnor UO_359 (O_359,N_2991,N_2955);
nand UO_360 (O_360,N_2968,N_2982);
and UO_361 (O_361,N_2952,N_2989);
nand UO_362 (O_362,N_2973,N_2998);
nor UO_363 (O_363,N_2951,N_2972);
nor UO_364 (O_364,N_2963,N_2957);
and UO_365 (O_365,N_2959,N_2993);
nor UO_366 (O_366,N_2958,N_2955);
nand UO_367 (O_367,N_2975,N_2952);
nor UO_368 (O_368,N_2974,N_2966);
or UO_369 (O_369,N_2954,N_2985);
xor UO_370 (O_370,N_2955,N_2994);
and UO_371 (O_371,N_2982,N_2980);
nor UO_372 (O_372,N_2976,N_2964);
xnor UO_373 (O_373,N_2979,N_2978);
and UO_374 (O_374,N_2982,N_2964);
and UO_375 (O_375,N_2997,N_2982);
or UO_376 (O_376,N_2996,N_2953);
or UO_377 (O_377,N_2958,N_2997);
or UO_378 (O_378,N_2979,N_2975);
and UO_379 (O_379,N_2978,N_2954);
nand UO_380 (O_380,N_2976,N_2956);
nand UO_381 (O_381,N_2963,N_2973);
xnor UO_382 (O_382,N_2974,N_2998);
nand UO_383 (O_383,N_2961,N_2982);
nand UO_384 (O_384,N_2983,N_2997);
and UO_385 (O_385,N_2950,N_2952);
xor UO_386 (O_386,N_2978,N_2956);
or UO_387 (O_387,N_2981,N_2993);
nand UO_388 (O_388,N_2966,N_2978);
nand UO_389 (O_389,N_2991,N_2983);
and UO_390 (O_390,N_2998,N_2988);
nor UO_391 (O_391,N_2960,N_2976);
nand UO_392 (O_392,N_2956,N_2991);
xor UO_393 (O_393,N_2980,N_2958);
and UO_394 (O_394,N_2960,N_2993);
nand UO_395 (O_395,N_2995,N_2957);
and UO_396 (O_396,N_2999,N_2974);
nand UO_397 (O_397,N_2979,N_2990);
nor UO_398 (O_398,N_2951,N_2995);
and UO_399 (O_399,N_2981,N_2991);
and UO_400 (O_400,N_2963,N_2985);
nor UO_401 (O_401,N_2950,N_2968);
nor UO_402 (O_402,N_2977,N_2950);
nor UO_403 (O_403,N_2958,N_2975);
nor UO_404 (O_404,N_2990,N_2995);
or UO_405 (O_405,N_2969,N_2974);
nor UO_406 (O_406,N_2992,N_2979);
xor UO_407 (O_407,N_2958,N_2981);
nor UO_408 (O_408,N_2953,N_2964);
xnor UO_409 (O_409,N_2986,N_2955);
nor UO_410 (O_410,N_2963,N_2992);
or UO_411 (O_411,N_2978,N_2981);
or UO_412 (O_412,N_2968,N_2992);
xor UO_413 (O_413,N_2967,N_2988);
or UO_414 (O_414,N_2958,N_2986);
nand UO_415 (O_415,N_2984,N_2975);
xnor UO_416 (O_416,N_2954,N_2952);
nand UO_417 (O_417,N_2999,N_2961);
xnor UO_418 (O_418,N_2970,N_2959);
nor UO_419 (O_419,N_2990,N_2983);
or UO_420 (O_420,N_2951,N_2999);
and UO_421 (O_421,N_2951,N_2978);
and UO_422 (O_422,N_2966,N_2951);
and UO_423 (O_423,N_2996,N_2998);
nand UO_424 (O_424,N_2964,N_2986);
nand UO_425 (O_425,N_2998,N_2989);
nor UO_426 (O_426,N_2967,N_2960);
nand UO_427 (O_427,N_2999,N_2978);
nand UO_428 (O_428,N_2969,N_2986);
nand UO_429 (O_429,N_2968,N_2963);
and UO_430 (O_430,N_2974,N_2962);
or UO_431 (O_431,N_2971,N_2980);
and UO_432 (O_432,N_2958,N_2967);
nor UO_433 (O_433,N_2994,N_2983);
nor UO_434 (O_434,N_2960,N_2997);
and UO_435 (O_435,N_2979,N_2954);
and UO_436 (O_436,N_2984,N_2983);
and UO_437 (O_437,N_2969,N_2952);
nand UO_438 (O_438,N_2958,N_2983);
and UO_439 (O_439,N_2974,N_2994);
xnor UO_440 (O_440,N_2958,N_2988);
or UO_441 (O_441,N_2977,N_2997);
and UO_442 (O_442,N_2999,N_2952);
and UO_443 (O_443,N_2951,N_2988);
and UO_444 (O_444,N_2962,N_2966);
or UO_445 (O_445,N_2989,N_2973);
xnor UO_446 (O_446,N_2983,N_2981);
and UO_447 (O_447,N_2997,N_2962);
and UO_448 (O_448,N_2971,N_2992);
or UO_449 (O_449,N_2969,N_2995);
nor UO_450 (O_450,N_2962,N_2991);
and UO_451 (O_451,N_2965,N_2968);
nand UO_452 (O_452,N_2964,N_2994);
or UO_453 (O_453,N_2987,N_2992);
xnor UO_454 (O_454,N_2970,N_2998);
nor UO_455 (O_455,N_2988,N_2977);
and UO_456 (O_456,N_2996,N_2972);
nor UO_457 (O_457,N_2989,N_2959);
or UO_458 (O_458,N_2959,N_2982);
nand UO_459 (O_459,N_2974,N_2958);
xor UO_460 (O_460,N_2969,N_2965);
xor UO_461 (O_461,N_2998,N_2968);
and UO_462 (O_462,N_2956,N_2964);
and UO_463 (O_463,N_2999,N_2972);
and UO_464 (O_464,N_2990,N_2993);
nor UO_465 (O_465,N_2955,N_2988);
xnor UO_466 (O_466,N_2970,N_2952);
and UO_467 (O_467,N_2964,N_2997);
nand UO_468 (O_468,N_2977,N_2957);
xnor UO_469 (O_469,N_2988,N_2965);
nor UO_470 (O_470,N_2988,N_2953);
nand UO_471 (O_471,N_2977,N_2991);
nand UO_472 (O_472,N_2959,N_2984);
and UO_473 (O_473,N_2989,N_2950);
and UO_474 (O_474,N_2970,N_2987);
nand UO_475 (O_475,N_2956,N_2972);
xnor UO_476 (O_476,N_2966,N_2995);
xor UO_477 (O_477,N_2979,N_2969);
xor UO_478 (O_478,N_2962,N_2968);
nor UO_479 (O_479,N_2985,N_2997);
nand UO_480 (O_480,N_2968,N_2971);
and UO_481 (O_481,N_2968,N_2978);
xnor UO_482 (O_482,N_2968,N_2974);
or UO_483 (O_483,N_2956,N_2973);
or UO_484 (O_484,N_2973,N_2967);
nor UO_485 (O_485,N_2993,N_2997);
or UO_486 (O_486,N_2967,N_2994);
and UO_487 (O_487,N_2976,N_2983);
and UO_488 (O_488,N_2988,N_2994);
or UO_489 (O_489,N_2953,N_2963);
nand UO_490 (O_490,N_2999,N_2950);
xor UO_491 (O_491,N_2969,N_2962);
nand UO_492 (O_492,N_2987,N_2953);
nor UO_493 (O_493,N_2956,N_2995);
xor UO_494 (O_494,N_2982,N_2985);
nand UO_495 (O_495,N_2990,N_2962);
and UO_496 (O_496,N_2980,N_2985);
nand UO_497 (O_497,N_2980,N_2954);
nor UO_498 (O_498,N_2957,N_2961);
and UO_499 (O_499,N_2989,N_2999);
endmodule