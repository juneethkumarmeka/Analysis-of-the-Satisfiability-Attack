module basic_500_3000_500_5_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_211,In_332);
nand U1 (N_1,In_304,In_461);
or U2 (N_2,In_421,In_83);
xor U3 (N_3,In_121,In_56);
xnor U4 (N_4,In_440,In_334);
and U5 (N_5,In_169,In_23);
nor U6 (N_6,In_66,In_87);
xnor U7 (N_7,In_481,In_415);
xor U8 (N_8,In_132,In_371);
nor U9 (N_9,In_271,In_99);
and U10 (N_10,In_310,In_411);
xnor U11 (N_11,In_399,In_351);
xnor U12 (N_12,In_179,In_320);
xor U13 (N_13,In_424,In_153);
xor U14 (N_14,In_284,In_64);
and U15 (N_15,In_115,In_196);
xnor U16 (N_16,In_472,In_491);
xor U17 (N_17,In_279,In_14);
xnor U18 (N_18,In_376,In_344);
or U19 (N_19,In_474,In_58);
or U20 (N_20,In_378,In_268);
nand U21 (N_21,In_273,In_57);
nand U22 (N_22,In_217,In_362);
or U23 (N_23,In_435,In_164);
xnor U24 (N_24,In_293,In_408);
nor U25 (N_25,In_163,In_251);
nand U26 (N_26,In_100,In_6);
xor U27 (N_27,In_463,In_88);
or U28 (N_28,In_390,In_219);
or U29 (N_29,In_89,In_433);
nor U30 (N_30,In_84,In_50);
xnor U31 (N_31,In_29,In_246);
or U32 (N_32,In_48,In_456);
or U33 (N_33,In_45,In_395);
nor U34 (N_34,In_479,In_85);
xnor U35 (N_35,In_483,In_361);
and U36 (N_36,In_436,In_218);
nand U37 (N_37,In_488,In_135);
nor U38 (N_38,In_499,In_37);
nand U39 (N_39,In_226,In_450);
or U40 (N_40,In_46,In_368);
nor U41 (N_41,In_462,In_72);
nor U42 (N_42,In_190,In_397);
nor U43 (N_43,In_314,In_144);
nor U44 (N_44,In_276,In_119);
nor U45 (N_45,In_400,In_496);
and U46 (N_46,In_471,In_322);
nor U47 (N_47,In_283,In_125);
and U48 (N_48,In_467,In_487);
nor U49 (N_49,In_10,In_188);
nand U50 (N_50,In_384,In_228);
nor U51 (N_51,In_388,In_297);
and U52 (N_52,In_470,In_262);
nor U53 (N_53,In_43,In_128);
and U54 (N_54,In_137,In_401);
nor U55 (N_55,In_382,In_221);
or U56 (N_56,In_156,In_51);
or U57 (N_57,In_103,In_489);
and U58 (N_58,In_212,In_292);
and U59 (N_59,In_392,In_347);
or U60 (N_60,In_73,In_389);
or U61 (N_61,In_383,In_363);
xor U62 (N_62,In_59,In_231);
nor U63 (N_63,In_187,In_272);
nand U64 (N_64,In_107,In_138);
nand U65 (N_65,In_140,In_108);
nand U66 (N_66,In_189,In_86);
or U67 (N_67,In_186,In_431);
nand U68 (N_68,In_303,In_475);
nor U69 (N_69,In_166,In_194);
xor U70 (N_70,In_39,In_12);
xnor U71 (N_71,In_373,In_213);
xor U72 (N_72,In_13,In_236);
nand U73 (N_73,In_274,In_198);
nand U74 (N_74,In_305,In_277);
xnor U75 (N_75,In_33,In_35);
and U76 (N_76,In_148,In_18);
nand U77 (N_77,In_91,In_340);
and U78 (N_78,In_124,In_230);
xnor U79 (N_79,In_430,In_101);
and U80 (N_80,In_4,In_63);
xnor U81 (N_81,In_206,In_321);
nor U82 (N_82,In_146,In_345);
or U83 (N_83,In_437,In_337);
nand U84 (N_84,In_282,In_466);
xor U85 (N_85,In_242,In_453);
xor U86 (N_86,In_403,In_323);
or U87 (N_87,In_75,In_417);
nor U88 (N_88,In_495,In_289);
and U89 (N_89,In_42,In_405);
nor U90 (N_90,In_404,In_315);
or U91 (N_91,In_357,In_497);
xnor U92 (N_92,In_105,In_182);
xnor U93 (N_93,In_478,In_386);
nand U94 (N_94,In_61,In_239);
nor U95 (N_95,In_53,In_222);
xor U96 (N_96,In_252,In_36);
nand U97 (N_97,In_191,In_302);
or U98 (N_98,In_342,In_449);
nand U99 (N_99,In_192,In_260);
and U100 (N_100,In_16,In_377);
nand U101 (N_101,In_258,In_327);
and U102 (N_102,In_459,In_142);
and U103 (N_103,In_193,In_269);
nor U104 (N_104,In_253,In_387);
nor U105 (N_105,In_241,In_468);
and U106 (N_106,In_157,In_328);
and U107 (N_107,In_299,In_126);
nand U108 (N_108,In_110,In_17);
nor U109 (N_109,In_71,In_141);
and U110 (N_110,In_224,In_233);
or U111 (N_111,In_358,In_133);
xnor U112 (N_112,In_195,In_95);
and U113 (N_113,In_1,In_365);
nor U114 (N_114,In_280,In_367);
nand U115 (N_115,In_353,In_385);
nor U116 (N_116,In_354,In_234);
xnor U117 (N_117,In_446,In_352);
nor U118 (N_118,In_38,In_264);
and U119 (N_119,In_287,In_341);
or U120 (N_120,In_174,In_47);
nor U121 (N_121,In_24,In_476);
or U122 (N_122,In_123,In_288);
or U123 (N_123,In_22,In_129);
nand U124 (N_124,In_8,In_469);
or U125 (N_125,In_9,In_177);
nor U126 (N_126,In_396,In_199);
nor U127 (N_127,In_21,In_216);
or U128 (N_128,In_366,In_202);
xor U129 (N_129,In_257,In_55);
nand U130 (N_130,In_170,In_145);
nor U131 (N_131,In_7,In_432);
and U132 (N_132,In_444,In_171);
xnor U133 (N_133,In_423,In_318);
and U134 (N_134,In_448,In_154);
nand U135 (N_135,In_291,In_498);
and U136 (N_136,In_243,In_457);
and U137 (N_137,In_374,In_316);
nor U138 (N_138,In_152,In_197);
and U139 (N_139,In_434,In_317);
or U140 (N_140,In_313,In_494);
nand U141 (N_141,In_44,In_398);
or U142 (N_142,In_102,In_225);
xor U143 (N_143,In_215,In_116);
xnor U144 (N_144,In_369,In_406);
nand U145 (N_145,In_158,In_290);
nor U146 (N_146,In_52,In_90);
nor U147 (N_147,In_147,In_98);
and U148 (N_148,In_130,In_200);
or U149 (N_149,In_161,In_301);
xnor U150 (N_150,In_324,In_210);
nand U151 (N_151,In_261,In_412);
nand U152 (N_152,In_355,In_203);
or U153 (N_153,In_267,In_300);
nor U154 (N_154,In_247,In_379);
nand U155 (N_155,In_455,In_5);
nor U156 (N_156,In_410,In_482);
nor U157 (N_157,In_178,In_70);
nor U158 (N_158,In_402,In_428);
xor U159 (N_159,In_11,In_65);
xor U160 (N_160,In_254,In_442);
or U161 (N_161,In_28,In_360);
nor U162 (N_162,In_275,In_480);
xnor U163 (N_163,In_372,In_307);
nor U164 (N_164,In_113,In_40);
and U165 (N_165,In_165,In_460);
or U166 (N_166,In_441,In_114);
nand U167 (N_167,In_364,In_319);
or U168 (N_168,In_419,In_41);
or U169 (N_169,In_19,In_20);
and U170 (N_170,In_270,In_370);
and U171 (N_171,In_67,In_325);
or U172 (N_172,In_2,In_60);
or U173 (N_173,In_69,In_168);
xnor U174 (N_174,In_485,In_172);
xor U175 (N_175,In_92,In_32);
nor U176 (N_176,In_34,In_127);
and U177 (N_177,In_308,In_31);
or U178 (N_178,In_248,In_335);
xor U179 (N_179,In_68,In_160);
or U180 (N_180,In_349,In_429);
nor U181 (N_181,In_244,In_492);
or U182 (N_182,In_209,In_74);
or U183 (N_183,In_205,In_420);
and U184 (N_184,In_416,In_159);
or U185 (N_185,In_484,In_30);
and U186 (N_186,In_201,In_93);
nand U187 (N_187,In_391,In_312);
nor U188 (N_188,In_438,In_78);
nor U189 (N_189,In_311,In_413);
nand U190 (N_190,In_104,In_106);
or U191 (N_191,In_134,In_407);
xor U192 (N_192,In_204,In_296);
nand U193 (N_193,In_256,In_486);
xor U194 (N_194,In_167,In_62);
nand U195 (N_195,In_162,In_359);
or U196 (N_196,In_139,In_298);
xnor U197 (N_197,In_350,In_81);
and U198 (N_198,In_250,In_281);
and U199 (N_199,In_454,In_265);
nor U200 (N_200,In_426,In_339);
nor U201 (N_201,In_381,In_111);
nand U202 (N_202,In_375,In_15);
and U203 (N_203,In_229,In_477);
or U204 (N_204,In_208,In_285);
xnor U205 (N_205,In_25,In_94);
nand U206 (N_206,In_295,In_173);
nor U207 (N_207,In_27,In_185);
xnor U208 (N_208,In_235,In_136);
and U209 (N_209,In_286,In_180);
and U210 (N_210,In_309,In_249);
and U211 (N_211,In_330,In_394);
or U212 (N_212,In_445,In_175);
xnor U213 (N_213,In_96,In_490);
and U214 (N_214,In_0,In_447);
or U215 (N_215,In_150,In_263);
or U216 (N_216,In_26,In_76);
xor U217 (N_217,In_343,In_338);
and U218 (N_218,In_356,In_266);
nor U219 (N_219,In_331,In_183);
and U220 (N_220,In_443,In_184);
xor U221 (N_221,In_155,In_149);
or U222 (N_222,In_465,In_336);
nor U223 (N_223,In_418,In_227);
nand U224 (N_224,In_458,In_3);
or U225 (N_225,In_131,In_427);
nand U226 (N_226,In_223,In_151);
nor U227 (N_227,In_259,In_77);
nor U228 (N_228,In_473,In_439);
and U229 (N_229,In_380,In_329);
xor U230 (N_230,In_425,In_245);
nand U231 (N_231,In_238,In_122);
or U232 (N_232,In_326,In_214);
nor U233 (N_233,In_232,In_207);
and U234 (N_234,In_54,In_333);
and U235 (N_235,In_393,In_97);
nor U236 (N_236,In_181,In_176);
xor U237 (N_237,In_109,In_409);
or U238 (N_238,In_414,In_117);
and U239 (N_239,In_422,In_143);
xor U240 (N_240,In_464,In_237);
and U241 (N_241,In_112,In_120);
or U242 (N_242,In_118,In_255);
or U243 (N_243,In_452,In_82);
xor U244 (N_244,In_240,In_220);
or U245 (N_245,In_306,In_49);
or U246 (N_246,In_294,In_278);
or U247 (N_247,In_451,In_79);
and U248 (N_248,In_346,In_80);
nand U249 (N_249,In_493,In_348);
nor U250 (N_250,In_97,In_291);
and U251 (N_251,In_195,In_139);
nand U252 (N_252,In_351,In_343);
and U253 (N_253,In_384,In_495);
nor U254 (N_254,In_202,In_340);
xnor U255 (N_255,In_423,In_154);
nor U256 (N_256,In_415,In_348);
and U257 (N_257,In_302,In_408);
or U258 (N_258,In_170,In_13);
xnor U259 (N_259,In_199,In_119);
nand U260 (N_260,In_174,In_62);
or U261 (N_261,In_104,In_199);
and U262 (N_262,In_441,In_41);
or U263 (N_263,In_296,In_340);
nor U264 (N_264,In_297,In_220);
nor U265 (N_265,In_468,In_116);
or U266 (N_266,In_132,In_201);
nand U267 (N_267,In_67,In_283);
xnor U268 (N_268,In_342,In_293);
or U269 (N_269,In_153,In_365);
and U270 (N_270,In_21,In_6);
or U271 (N_271,In_191,In_100);
or U272 (N_272,In_127,In_395);
nor U273 (N_273,In_138,In_21);
nor U274 (N_274,In_453,In_97);
and U275 (N_275,In_50,In_56);
or U276 (N_276,In_45,In_85);
xor U277 (N_277,In_127,In_407);
nand U278 (N_278,In_439,In_31);
nor U279 (N_279,In_321,In_256);
and U280 (N_280,In_72,In_215);
nand U281 (N_281,In_313,In_202);
and U282 (N_282,In_156,In_35);
nand U283 (N_283,In_409,In_155);
xnor U284 (N_284,In_329,In_255);
xor U285 (N_285,In_315,In_373);
nand U286 (N_286,In_346,In_485);
nor U287 (N_287,In_289,In_138);
nand U288 (N_288,In_152,In_432);
nand U289 (N_289,In_171,In_353);
nor U290 (N_290,In_260,In_335);
and U291 (N_291,In_117,In_404);
xor U292 (N_292,In_382,In_234);
nor U293 (N_293,In_246,In_133);
nand U294 (N_294,In_147,In_388);
nand U295 (N_295,In_101,In_282);
nand U296 (N_296,In_338,In_275);
nor U297 (N_297,In_134,In_47);
and U298 (N_298,In_295,In_26);
xor U299 (N_299,In_479,In_293);
and U300 (N_300,In_96,In_64);
or U301 (N_301,In_473,In_188);
nand U302 (N_302,In_407,In_240);
nor U303 (N_303,In_50,In_93);
or U304 (N_304,In_4,In_394);
and U305 (N_305,In_451,In_323);
xor U306 (N_306,In_440,In_140);
xnor U307 (N_307,In_181,In_371);
nor U308 (N_308,In_185,In_190);
and U309 (N_309,In_53,In_403);
or U310 (N_310,In_88,In_485);
or U311 (N_311,In_123,In_297);
or U312 (N_312,In_95,In_39);
or U313 (N_313,In_326,In_347);
xnor U314 (N_314,In_337,In_230);
and U315 (N_315,In_60,In_490);
nand U316 (N_316,In_282,In_42);
nand U317 (N_317,In_208,In_255);
xnor U318 (N_318,In_192,In_76);
nand U319 (N_319,In_36,In_494);
nor U320 (N_320,In_75,In_486);
nor U321 (N_321,In_212,In_258);
or U322 (N_322,In_376,In_472);
nor U323 (N_323,In_181,In_305);
and U324 (N_324,In_496,In_161);
nor U325 (N_325,In_200,In_410);
or U326 (N_326,In_394,In_216);
nor U327 (N_327,In_207,In_389);
and U328 (N_328,In_51,In_254);
nor U329 (N_329,In_43,In_429);
and U330 (N_330,In_52,In_127);
or U331 (N_331,In_254,In_3);
nor U332 (N_332,In_132,In_143);
nand U333 (N_333,In_46,In_140);
or U334 (N_334,In_144,In_354);
nand U335 (N_335,In_353,In_496);
or U336 (N_336,In_8,In_136);
or U337 (N_337,In_133,In_73);
nand U338 (N_338,In_133,In_482);
and U339 (N_339,In_280,In_331);
or U340 (N_340,In_458,In_386);
nand U341 (N_341,In_460,In_140);
and U342 (N_342,In_117,In_17);
and U343 (N_343,In_146,In_429);
or U344 (N_344,In_201,In_494);
or U345 (N_345,In_233,In_304);
and U346 (N_346,In_118,In_422);
xnor U347 (N_347,In_421,In_334);
and U348 (N_348,In_183,In_58);
nor U349 (N_349,In_367,In_366);
or U350 (N_350,In_247,In_45);
nor U351 (N_351,In_297,In_197);
and U352 (N_352,In_307,In_417);
and U353 (N_353,In_412,In_21);
or U354 (N_354,In_159,In_5);
nor U355 (N_355,In_91,In_274);
nand U356 (N_356,In_241,In_47);
and U357 (N_357,In_66,In_424);
nor U358 (N_358,In_51,In_326);
and U359 (N_359,In_96,In_399);
and U360 (N_360,In_409,In_371);
nor U361 (N_361,In_484,In_320);
and U362 (N_362,In_38,In_384);
xnor U363 (N_363,In_16,In_191);
xnor U364 (N_364,In_85,In_101);
nor U365 (N_365,In_198,In_298);
and U366 (N_366,In_171,In_359);
or U367 (N_367,In_126,In_377);
or U368 (N_368,In_11,In_82);
and U369 (N_369,In_184,In_300);
nor U370 (N_370,In_234,In_433);
and U371 (N_371,In_462,In_146);
xnor U372 (N_372,In_447,In_246);
and U373 (N_373,In_379,In_332);
nand U374 (N_374,In_111,In_379);
nand U375 (N_375,In_121,In_438);
and U376 (N_376,In_129,In_81);
and U377 (N_377,In_57,In_112);
nand U378 (N_378,In_463,In_372);
or U379 (N_379,In_64,In_315);
xor U380 (N_380,In_137,In_98);
nor U381 (N_381,In_207,In_351);
nand U382 (N_382,In_86,In_147);
and U383 (N_383,In_272,In_466);
nor U384 (N_384,In_314,In_444);
or U385 (N_385,In_418,In_212);
and U386 (N_386,In_319,In_208);
nand U387 (N_387,In_221,In_240);
nor U388 (N_388,In_189,In_470);
nor U389 (N_389,In_314,In_178);
nand U390 (N_390,In_140,In_117);
and U391 (N_391,In_474,In_361);
and U392 (N_392,In_133,In_203);
or U393 (N_393,In_327,In_230);
nor U394 (N_394,In_248,In_218);
or U395 (N_395,In_364,In_97);
and U396 (N_396,In_446,In_20);
and U397 (N_397,In_237,In_153);
nand U398 (N_398,In_89,In_412);
or U399 (N_399,In_40,In_354);
or U400 (N_400,In_279,In_65);
nand U401 (N_401,In_489,In_17);
xor U402 (N_402,In_155,In_98);
nand U403 (N_403,In_296,In_289);
xor U404 (N_404,In_436,In_206);
nand U405 (N_405,In_360,In_151);
and U406 (N_406,In_402,In_153);
nor U407 (N_407,In_3,In_181);
nor U408 (N_408,In_389,In_70);
nand U409 (N_409,In_192,In_212);
and U410 (N_410,In_475,In_265);
xor U411 (N_411,In_35,In_141);
xor U412 (N_412,In_62,In_459);
nand U413 (N_413,In_451,In_420);
xor U414 (N_414,In_491,In_126);
nand U415 (N_415,In_393,In_382);
xor U416 (N_416,In_362,In_324);
xnor U417 (N_417,In_226,In_426);
nor U418 (N_418,In_91,In_228);
and U419 (N_419,In_138,In_368);
or U420 (N_420,In_77,In_305);
and U421 (N_421,In_468,In_205);
nor U422 (N_422,In_79,In_243);
and U423 (N_423,In_472,In_139);
nand U424 (N_424,In_255,In_376);
or U425 (N_425,In_475,In_367);
and U426 (N_426,In_263,In_380);
and U427 (N_427,In_77,In_368);
nand U428 (N_428,In_420,In_148);
nor U429 (N_429,In_261,In_427);
nor U430 (N_430,In_407,In_75);
or U431 (N_431,In_141,In_7);
xnor U432 (N_432,In_479,In_52);
xor U433 (N_433,In_121,In_339);
and U434 (N_434,In_150,In_152);
xnor U435 (N_435,In_396,In_84);
nor U436 (N_436,In_33,In_415);
and U437 (N_437,In_372,In_251);
and U438 (N_438,In_6,In_451);
or U439 (N_439,In_68,In_244);
and U440 (N_440,In_214,In_419);
xor U441 (N_441,In_450,In_23);
or U442 (N_442,In_68,In_263);
or U443 (N_443,In_14,In_64);
or U444 (N_444,In_278,In_7);
nor U445 (N_445,In_171,In_373);
nand U446 (N_446,In_408,In_22);
or U447 (N_447,In_158,In_107);
nand U448 (N_448,In_34,In_89);
xnor U449 (N_449,In_264,In_397);
nor U450 (N_450,In_62,In_395);
xor U451 (N_451,In_26,In_384);
nor U452 (N_452,In_87,In_481);
xnor U453 (N_453,In_255,In_439);
and U454 (N_454,In_260,In_328);
and U455 (N_455,In_129,In_349);
and U456 (N_456,In_240,In_171);
xor U457 (N_457,In_340,In_76);
xor U458 (N_458,In_333,In_415);
and U459 (N_459,In_200,In_445);
and U460 (N_460,In_241,In_200);
or U461 (N_461,In_271,In_176);
nor U462 (N_462,In_315,In_137);
xor U463 (N_463,In_139,In_396);
xnor U464 (N_464,In_318,In_203);
nand U465 (N_465,In_41,In_481);
nor U466 (N_466,In_102,In_395);
nand U467 (N_467,In_132,In_364);
xor U468 (N_468,In_61,In_325);
and U469 (N_469,In_389,In_278);
nand U470 (N_470,In_322,In_474);
xor U471 (N_471,In_478,In_167);
nand U472 (N_472,In_70,In_9);
xor U473 (N_473,In_23,In_166);
or U474 (N_474,In_429,In_361);
nand U475 (N_475,In_307,In_136);
or U476 (N_476,In_321,In_44);
xor U477 (N_477,In_92,In_315);
nor U478 (N_478,In_457,In_358);
or U479 (N_479,In_231,In_324);
xnor U480 (N_480,In_23,In_499);
nand U481 (N_481,In_60,In_277);
nand U482 (N_482,In_300,In_149);
or U483 (N_483,In_383,In_78);
nor U484 (N_484,In_145,In_220);
nor U485 (N_485,In_360,In_375);
nand U486 (N_486,In_360,In_381);
xnor U487 (N_487,In_332,In_185);
and U488 (N_488,In_142,In_480);
xor U489 (N_489,In_263,In_113);
xor U490 (N_490,In_199,In_160);
or U491 (N_491,In_80,In_392);
or U492 (N_492,In_109,In_305);
nand U493 (N_493,In_223,In_60);
nand U494 (N_494,In_431,In_304);
and U495 (N_495,In_199,In_211);
nor U496 (N_496,In_272,In_425);
or U497 (N_497,In_414,In_375);
nor U498 (N_498,In_393,In_319);
nand U499 (N_499,In_2,In_1);
nand U500 (N_500,In_204,In_132);
and U501 (N_501,In_105,In_183);
nor U502 (N_502,In_406,In_416);
xnor U503 (N_503,In_435,In_98);
nand U504 (N_504,In_398,In_274);
nand U505 (N_505,In_428,In_448);
or U506 (N_506,In_368,In_444);
nor U507 (N_507,In_267,In_399);
and U508 (N_508,In_386,In_14);
xnor U509 (N_509,In_66,In_476);
nor U510 (N_510,In_489,In_16);
and U511 (N_511,In_132,In_30);
nor U512 (N_512,In_371,In_3);
or U513 (N_513,In_12,In_492);
xor U514 (N_514,In_70,In_196);
xnor U515 (N_515,In_312,In_20);
nor U516 (N_516,In_374,In_111);
nand U517 (N_517,In_50,In_346);
nand U518 (N_518,In_430,In_248);
nor U519 (N_519,In_26,In_271);
and U520 (N_520,In_149,In_279);
xnor U521 (N_521,In_328,In_249);
or U522 (N_522,In_364,In_465);
nor U523 (N_523,In_493,In_484);
nand U524 (N_524,In_163,In_468);
and U525 (N_525,In_484,In_326);
or U526 (N_526,In_104,In_135);
or U527 (N_527,In_152,In_224);
nor U528 (N_528,In_207,In_212);
and U529 (N_529,In_47,In_401);
and U530 (N_530,In_69,In_404);
and U531 (N_531,In_241,In_378);
xor U532 (N_532,In_200,In_180);
or U533 (N_533,In_124,In_80);
xnor U534 (N_534,In_22,In_445);
or U535 (N_535,In_107,In_314);
nand U536 (N_536,In_462,In_52);
and U537 (N_537,In_465,In_41);
xnor U538 (N_538,In_449,In_64);
nor U539 (N_539,In_454,In_330);
nand U540 (N_540,In_183,In_483);
or U541 (N_541,In_252,In_96);
or U542 (N_542,In_261,In_464);
and U543 (N_543,In_469,In_65);
and U544 (N_544,In_269,In_112);
nor U545 (N_545,In_493,In_324);
xor U546 (N_546,In_10,In_425);
nor U547 (N_547,In_444,In_120);
nand U548 (N_548,In_332,In_436);
nor U549 (N_549,In_135,In_344);
nor U550 (N_550,In_267,In_394);
nor U551 (N_551,In_92,In_103);
xnor U552 (N_552,In_247,In_354);
nand U553 (N_553,In_73,In_481);
nand U554 (N_554,In_290,In_222);
xnor U555 (N_555,In_121,In_125);
xor U556 (N_556,In_58,In_80);
nor U557 (N_557,In_434,In_0);
and U558 (N_558,In_283,In_363);
or U559 (N_559,In_450,In_150);
nand U560 (N_560,In_419,In_2);
and U561 (N_561,In_431,In_127);
xnor U562 (N_562,In_82,In_424);
xnor U563 (N_563,In_175,In_427);
xnor U564 (N_564,In_177,In_211);
xor U565 (N_565,In_95,In_233);
or U566 (N_566,In_136,In_481);
xor U567 (N_567,In_387,In_386);
or U568 (N_568,In_260,In_184);
and U569 (N_569,In_197,In_6);
nor U570 (N_570,In_358,In_440);
and U571 (N_571,In_131,In_64);
or U572 (N_572,In_107,In_168);
nand U573 (N_573,In_452,In_201);
nand U574 (N_574,In_357,In_207);
or U575 (N_575,In_176,In_436);
nand U576 (N_576,In_199,In_152);
nand U577 (N_577,In_273,In_433);
or U578 (N_578,In_237,In_61);
and U579 (N_579,In_147,In_287);
nand U580 (N_580,In_38,In_98);
xnor U581 (N_581,In_119,In_319);
nor U582 (N_582,In_52,In_222);
or U583 (N_583,In_96,In_90);
nand U584 (N_584,In_0,In_250);
and U585 (N_585,In_5,In_428);
or U586 (N_586,In_383,In_189);
nand U587 (N_587,In_100,In_220);
and U588 (N_588,In_176,In_240);
nand U589 (N_589,In_361,In_113);
or U590 (N_590,In_300,In_46);
and U591 (N_591,In_329,In_113);
xor U592 (N_592,In_488,In_253);
and U593 (N_593,In_73,In_23);
nand U594 (N_594,In_8,In_325);
nand U595 (N_595,In_172,In_175);
or U596 (N_596,In_105,In_111);
nand U597 (N_597,In_174,In_165);
and U598 (N_598,In_201,In_387);
or U599 (N_599,In_269,In_172);
and U600 (N_600,N_133,N_278);
or U601 (N_601,N_544,N_367);
and U602 (N_602,N_120,N_210);
nand U603 (N_603,N_425,N_522);
or U604 (N_604,N_272,N_294);
and U605 (N_605,N_274,N_32);
nand U606 (N_606,N_22,N_213);
xnor U607 (N_607,N_434,N_387);
and U608 (N_608,N_147,N_591);
nor U609 (N_609,N_471,N_26);
xor U610 (N_610,N_571,N_288);
and U611 (N_611,N_577,N_500);
nand U612 (N_612,N_372,N_15);
nand U613 (N_613,N_469,N_146);
xnor U614 (N_614,N_240,N_221);
xor U615 (N_615,N_583,N_145);
and U616 (N_616,N_142,N_590);
or U617 (N_617,N_325,N_289);
xnor U618 (N_618,N_47,N_118);
or U619 (N_619,N_124,N_198);
xnor U620 (N_620,N_230,N_308);
nand U621 (N_621,N_380,N_297);
nor U622 (N_622,N_549,N_323);
and U623 (N_623,N_4,N_324);
nand U624 (N_624,N_414,N_113);
xor U625 (N_625,N_537,N_538);
or U626 (N_626,N_354,N_438);
and U627 (N_627,N_182,N_532);
and U628 (N_628,N_542,N_408);
nor U629 (N_629,N_62,N_72);
xor U630 (N_630,N_29,N_448);
nor U631 (N_631,N_334,N_228);
xor U632 (N_632,N_348,N_150);
and U633 (N_633,N_135,N_598);
and U634 (N_634,N_444,N_239);
nand U635 (N_635,N_467,N_59);
or U636 (N_636,N_580,N_291);
nor U637 (N_637,N_151,N_319);
nor U638 (N_638,N_514,N_546);
nor U639 (N_639,N_498,N_117);
nor U640 (N_640,N_392,N_31);
nor U641 (N_641,N_592,N_106);
and U642 (N_642,N_49,N_183);
and U643 (N_643,N_488,N_474);
nor U644 (N_644,N_231,N_77);
nand U645 (N_645,N_365,N_171);
and U646 (N_646,N_364,N_395);
nor U647 (N_647,N_588,N_163);
xor U648 (N_648,N_453,N_84);
and U649 (N_649,N_557,N_69);
nand U650 (N_650,N_45,N_115);
or U651 (N_651,N_369,N_521);
and U652 (N_652,N_505,N_200);
xnor U653 (N_653,N_341,N_596);
or U654 (N_654,N_340,N_470);
or U655 (N_655,N_197,N_275);
nor U656 (N_656,N_559,N_545);
and U657 (N_657,N_122,N_597);
or U658 (N_658,N_480,N_349);
xnor U659 (N_659,N_258,N_377);
or U660 (N_660,N_180,N_271);
or U661 (N_661,N_292,N_357);
and U662 (N_662,N_322,N_335);
nand U663 (N_663,N_581,N_24);
nor U664 (N_664,N_23,N_130);
and U665 (N_665,N_279,N_98);
xor U666 (N_666,N_35,N_86);
nor U667 (N_667,N_534,N_304);
xnor U668 (N_668,N_519,N_423);
or U669 (N_669,N_28,N_393);
xor U670 (N_670,N_137,N_497);
nand U671 (N_671,N_5,N_424);
or U672 (N_672,N_277,N_513);
nor U673 (N_673,N_208,N_572);
and U674 (N_674,N_83,N_55);
xor U675 (N_675,N_104,N_337);
and U676 (N_676,N_1,N_579);
nor U677 (N_677,N_458,N_389);
nor U678 (N_678,N_490,N_344);
and U679 (N_679,N_242,N_381);
and U680 (N_680,N_456,N_44);
xnor U681 (N_681,N_290,N_310);
or U682 (N_682,N_382,N_516);
and U683 (N_683,N_353,N_515);
and U684 (N_684,N_529,N_578);
and U685 (N_685,N_398,N_595);
nand U686 (N_686,N_539,N_114);
or U687 (N_687,N_184,N_276);
nor U688 (N_688,N_193,N_384);
nand U689 (N_689,N_439,N_233);
nor U690 (N_690,N_227,N_352);
xnor U691 (N_691,N_134,N_431);
xor U692 (N_692,N_533,N_76);
nand U693 (N_693,N_174,N_191);
nand U694 (N_694,N_298,N_587);
nand U695 (N_695,N_586,N_493);
nand U696 (N_696,N_252,N_415);
or U697 (N_697,N_40,N_573);
or U698 (N_698,N_442,N_375);
nor U699 (N_699,N_87,N_351);
and U700 (N_700,N_284,N_269);
xnor U701 (N_701,N_91,N_373);
xor U702 (N_702,N_136,N_58);
or U703 (N_703,N_41,N_419);
or U704 (N_704,N_259,N_565);
or U705 (N_705,N_479,N_251);
or U706 (N_706,N_440,N_237);
nor U707 (N_707,N_201,N_396);
nor U708 (N_708,N_313,N_478);
xnor U709 (N_709,N_404,N_202);
or U710 (N_710,N_388,N_207);
or U711 (N_711,N_312,N_574);
nor U712 (N_712,N_486,N_394);
or U713 (N_713,N_222,N_46);
nor U714 (N_714,N_543,N_132);
nor U715 (N_715,N_93,N_386);
or U716 (N_716,N_52,N_236);
and U717 (N_717,N_260,N_492);
nor U718 (N_718,N_75,N_64);
nor U719 (N_719,N_90,N_528);
and U720 (N_720,N_166,N_331);
nor U721 (N_721,N_74,N_105);
nor U722 (N_722,N_244,N_125);
or U723 (N_723,N_306,N_356);
xnor U724 (N_724,N_599,N_320);
xor U725 (N_725,N_422,N_461);
nor U726 (N_726,N_282,N_451);
xnor U727 (N_727,N_441,N_346);
nor U728 (N_728,N_165,N_266);
and U729 (N_729,N_462,N_343);
nor U730 (N_730,N_280,N_447);
xor U731 (N_731,N_333,N_303);
nand U732 (N_732,N_9,N_0);
xnor U733 (N_733,N_400,N_195);
and U734 (N_734,N_78,N_556);
or U735 (N_735,N_168,N_378);
nand U736 (N_736,N_33,N_273);
nand U737 (N_737,N_65,N_501);
nor U738 (N_738,N_216,N_170);
nand U739 (N_739,N_296,N_121);
or U740 (N_740,N_428,N_407);
or U741 (N_741,N_108,N_358);
nor U742 (N_742,N_494,N_39);
nor U743 (N_743,N_156,N_531);
or U744 (N_744,N_265,N_570);
or U745 (N_745,N_229,N_558);
nor U746 (N_746,N_164,N_432);
xnor U747 (N_747,N_92,N_16);
nor U748 (N_748,N_552,N_116);
and U749 (N_749,N_487,N_548);
nand U750 (N_750,N_249,N_88);
nor U751 (N_751,N_67,N_502);
or U752 (N_752,N_109,N_219);
or U753 (N_753,N_550,N_185);
or U754 (N_754,N_148,N_30);
nor U755 (N_755,N_504,N_568);
or U756 (N_756,N_60,N_594);
nand U757 (N_757,N_466,N_158);
xor U758 (N_758,N_68,N_263);
nand U759 (N_759,N_245,N_25);
xor U760 (N_760,N_175,N_336);
nor U761 (N_761,N_17,N_270);
and U762 (N_762,N_405,N_359);
nand U763 (N_763,N_100,N_347);
nand U764 (N_764,N_141,N_192);
nand U765 (N_765,N_172,N_547);
or U766 (N_766,N_443,N_264);
or U767 (N_767,N_436,N_140);
or U768 (N_768,N_311,N_473);
nand U769 (N_769,N_330,N_567);
xor U770 (N_770,N_411,N_173);
and U771 (N_771,N_287,N_126);
or U772 (N_772,N_293,N_307);
nor U773 (N_773,N_257,N_302);
and U774 (N_774,N_187,N_226);
xor U775 (N_775,N_194,N_243);
xnor U776 (N_776,N_34,N_540);
and U777 (N_777,N_262,N_256);
nor U778 (N_778,N_555,N_309);
nor U779 (N_779,N_177,N_535);
nor U780 (N_780,N_261,N_564);
or U781 (N_781,N_220,N_518);
xor U782 (N_782,N_464,N_383);
nor U783 (N_783,N_169,N_246);
and U784 (N_784,N_268,N_433);
nor U785 (N_785,N_223,N_460);
nand U786 (N_786,N_162,N_397);
and U787 (N_787,N_224,N_454);
nor U788 (N_788,N_426,N_152);
nor U789 (N_789,N_523,N_7);
and U790 (N_790,N_318,N_102);
and U791 (N_791,N_566,N_332);
and U792 (N_792,N_430,N_153);
or U793 (N_793,N_362,N_110);
nand U794 (N_794,N_520,N_338);
and U795 (N_795,N_412,N_285);
or U796 (N_796,N_339,N_101);
nor U797 (N_797,N_360,N_154);
xnor U798 (N_798,N_370,N_112);
nor U799 (N_799,N_89,N_329);
xnor U800 (N_800,N_85,N_495);
xor U801 (N_801,N_551,N_584);
nor U802 (N_802,N_496,N_80);
and U803 (N_803,N_81,N_476);
nor U804 (N_804,N_96,N_321);
xnor U805 (N_805,N_399,N_61);
and U806 (N_806,N_131,N_218);
nand U807 (N_807,N_286,N_11);
nor U808 (N_808,N_119,N_211);
xnor U809 (N_809,N_452,N_209);
nor U810 (N_810,N_12,N_199);
or U811 (N_811,N_526,N_235);
xnor U812 (N_812,N_160,N_512);
xor U813 (N_813,N_123,N_79);
or U814 (N_814,N_316,N_305);
xor U815 (N_815,N_481,N_129);
nand U816 (N_816,N_477,N_582);
nand U817 (N_817,N_484,N_234);
and U818 (N_818,N_485,N_576);
nor U819 (N_819,N_36,N_585);
xnor U820 (N_820,N_449,N_253);
and U821 (N_821,N_128,N_575);
or U822 (N_822,N_517,N_524);
xnor U823 (N_823,N_589,N_53);
nor U824 (N_824,N_181,N_390);
or U825 (N_825,N_37,N_376);
nor U826 (N_826,N_10,N_463);
and U827 (N_827,N_315,N_3);
xor U828 (N_828,N_435,N_155);
and U829 (N_829,N_299,N_73);
nor U830 (N_830,N_6,N_50);
nand U831 (N_831,N_176,N_314);
xor U832 (N_832,N_48,N_281);
and U833 (N_833,N_161,N_295);
nor U834 (N_834,N_379,N_465);
and U835 (N_835,N_525,N_374);
or U836 (N_836,N_507,N_506);
xnor U837 (N_837,N_94,N_541);
and U838 (N_838,N_569,N_418);
nand U839 (N_839,N_491,N_188);
and U840 (N_840,N_317,N_403);
nand U841 (N_841,N_127,N_250);
and U842 (N_842,N_149,N_429);
nor U843 (N_843,N_593,N_366);
xor U844 (N_844,N_247,N_189);
and U845 (N_845,N_416,N_472);
or U846 (N_846,N_437,N_527);
and U847 (N_847,N_361,N_483);
nand U848 (N_848,N_238,N_326);
xnor U849 (N_849,N_482,N_232);
or U850 (N_850,N_97,N_159);
xor U851 (N_851,N_21,N_459);
nor U852 (N_852,N_421,N_13);
xor U853 (N_853,N_203,N_450);
nand U854 (N_854,N_475,N_196);
nor U855 (N_855,N_371,N_509);
nor U856 (N_856,N_489,N_511);
and U857 (N_857,N_508,N_178);
nor U858 (N_858,N_71,N_560);
nand U859 (N_859,N_385,N_19);
or U860 (N_860,N_14,N_157);
nor U861 (N_861,N_345,N_536);
and U862 (N_862,N_457,N_215);
and U863 (N_863,N_327,N_401);
or U864 (N_864,N_57,N_255);
and U865 (N_865,N_205,N_563);
nor U866 (N_866,N_363,N_42);
nor U867 (N_867,N_139,N_410);
nor U868 (N_868,N_38,N_300);
nand U869 (N_869,N_43,N_204);
or U870 (N_870,N_186,N_107);
nor U871 (N_871,N_103,N_143);
or U872 (N_872,N_561,N_214);
and U873 (N_873,N_409,N_455);
nor U874 (N_874,N_562,N_413);
or U875 (N_875,N_445,N_54);
nor U876 (N_876,N_225,N_510);
xor U877 (N_877,N_503,N_70);
nand U878 (N_878,N_63,N_554);
nand U879 (N_879,N_190,N_241);
nor U880 (N_880,N_406,N_82);
or U881 (N_881,N_212,N_217);
and U882 (N_882,N_51,N_27);
xor U883 (N_883,N_66,N_342);
and U884 (N_884,N_468,N_446);
nand U885 (N_885,N_499,N_355);
xor U886 (N_886,N_138,N_8);
nor U887 (N_887,N_350,N_95);
nor U888 (N_888,N_283,N_20);
nand U889 (N_889,N_248,N_368);
nor U890 (N_890,N_328,N_56);
xnor U891 (N_891,N_301,N_391);
and U892 (N_892,N_530,N_167);
and U893 (N_893,N_417,N_254);
nand U894 (N_894,N_420,N_427);
nor U895 (N_895,N_111,N_206);
or U896 (N_896,N_144,N_99);
nand U897 (N_897,N_18,N_2);
or U898 (N_898,N_553,N_267);
and U899 (N_899,N_402,N_179);
nor U900 (N_900,N_263,N_597);
and U901 (N_901,N_579,N_172);
or U902 (N_902,N_361,N_282);
and U903 (N_903,N_474,N_404);
nand U904 (N_904,N_175,N_548);
nor U905 (N_905,N_291,N_152);
nor U906 (N_906,N_422,N_60);
nand U907 (N_907,N_184,N_56);
xnor U908 (N_908,N_421,N_269);
nor U909 (N_909,N_141,N_107);
nand U910 (N_910,N_14,N_175);
nor U911 (N_911,N_22,N_350);
nand U912 (N_912,N_137,N_152);
or U913 (N_913,N_174,N_377);
xor U914 (N_914,N_171,N_595);
or U915 (N_915,N_183,N_56);
xnor U916 (N_916,N_95,N_216);
xor U917 (N_917,N_446,N_399);
and U918 (N_918,N_339,N_428);
nor U919 (N_919,N_361,N_348);
xor U920 (N_920,N_432,N_125);
or U921 (N_921,N_303,N_144);
and U922 (N_922,N_357,N_39);
nor U923 (N_923,N_149,N_23);
and U924 (N_924,N_11,N_372);
and U925 (N_925,N_218,N_213);
and U926 (N_926,N_192,N_362);
nand U927 (N_927,N_8,N_208);
and U928 (N_928,N_588,N_415);
or U929 (N_929,N_238,N_258);
and U930 (N_930,N_63,N_164);
xnor U931 (N_931,N_349,N_149);
and U932 (N_932,N_189,N_484);
nor U933 (N_933,N_158,N_229);
xor U934 (N_934,N_491,N_514);
and U935 (N_935,N_79,N_466);
nand U936 (N_936,N_137,N_379);
xnor U937 (N_937,N_258,N_342);
and U938 (N_938,N_492,N_169);
and U939 (N_939,N_336,N_516);
nand U940 (N_940,N_121,N_485);
or U941 (N_941,N_445,N_423);
and U942 (N_942,N_532,N_112);
and U943 (N_943,N_569,N_526);
or U944 (N_944,N_533,N_237);
nand U945 (N_945,N_219,N_528);
or U946 (N_946,N_514,N_404);
nor U947 (N_947,N_514,N_480);
nor U948 (N_948,N_411,N_513);
xor U949 (N_949,N_402,N_141);
and U950 (N_950,N_404,N_333);
and U951 (N_951,N_212,N_264);
and U952 (N_952,N_553,N_95);
or U953 (N_953,N_367,N_511);
nor U954 (N_954,N_374,N_390);
and U955 (N_955,N_221,N_350);
nor U956 (N_956,N_41,N_431);
and U957 (N_957,N_369,N_444);
xor U958 (N_958,N_26,N_35);
nor U959 (N_959,N_446,N_386);
xnor U960 (N_960,N_163,N_426);
xor U961 (N_961,N_237,N_111);
xor U962 (N_962,N_251,N_495);
or U963 (N_963,N_59,N_487);
nor U964 (N_964,N_366,N_381);
xor U965 (N_965,N_141,N_506);
nand U966 (N_966,N_260,N_110);
or U967 (N_967,N_286,N_348);
and U968 (N_968,N_5,N_439);
nor U969 (N_969,N_519,N_175);
or U970 (N_970,N_431,N_62);
xnor U971 (N_971,N_531,N_217);
or U972 (N_972,N_482,N_362);
xnor U973 (N_973,N_117,N_528);
xor U974 (N_974,N_572,N_180);
and U975 (N_975,N_1,N_264);
and U976 (N_976,N_369,N_306);
and U977 (N_977,N_347,N_556);
nand U978 (N_978,N_504,N_213);
nand U979 (N_979,N_454,N_122);
or U980 (N_980,N_351,N_75);
nor U981 (N_981,N_568,N_86);
nor U982 (N_982,N_307,N_5);
and U983 (N_983,N_36,N_28);
and U984 (N_984,N_325,N_542);
xor U985 (N_985,N_429,N_247);
nand U986 (N_986,N_235,N_510);
xnor U987 (N_987,N_69,N_229);
and U988 (N_988,N_273,N_325);
nor U989 (N_989,N_53,N_56);
or U990 (N_990,N_587,N_145);
nand U991 (N_991,N_96,N_316);
nand U992 (N_992,N_165,N_448);
xnor U993 (N_993,N_122,N_5);
xor U994 (N_994,N_262,N_517);
or U995 (N_995,N_190,N_436);
xnor U996 (N_996,N_506,N_67);
or U997 (N_997,N_98,N_518);
or U998 (N_998,N_353,N_217);
and U999 (N_999,N_449,N_136);
nor U1000 (N_1000,N_75,N_569);
or U1001 (N_1001,N_577,N_234);
nand U1002 (N_1002,N_302,N_424);
xnor U1003 (N_1003,N_52,N_592);
nor U1004 (N_1004,N_404,N_578);
or U1005 (N_1005,N_418,N_212);
nand U1006 (N_1006,N_371,N_359);
or U1007 (N_1007,N_598,N_37);
or U1008 (N_1008,N_486,N_530);
nor U1009 (N_1009,N_48,N_390);
xnor U1010 (N_1010,N_234,N_68);
or U1011 (N_1011,N_376,N_497);
nor U1012 (N_1012,N_203,N_363);
and U1013 (N_1013,N_550,N_574);
or U1014 (N_1014,N_385,N_17);
nand U1015 (N_1015,N_84,N_466);
nor U1016 (N_1016,N_117,N_303);
xor U1017 (N_1017,N_576,N_589);
or U1018 (N_1018,N_314,N_34);
and U1019 (N_1019,N_161,N_581);
nor U1020 (N_1020,N_519,N_14);
nor U1021 (N_1021,N_570,N_480);
nor U1022 (N_1022,N_131,N_549);
nand U1023 (N_1023,N_152,N_458);
or U1024 (N_1024,N_197,N_254);
nand U1025 (N_1025,N_386,N_498);
nor U1026 (N_1026,N_162,N_245);
or U1027 (N_1027,N_243,N_66);
xnor U1028 (N_1028,N_449,N_184);
nand U1029 (N_1029,N_191,N_159);
nand U1030 (N_1030,N_159,N_485);
and U1031 (N_1031,N_339,N_594);
and U1032 (N_1032,N_439,N_467);
and U1033 (N_1033,N_242,N_561);
xnor U1034 (N_1034,N_376,N_557);
xor U1035 (N_1035,N_155,N_565);
xor U1036 (N_1036,N_433,N_498);
and U1037 (N_1037,N_103,N_145);
xor U1038 (N_1038,N_38,N_583);
nor U1039 (N_1039,N_566,N_61);
xor U1040 (N_1040,N_296,N_292);
or U1041 (N_1041,N_467,N_454);
and U1042 (N_1042,N_80,N_222);
or U1043 (N_1043,N_363,N_190);
and U1044 (N_1044,N_219,N_33);
xor U1045 (N_1045,N_423,N_407);
nor U1046 (N_1046,N_597,N_524);
and U1047 (N_1047,N_483,N_367);
xnor U1048 (N_1048,N_12,N_512);
and U1049 (N_1049,N_178,N_365);
nor U1050 (N_1050,N_261,N_190);
xor U1051 (N_1051,N_96,N_253);
nand U1052 (N_1052,N_283,N_455);
and U1053 (N_1053,N_592,N_269);
nor U1054 (N_1054,N_429,N_185);
and U1055 (N_1055,N_539,N_425);
or U1056 (N_1056,N_266,N_486);
or U1057 (N_1057,N_559,N_350);
xor U1058 (N_1058,N_413,N_116);
and U1059 (N_1059,N_337,N_17);
or U1060 (N_1060,N_144,N_308);
xor U1061 (N_1061,N_84,N_382);
nor U1062 (N_1062,N_564,N_223);
or U1063 (N_1063,N_227,N_407);
xnor U1064 (N_1064,N_372,N_117);
or U1065 (N_1065,N_443,N_98);
nand U1066 (N_1066,N_342,N_405);
and U1067 (N_1067,N_221,N_159);
nand U1068 (N_1068,N_236,N_298);
and U1069 (N_1069,N_131,N_242);
xor U1070 (N_1070,N_525,N_394);
nor U1071 (N_1071,N_298,N_165);
nand U1072 (N_1072,N_418,N_449);
nor U1073 (N_1073,N_569,N_553);
nand U1074 (N_1074,N_160,N_409);
or U1075 (N_1075,N_153,N_146);
xor U1076 (N_1076,N_380,N_112);
xor U1077 (N_1077,N_537,N_58);
xor U1078 (N_1078,N_338,N_77);
or U1079 (N_1079,N_138,N_124);
nor U1080 (N_1080,N_386,N_401);
or U1081 (N_1081,N_597,N_554);
nor U1082 (N_1082,N_28,N_136);
nand U1083 (N_1083,N_575,N_468);
or U1084 (N_1084,N_235,N_127);
nand U1085 (N_1085,N_441,N_127);
xnor U1086 (N_1086,N_66,N_527);
and U1087 (N_1087,N_456,N_599);
nand U1088 (N_1088,N_319,N_202);
nand U1089 (N_1089,N_16,N_260);
xor U1090 (N_1090,N_17,N_4);
and U1091 (N_1091,N_568,N_251);
nand U1092 (N_1092,N_395,N_88);
or U1093 (N_1093,N_139,N_50);
xor U1094 (N_1094,N_418,N_582);
nor U1095 (N_1095,N_565,N_389);
nor U1096 (N_1096,N_383,N_573);
nor U1097 (N_1097,N_425,N_11);
and U1098 (N_1098,N_245,N_424);
nand U1099 (N_1099,N_43,N_141);
nor U1100 (N_1100,N_306,N_373);
or U1101 (N_1101,N_39,N_376);
and U1102 (N_1102,N_159,N_164);
xor U1103 (N_1103,N_502,N_183);
xnor U1104 (N_1104,N_341,N_56);
nand U1105 (N_1105,N_422,N_512);
nand U1106 (N_1106,N_435,N_549);
and U1107 (N_1107,N_123,N_327);
xnor U1108 (N_1108,N_88,N_26);
and U1109 (N_1109,N_404,N_68);
and U1110 (N_1110,N_591,N_401);
nand U1111 (N_1111,N_67,N_118);
nor U1112 (N_1112,N_350,N_323);
nand U1113 (N_1113,N_4,N_70);
and U1114 (N_1114,N_63,N_399);
nor U1115 (N_1115,N_132,N_434);
nand U1116 (N_1116,N_533,N_531);
xor U1117 (N_1117,N_311,N_16);
and U1118 (N_1118,N_334,N_277);
and U1119 (N_1119,N_303,N_416);
nor U1120 (N_1120,N_131,N_192);
nor U1121 (N_1121,N_169,N_472);
and U1122 (N_1122,N_575,N_550);
and U1123 (N_1123,N_202,N_541);
nand U1124 (N_1124,N_156,N_68);
or U1125 (N_1125,N_555,N_151);
or U1126 (N_1126,N_69,N_364);
or U1127 (N_1127,N_401,N_555);
or U1128 (N_1128,N_321,N_88);
nor U1129 (N_1129,N_281,N_105);
or U1130 (N_1130,N_83,N_158);
nor U1131 (N_1131,N_234,N_315);
nor U1132 (N_1132,N_570,N_518);
nand U1133 (N_1133,N_355,N_531);
nor U1134 (N_1134,N_106,N_580);
nor U1135 (N_1135,N_103,N_104);
and U1136 (N_1136,N_483,N_249);
xnor U1137 (N_1137,N_74,N_481);
and U1138 (N_1138,N_236,N_349);
or U1139 (N_1139,N_260,N_175);
or U1140 (N_1140,N_133,N_60);
nand U1141 (N_1141,N_156,N_288);
or U1142 (N_1142,N_106,N_154);
xnor U1143 (N_1143,N_447,N_333);
or U1144 (N_1144,N_310,N_438);
xnor U1145 (N_1145,N_336,N_594);
or U1146 (N_1146,N_204,N_217);
xnor U1147 (N_1147,N_421,N_178);
and U1148 (N_1148,N_595,N_482);
or U1149 (N_1149,N_12,N_112);
nand U1150 (N_1150,N_59,N_563);
and U1151 (N_1151,N_502,N_389);
nor U1152 (N_1152,N_72,N_366);
and U1153 (N_1153,N_327,N_200);
nor U1154 (N_1154,N_30,N_12);
nand U1155 (N_1155,N_69,N_199);
nand U1156 (N_1156,N_290,N_401);
xnor U1157 (N_1157,N_114,N_20);
nor U1158 (N_1158,N_17,N_445);
xor U1159 (N_1159,N_587,N_380);
nand U1160 (N_1160,N_112,N_243);
and U1161 (N_1161,N_448,N_37);
xor U1162 (N_1162,N_246,N_466);
nand U1163 (N_1163,N_359,N_463);
nand U1164 (N_1164,N_30,N_264);
or U1165 (N_1165,N_83,N_431);
xnor U1166 (N_1166,N_494,N_45);
or U1167 (N_1167,N_32,N_0);
nor U1168 (N_1168,N_198,N_167);
xnor U1169 (N_1169,N_16,N_326);
xnor U1170 (N_1170,N_596,N_149);
xor U1171 (N_1171,N_463,N_258);
nor U1172 (N_1172,N_389,N_559);
and U1173 (N_1173,N_432,N_232);
nor U1174 (N_1174,N_465,N_577);
and U1175 (N_1175,N_316,N_526);
nor U1176 (N_1176,N_169,N_322);
and U1177 (N_1177,N_392,N_129);
or U1178 (N_1178,N_85,N_75);
nand U1179 (N_1179,N_578,N_0);
nand U1180 (N_1180,N_402,N_16);
xor U1181 (N_1181,N_253,N_106);
and U1182 (N_1182,N_68,N_195);
nor U1183 (N_1183,N_31,N_48);
or U1184 (N_1184,N_281,N_361);
xnor U1185 (N_1185,N_461,N_168);
or U1186 (N_1186,N_421,N_529);
xor U1187 (N_1187,N_556,N_520);
nand U1188 (N_1188,N_520,N_463);
or U1189 (N_1189,N_570,N_126);
or U1190 (N_1190,N_99,N_341);
nand U1191 (N_1191,N_423,N_169);
nand U1192 (N_1192,N_17,N_467);
nand U1193 (N_1193,N_160,N_145);
and U1194 (N_1194,N_538,N_28);
and U1195 (N_1195,N_298,N_579);
and U1196 (N_1196,N_558,N_385);
xor U1197 (N_1197,N_50,N_399);
or U1198 (N_1198,N_246,N_170);
or U1199 (N_1199,N_528,N_379);
nand U1200 (N_1200,N_1172,N_676);
nor U1201 (N_1201,N_1088,N_1198);
or U1202 (N_1202,N_682,N_653);
nor U1203 (N_1203,N_940,N_689);
nor U1204 (N_1204,N_741,N_911);
xor U1205 (N_1205,N_1097,N_1092);
or U1206 (N_1206,N_783,N_1114);
xor U1207 (N_1207,N_946,N_1080);
and U1208 (N_1208,N_810,N_996);
and U1209 (N_1209,N_821,N_842);
nor U1210 (N_1210,N_883,N_1169);
nor U1211 (N_1211,N_879,N_920);
nand U1212 (N_1212,N_1012,N_1022);
nand U1213 (N_1213,N_975,N_872);
and U1214 (N_1214,N_1143,N_745);
xnor U1215 (N_1215,N_943,N_750);
nor U1216 (N_1216,N_933,N_1007);
nand U1217 (N_1217,N_735,N_812);
and U1218 (N_1218,N_1094,N_1189);
nor U1219 (N_1219,N_1133,N_944);
nand U1220 (N_1220,N_1016,N_966);
nor U1221 (N_1221,N_792,N_1112);
or U1222 (N_1222,N_997,N_774);
and U1223 (N_1223,N_1194,N_1176);
and U1224 (N_1224,N_731,N_748);
nor U1225 (N_1225,N_992,N_804);
nand U1226 (N_1226,N_727,N_611);
nor U1227 (N_1227,N_801,N_712);
nor U1228 (N_1228,N_695,N_616);
nand U1229 (N_1229,N_891,N_1127);
and U1230 (N_1230,N_781,N_893);
xor U1231 (N_1231,N_1170,N_962);
and U1232 (N_1232,N_818,N_838);
and U1233 (N_1233,N_1062,N_1124);
and U1234 (N_1234,N_765,N_1011);
and U1235 (N_1235,N_1180,N_1183);
nand U1236 (N_1236,N_656,N_779);
xor U1237 (N_1237,N_685,N_1049);
nor U1238 (N_1238,N_1178,N_910);
nor U1239 (N_1239,N_1041,N_754);
xnor U1240 (N_1240,N_699,N_669);
xnor U1241 (N_1241,N_1040,N_841);
nand U1242 (N_1242,N_1024,N_1017);
nor U1243 (N_1243,N_1069,N_915);
nand U1244 (N_1244,N_832,N_1056);
xnor U1245 (N_1245,N_967,N_854);
nand U1246 (N_1246,N_925,N_899);
nand U1247 (N_1247,N_850,N_973);
nor U1248 (N_1248,N_835,N_787);
nor U1249 (N_1249,N_1038,N_683);
nor U1250 (N_1250,N_776,N_980);
nor U1251 (N_1251,N_1125,N_620);
nand U1252 (N_1252,N_937,N_717);
and U1253 (N_1253,N_1005,N_1117);
or U1254 (N_1254,N_635,N_1000);
or U1255 (N_1255,N_797,N_1107);
and U1256 (N_1256,N_789,N_874);
and U1257 (N_1257,N_978,N_723);
or U1258 (N_1258,N_982,N_1013);
or U1259 (N_1259,N_1050,N_619);
and U1260 (N_1260,N_896,N_1009);
xnor U1261 (N_1261,N_941,N_607);
or U1262 (N_1262,N_1190,N_860);
nor U1263 (N_1263,N_1028,N_672);
xnor U1264 (N_1264,N_710,N_684);
nor U1265 (N_1265,N_953,N_1126);
xnor U1266 (N_1266,N_848,N_858);
or U1267 (N_1267,N_708,N_764);
nand U1268 (N_1268,N_1046,N_746);
and U1269 (N_1269,N_959,N_831);
nand U1270 (N_1270,N_800,N_756);
xor U1271 (N_1271,N_1100,N_1149);
nor U1272 (N_1272,N_1096,N_809);
nand U1273 (N_1273,N_785,N_788);
nor U1274 (N_1274,N_1191,N_798);
or U1275 (N_1275,N_1072,N_903);
nand U1276 (N_1276,N_902,N_930);
and U1277 (N_1277,N_1175,N_1104);
nor U1278 (N_1278,N_1150,N_771);
nand U1279 (N_1279,N_970,N_1071);
or U1280 (N_1280,N_637,N_1047);
or U1281 (N_1281,N_1018,N_1148);
nand U1282 (N_1282,N_1023,N_948);
nor U1283 (N_1283,N_766,N_1098);
xor U1284 (N_1284,N_987,N_1177);
and U1285 (N_1285,N_752,N_1020);
nor U1286 (N_1286,N_968,N_906);
or U1287 (N_1287,N_989,N_1137);
nor U1288 (N_1288,N_759,N_836);
or U1289 (N_1289,N_1151,N_1109);
nand U1290 (N_1290,N_1136,N_1052);
and U1291 (N_1291,N_1043,N_972);
nand U1292 (N_1292,N_1179,N_998);
nor U1293 (N_1293,N_927,N_1061);
xor U1294 (N_1294,N_1037,N_782);
nand U1295 (N_1295,N_1131,N_839);
nand U1296 (N_1296,N_626,N_868);
nand U1297 (N_1297,N_627,N_1087);
and U1298 (N_1298,N_844,N_816);
nand U1299 (N_1299,N_995,N_1103);
or U1300 (N_1300,N_734,N_887);
and U1301 (N_1301,N_621,N_1078);
nor U1302 (N_1302,N_612,N_659);
nor U1303 (N_1303,N_1010,N_647);
nor U1304 (N_1304,N_665,N_608);
nand U1305 (N_1305,N_675,N_743);
nor U1306 (N_1306,N_1164,N_681);
and U1307 (N_1307,N_1014,N_1066);
xnor U1308 (N_1308,N_1030,N_1161);
nand U1309 (N_1309,N_1168,N_956);
or U1310 (N_1310,N_852,N_1163);
nor U1311 (N_1311,N_863,N_739);
nand U1312 (N_1312,N_965,N_613);
and U1313 (N_1313,N_871,N_1081);
nand U1314 (N_1314,N_606,N_1110);
and U1315 (N_1315,N_805,N_691);
nor U1316 (N_1316,N_916,N_1145);
xor U1317 (N_1317,N_1075,N_1188);
xnor U1318 (N_1318,N_870,N_722);
and U1319 (N_1319,N_737,N_1082);
and U1320 (N_1320,N_1048,N_753);
nor U1321 (N_1321,N_640,N_859);
and U1322 (N_1322,N_985,N_904);
and U1323 (N_1323,N_677,N_952);
nor U1324 (N_1324,N_964,N_1006);
xnor U1325 (N_1325,N_1058,N_668);
nor U1326 (N_1326,N_1192,N_1002);
nor U1327 (N_1327,N_1051,N_977);
nor U1328 (N_1328,N_1157,N_1174);
xor U1329 (N_1329,N_811,N_740);
nor U1330 (N_1330,N_924,N_1057);
nor U1331 (N_1331,N_724,N_882);
nor U1332 (N_1332,N_1134,N_630);
or U1333 (N_1333,N_654,N_690);
nand U1334 (N_1334,N_1003,N_815);
xor U1335 (N_1335,N_849,N_875);
nand U1336 (N_1336,N_971,N_813);
xnor U1337 (N_1337,N_846,N_945);
xor U1338 (N_1338,N_905,N_1166);
nor U1339 (N_1339,N_625,N_999);
or U1340 (N_1340,N_1102,N_1029);
xnor U1341 (N_1341,N_921,N_1106);
and U1342 (N_1342,N_1154,N_961);
nand U1343 (N_1343,N_778,N_796);
xnor U1344 (N_1344,N_707,N_725);
nor U1345 (N_1345,N_1132,N_803);
and U1346 (N_1346,N_715,N_1083);
and U1347 (N_1347,N_762,N_826);
xnor U1348 (N_1348,N_622,N_709);
and U1349 (N_1349,N_802,N_888);
and U1350 (N_1350,N_628,N_1152);
nand U1351 (N_1351,N_917,N_751);
xor U1352 (N_1352,N_876,N_929);
and U1353 (N_1353,N_1021,N_742);
or U1354 (N_1354,N_1077,N_807);
or U1355 (N_1355,N_1036,N_869);
xnor U1356 (N_1356,N_960,N_909);
and U1357 (N_1357,N_991,N_856);
xnor U1358 (N_1358,N_827,N_678);
xor U1359 (N_1359,N_958,N_1095);
or U1360 (N_1360,N_674,N_901);
or U1361 (N_1361,N_1032,N_704);
nand U1362 (N_1362,N_733,N_918);
nand U1363 (N_1363,N_655,N_892);
xnor U1364 (N_1364,N_913,N_794);
and U1365 (N_1365,N_729,N_1019);
xnor U1366 (N_1366,N_763,N_866);
or U1367 (N_1367,N_1001,N_772);
and U1368 (N_1368,N_889,N_825);
or U1369 (N_1369,N_760,N_954);
nor U1370 (N_1370,N_862,N_1027);
xor U1371 (N_1371,N_1045,N_664);
nand U1372 (N_1372,N_719,N_749);
and U1373 (N_1373,N_736,N_713);
xnor U1374 (N_1374,N_1119,N_702);
nand U1375 (N_1375,N_926,N_663);
nand U1376 (N_1376,N_650,N_658);
nand U1377 (N_1377,N_1173,N_1186);
nor U1378 (N_1378,N_1090,N_614);
nor U1379 (N_1379,N_1146,N_636);
and U1380 (N_1380,N_609,N_1093);
nor U1381 (N_1381,N_1113,N_932);
nor U1382 (N_1382,N_963,N_738);
xor U1383 (N_1383,N_728,N_651);
and U1384 (N_1384,N_1064,N_617);
or U1385 (N_1385,N_806,N_1167);
and U1386 (N_1386,N_857,N_1115);
or U1387 (N_1387,N_1084,N_657);
nor U1388 (N_1388,N_824,N_928);
xor U1389 (N_1389,N_652,N_1073);
or U1390 (N_1390,N_1139,N_755);
or U1391 (N_1391,N_974,N_1141);
and U1392 (N_1392,N_720,N_1197);
or U1393 (N_1393,N_1122,N_679);
nor U1394 (N_1394,N_885,N_829);
and U1395 (N_1395,N_984,N_853);
xnor U1396 (N_1396,N_1065,N_604);
nor U1397 (N_1397,N_747,N_1147);
nor U1398 (N_1398,N_1160,N_1116);
xor U1399 (N_1399,N_934,N_670);
and U1400 (N_1400,N_808,N_1158);
nand U1401 (N_1401,N_979,N_730);
and U1402 (N_1402,N_1079,N_1060);
and U1403 (N_1403,N_895,N_703);
xnor U1404 (N_1404,N_1015,N_923);
or U1405 (N_1405,N_908,N_649);
nor U1406 (N_1406,N_1181,N_680);
xor U1407 (N_1407,N_897,N_1053);
nor U1408 (N_1408,N_942,N_830);
or U1409 (N_1409,N_988,N_957);
and U1410 (N_1410,N_912,N_1165);
nand U1411 (N_1411,N_744,N_1108);
and U1412 (N_1412,N_634,N_1121);
xor U1413 (N_1413,N_851,N_768);
or U1414 (N_1414,N_1063,N_983);
nor U1415 (N_1415,N_855,N_981);
xnor U1416 (N_1416,N_757,N_600);
nand U1417 (N_1417,N_1034,N_1123);
nor U1418 (N_1418,N_721,N_1140);
nor U1419 (N_1419,N_666,N_994);
and U1420 (N_1420,N_890,N_791);
xnor U1421 (N_1421,N_1031,N_873);
xnor U1422 (N_1422,N_688,N_633);
or U1423 (N_1423,N_1156,N_1026);
nand U1424 (N_1424,N_645,N_1111);
nand U1425 (N_1425,N_775,N_706);
and U1426 (N_1426,N_814,N_769);
xor U1427 (N_1427,N_1155,N_1135);
nand U1428 (N_1428,N_898,N_1130);
nor U1429 (N_1429,N_1008,N_990);
xor U1430 (N_1430,N_714,N_732);
nor U1431 (N_1431,N_777,N_1099);
and U1432 (N_1432,N_716,N_641);
and U1433 (N_1433,N_1162,N_711);
or U1434 (N_1434,N_881,N_955);
and U1435 (N_1435,N_1035,N_793);
and U1436 (N_1436,N_845,N_864);
xnor U1437 (N_1437,N_1182,N_938);
nand U1438 (N_1438,N_660,N_820);
nand U1439 (N_1439,N_692,N_1044);
or U1440 (N_1440,N_865,N_726);
and U1441 (N_1441,N_799,N_605);
nor U1442 (N_1442,N_914,N_615);
xor U1443 (N_1443,N_1074,N_758);
or U1444 (N_1444,N_632,N_700);
nor U1445 (N_1445,N_610,N_1195);
xnor U1446 (N_1446,N_642,N_837);
nor U1447 (N_1447,N_1101,N_878);
nand U1448 (N_1448,N_1039,N_828);
and U1449 (N_1449,N_833,N_1199);
and U1450 (N_1450,N_786,N_986);
xnor U1451 (N_1451,N_1196,N_947);
and U1452 (N_1452,N_935,N_1091);
nand U1453 (N_1453,N_687,N_705);
xnor U1454 (N_1454,N_1042,N_843);
and U1455 (N_1455,N_1129,N_907);
xnor U1456 (N_1456,N_639,N_1144);
and U1457 (N_1457,N_819,N_894);
nand U1458 (N_1458,N_1153,N_939);
nor U1459 (N_1459,N_1076,N_1054);
xnor U1460 (N_1460,N_773,N_623);
xnor U1461 (N_1461,N_861,N_1004);
nand U1462 (N_1462,N_693,N_1159);
xnor U1463 (N_1463,N_817,N_1105);
xor U1464 (N_1464,N_780,N_1171);
nand U1465 (N_1465,N_1120,N_880);
nor U1466 (N_1466,N_1128,N_701);
nand U1467 (N_1467,N_1068,N_644);
and U1468 (N_1468,N_949,N_618);
xnor U1469 (N_1469,N_686,N_718);
and U1470 (N_1470,N_1085,N_671);
nor U1471 (N_1471,N_1089,N_886);
or U1472 (N_1472,N_1187,N_840);
and U1473 (N_1473,N_696,N_1070);
and U1474 (N_1474,N_936,N_1033);
nor U1475 (N_1475,N_1138,N_648);
or U1476 (N_1476,N_922,N_698);
or U1477 (N_1477,N_667,N_643);
or U1478 (N_1478,N_822,N_1067);
or U1479 (N_1479,N_790,N_1142);
or U1480 (N_1480,N_624,N_1025);
nand U1481 (N_1481,N_1059,N_823);
xor U1482 (N_1482,N_761,N_770);
nor U1483 (N_1483,N_950,N_601);
xor U1484 (N_1484,N_784,N_919);
xor U1485 (N_1485,N_1055,N_661);
nor U1486 (N_1486,N_976,N_969);
nand U1487 (N_1487,N_629,N_767);
and U1488 (N_1488,N_1185,N_867);
nand U1489 (N_1489,N_694,N_638);
nand U1490 (N_1490,N_900,N_1118);
xor U1491 (N_1491,N_673,N_847);
xor U1492 (N_1492,N_931,N_602);
or U1493 (N_1493,N_1193,N_834);
and U1494 (N_1494,N_951,N_603);
nand U1495 (N_1495,N_697,N_1184);
xor U1496 (N_1496,N_795,N_662);
xor U1497 (N_1497,N_646,N_993);
and U1498 (N_1498,N_884,N_1086);
xnor U1499 (N_1499,N_877,N_631);
or U1500 (N_1500,N_733,N_1005);
and U1501 (N_1501,N_672,N_1135);
nor U1502 (N_1502,N_813,N_928);
nand U1503 (N_1503,N_735,N_1070);
or U1504 (N_1504,N_605,N_957);
and U1505 (N_1505,N_964,N_1176);
or U1506 (N_1506,N_1101,N_807);
nor U1507 (N_1507,N_648,N_1144);
or U1508 (N_1508,N_680,N_829);
nand U1509 (N_1509,N_705,N_1115);
or U1510 (N_1510,N_1195,N_701);
nor U1511 (N_1511,N_1045,N_1031);
nand U1512 (N_1512,N_691,N_1153);
or U1513 (N_1513,N_762,N_1085);
nand U1514 (N_1514,N_800,N_1027);
and U1515 (N_1515,N_611,N_1001);
nand U1516 (N_1516,N_821,N_995);
nand U1517 (N_1517,N_869,N_625);
or U1518 (N_1518,N_1121,N_914);
nand U1519 (N_1519,N_988,N_604);
nand U1520 (N_1520,N_686,N_997);
and U1521 (N_1521,N_1157,N_1164);
or U1522 (N_1522,N_986,N_869);
nor U1523 (N_1523,N_1059,N_839);
or U1524 (N_1524,N_1076,N_1129);
xnor U1525 (N_1525,N_1140,N_840);
nor U1526 (N_1526,N_710,N_1021);
or U1527 (N_1527,N_1049,N_734);
and U1528 (N_1528,N_897,N_875);
xnor U1529 (N_1529,N_916,N_808);
nand U1530 (N_1530,N_944,N_1008);
nand U1531 (N_1531,N_950,N_1010);
nand U1532 (N_1532,N_1152,N_746);
and U1533 (N_1533,N_1035,N_821);
nor U1534 (N_1534,N_1162,N_656);
or U1535 (N_1535,N_1133,N_796);
and U1536 (N_1536,N_603,N_629);
nand U1537 (N_1537,N_796,N_645);
and U1538 (N_1538,N_1194,N_856);
nor U1539 (N_1539,N_872,N_646);
xor U1540 (N_1540,N_1026,N_1037);
and U1541 (N_1541,N_1186,N_1058);
and U1542 (N_1542,N_1156,N_642);
and U1543 (N_1543,N_994,N_1048);
and U1544 (N_1544,N_604,N_688);
or U1545 (N_1545,N_1190,N_1197);
and U1546 (N_1546,N_1087,N_754);
and U1547 (N_1547,N_1051,N_929);
xor U1548 (N_1548,N_1077,N_1192);
or U1549 (N_1549,N_711,N_676);
nor U1550 (N_1550,N_1015,N_991);
nand U1551 (N_1551,N_759,N_735);
nor U1552 (N_1552,N_1077,N_780);
nand U1553 (N_1553,N_895,N_1182);
and U1554 (N_1554,N_777,N_749);
or U1555 (N_1555,N_1152,N_743);
nand U1556 (N_1556,N_1067,N_933);
nand U1557 (N_1557,N_802,N_781);
or U1558 (N_1558,N_780,N_1132);
xor U1559 (N_1559,N_949,N_1142);
and U1560 (N_1560,N_647,N_815);
or U1561 (N_1561,N_902,N_613);
xor U1562 (N_1562,N_968,N_817);
and U1563 (N_1563,N_1002,N_951);
xor U1564 (N_1564,N_974,N_662);
xor U1565 (N_1565,N_916,N_942);
or U1566 (N_1566,N_766,N_929);
xor U1567 (N_1567,N_962,N_1072);
and U1568 (N_1568,N_715,N_1185);
or U1569 (N_1569,N_683,N_1179);
nor U1570 (N_1570,N_849,N_870);
and U1571 (N_1571,N_1021,N_1092);
nand U1572 (N_1572,N_1165,N_1131);
nand U1573 (N_1573,N_809,N_646);
nand U1574 (N_1574,N_701,N_936);
nand U1575 (N_1575,N_948,N_754);
nor U1576 (N_1576,N_801,N_980);
and U1577 (N_1577,N_918,N_1060);
or U1578 (N_1578,N_711,N_826);
nor U1579 (N_1579,N_1111,N_880);
nor U1580 (N_1580,N_1120,N_1009);
nor U1581 (N_1581,N_964,N_870);
xnor U1582 (N_1582,N_865,N_1084);
or U1583 (N_1583,N_801,N_674);
and U1584 (N_1584,N_1142,N_887);
nor U1585 (N_1585,N_717,N_936);
nor U1586 (N_1586,N_1122,N_628);
and U1587 (N_1587,N_1068,N_998);
nor U1588 (N_1588,N_796,N_847);
nor U1589 (N_1589,N_619,N_848);
and U1590 (N_1590,N_1176,N_971);
nor U1591 (N_1591,N_949,N_843);
or U1592 (N_1592,N_734,N_862);
and U1593 (N_1593,N_1078,N_955);
or U1594 (N_1594,N_793,N_1122);
nor U1595 (N_1595,N_804,N_979);
nor U1596 (N_1596,N_658,N_826);
nand U1597 (N_1597,N_778,N_677);
xor U1598 (N_1598,N_1097,N_1008);
and U1599 (N_1599,N_925,N_1137);
and U1600 (N_1600,N_664,N_788);
and U1601 (N_1601,N_820,N_1090);
nand U1602 (N_1602,N_1169,N_817);
nand U1603 (N_1603,N_1129,N_696);
xor U1604 (N_1604,N_787,N_1156);
and U1605 (N_1605,N_771,N_1169);
xor U1606 (N_1606,N_994,N_606);
or U1607 (N_1607,N_931,N_1190);
xnor U1608 (N_1608,N_777,N_896);
nand U1609 (N_1609,N_617,N_844);
nor U1610 (N_1610,N_1082,N_1010);
and U1611 (N_1611,N_1110,N_764);
nand U1612 (N_1612,N_1009,N_760);
nand U1613 (N_1613,N_700,N_857);
and U1614 (N_1614,N_730,N_880);
nand U1615 (N_1615,N_1113,N_846);
xor U1616 (N_1616,N_842,N_1035);
nand U1617 (N_1617,N_725,N_1054);
or U1618 (N_1618,N_905,N_878);
or U1619 (N_1619,N_1066,N_1075);
nor U1620 (N_1620,N_902,N_1174);
or U1621 (N_1621,N_936,N_1185);
or U1622 (N_1622,N_868,N_1095);
nand U1623 (N_1623,N_837,N_1168);
or U1624 (N_1624,N_1049,N_1041);
nand U1625 (N_1625,N_762,N_888);
xnor U1626 (N_1626,N_659,N_1197);
and U1627 (N_1627,N_1036,N_1009);
xor U1628 (N_1628,N_1067,N_1127);
nor U1629 (N_1629,N_1117,N_607);
and U1630 (N_1630,N_1008,N_735);
nand U1631 (N_1631,N_836,N_668);
nor U1632 (N_1632,N_891,N_1021);
xor U1633 (N_1633,N_696,N_621);
and U1634 (N_1634,N_1008,N_806);
nor U1635 (N_1635,N_769,N_1180);
nor U1636 (N_1636,N_1082,N_995);
or U1637 (N_1637,N_835,N_1187);
nor U1638 (N_1638,N_1059,N_659);
nand U1639 (N_1639,N_698,N_1198);
and U1640 (N_1640,N_1092,N_776);
nand U1641 (N_1641,N_783,N_904);
and U1642 (N_1642,N_783,N_743);
xor U1643 (N_1643,N_638,N_862);
and U1644 (N_1644,N_902,N_804);
or U1645 (N_1645,N_1175,N_618);
nor U1646 (N_1646,N_787,N_832);
nor U1647 (N_1647,N_738,N_998);
nor U1648 (N_1648,N_857,N_1028);
xor U1649 (N_1649,N_1126,N_730);
nor U1650 (N_1650,N_895,N_1108);
and U1651 (N_1651,N_644,N_846);
or U1652 (N_1652,N_911,N_1198);
xor U1653 (N_1653,N_1042,N_709);
nand U1654 (N_1654,N_1159,N_714);
xor U1655 (N_1655,N_928,N_795);
xnor U1656 (N_1656,N_888,N_963);
and U1657 (N_1657,N_1050,N_729);
xor U1658 (N_1658,N_1148,N_726);
and U1659 (N_1659,N_693,N_1085);
nand U1660 (N_1660,N_876,N_1064);
or U1661 (N_1661,N_950,N_973);
or U1662 (N_1662,N_897,N_755);
nand U1663 (N_1663,N_831,N_634);
nand U1664 (N_1664,N_1172,N_975);
xor U1665 (N_1665,N_988,N_761);
or U1666 (N_1666,N_823,N_941);
and U1667 (N_1667,N_961,N_835);
nand U1668 (N_1668,N_854,N_887);
or U1669 (N_1669,N_724,N_916);
or U1670 (N_1670,N_901,N_1012);
and U1671 (N_1671,N_1129,N_1162);
or U1672 (N_1672,N_1015,N_1185);
or U1673 (N_1673,N_673,N_859);
or U1674 (N_1674,N_1058,N_736);
nand U1675 (N_1675,N_1182,N_973);
nor U1676 (N_1676,N_1122,N_1121);
or U1677 (N_1677,N_1112,N_856);
nor U1678 (N_1678,N_717,N_806);
or U1679 (N_1679,N_822,N_1155);
xor U1680 (N_1680,N_845,N_812);
nand U1681 (N_1681,N_1021,N_991);
nand U1682 (N_1682,N_1008,N_1172);
xor U1683 (N_1683,N_839,N_883);
nor U1684 (N_1684,N_994,N_651);
and U1685 (N_1685,N_1058,N_1106);
xnor U1686 (N_1686,N_952,N_962);
nor U1687 (N_1687,N_833,N_873);
and U1688 (N_1688,N_1194,N_903);
xnor U1689 (N_1689,N_676,N_644);
or U1690 (N_1690,N_693,N_810);
or U1691 (N_1691,N_936,N_645);
or U1692 (N_1692,N_911,N_899);
nand U1693 (N_1693,N_614,N_868);
nand U1694 (N_1694,N_997,N_710);
xor U1695 (N_1695,N_901,N_1098);
or U1696 (N_1696,N_771,N_1043);
and U1697 (N_1697,N_846,N_752);
nand U1698 (N_1698,N_1039,N_773);
xnor U1699 (N_1699,N_1150,N_965);
or U1700 (N_1700,N_1152,N_1192);
nor U1701 (N_1701,N_705,N_911);
or U1702 (N_1702,N_1036,N_622);
nor U1703 (N_1703,N_1153,N_832);
nor U1704 (N_1704,N_1199,N_1046);
or U1705 (N_1705,N_930,N_895);
nor U1706 (N_1706,N_1188,N_755);
and U1707 (N_1707,N_954,N_1163);
or U1708 (N_1708,N_671,N_815);
nor U1709 (N_1709,N_1049,N_836);
nor U1710 (N_1710,N_1139,N_1103);
xor U1711 (N_1711,N_616,N_717);
nand U1712 (N_1712,N_1001,N_1124);
and U1713 (N_1713,N_703,N_728);
nor U1714 (N_1714,N_1080,N_928);
xor U1715 (N_1715,N_715,N_1087);
and U1716 (N_1716,N_1068,N_760);
xnor U1717 (N_1717,N_819,N_1191);
or U1718 (N_1718,N_665,N_1135);
nand U1719 (N_1719,N_1037,N_844);
or U1720 (N_1720,N_1178,N_1074);
nor U1721 (N_1721,N_883,N_603);
xor U1722 (N_1722,N_837,N_1138);
nor U1723 (N_1723,N_882,N_877);
nor U1724 (N_1724,N_925,N_1152);
nand U1725 (N_1725,N_951,N_895);
and U1726 (N_1726,N_1182,N_865);
xnor U1727 (N_1727,N_759,N_1197);
or U1728 (N_1728,N_1148,N_949);
nor U1729 (N_1729,N_883,N_879);
nand U1730 (N_1730,N_801,N_727);
nand U1731 (N_1731,N_1139,N_761);
xor U1732 (N_1732,N_1102,N_1126);
nor U1733 (N_1733,N_787,N_801);
nor U1734 (N_1734,N_701,N_1081);
and U1735 (N_1735,N_932,N_1080);
or U1736 (N_1736,N_902,N_1081);
nand U1737 (N_1737,N_954,N_1005);
xnor U1738 (N_1738,N_1013,N_1198);
nor U1739 (N_1739,N_806,N_849);
or U1740 (N_1740,N_968,N_616);
xnor U1741 (N_1741,N_962,N_794);
nor U1742 (N_1742,N_1107,N_885);
nand U1743 (N_1743,N_1151,N_709);
xnor U1744 (N_1744,N_723,N_940);
xor U1745 (N_1745,N_737,N_1198);
and U1746 (N_1746,N_962,N_648);
and U1747 (N_1747,N_937,N_783);
nand U1748 (N_1748,N_1060,N_847);
and U1749 (N_1749,N_1006,N_1090);
nor U1750 (N_1750,N_1128,N_832);
or U1751 (N_1751,N_901,N_1151);
or U1752 (N_1752,N_710,N_1015);
or U1753 (N_1753,N_904,N_681);
nor U1754 (N_1754,N_623,N_613);
nor U1755 (N_1755,N_722,N_720);
xor U1756 (N_1756,N_621,N_1048);
nand U1757 (N_1757,N_828,N_869);
nand U1758 (N_1758,N_1194,N_1081);
xor U1759 (N_1759,N_909,N_1041);
xnor U1760 (N_1760,N_661,N_1191);
nand U1761 (N_1761,N_819,N_1032);
and U1762 (N_1762,N_751,N_995);
nor U1763 (N_1763,N_1115,N_835);
xnor U1764 (N_1764,N_886,N_896);
nand U1765 (N_1765,N_616,N_1040);
nand U1766 (N_1766,N_1183,N_611);
nor U1767 (N_1767,N_832,N_1052);
nor U1768 (N_1768,N_1170,N_1146);
nor U1769 (N_1769,N_1199,N_777);
and U1770 (N_1770,N_1164,N_1159);
xor U1771 (N_1771,N_1043,N_1029);
nor U1772 (N_1772,N_993,N_1073);
nand U1773 (N_1773,N_779,N_958);
nand U1774 (N_1774,N_870,N_610);
nor U1775 (N_1775,N_1163,N_1181);
or U1776 (N_1776,N_1088,N_894);
or U1777 (N_1777,N_1138,N_604);
nor U1778 (N_1778,N_877,N_1129);
nand U1779 (N_1779,N_1006,N_1049);
nand U1780 (N_1780,N_789,N_1036);
nand U1781 (N_1781,N_1128,N_720);
and U1782 (N_1782,N_1045,N_617);
and U1783 (N_1783,N_811,N_869);
nor U1784 (N_1784,N_682,N_900);
nor U1785 (N_1785,N_1112,N_1151);
xor U1786 (N_1786,N_1050,N_820);
xor U1787 (N_1787,N_816,N_612);
nand U1788 (N_1788,N_926,N_994);
xor U1789 (N_1789,N_1125,N_838);
nor U1790 (N_1790,N_878,N_1082);
nor U1791 (N_1791,N_1195,N_720);
and U1792 (N_1792,N_1170,N_813);
nor U1793 (N_1793,N_728,N_881);
xnor U1794 (N_1794,N_1186,N_1100);
xor U1795 (N_1795,N_1159,N_793);
xnor U1796 (N_1796,N_1011,N_610);
and U1797 (N_1797,N_1022,N_1054);
nand U1798 (N_1798,N_790,N_643);
nor U1799 (N_1799,N_1106,N_941);
nand U1800 (N_1800,N_1273,N_1411);
nand U1801 (N_1801,N_1401,N_1288);
or U1802 (N_1802,N_1731,N_1278);
nand U1803 (N_1803,N_1769,N_1221);
nor U1804 (N_1804,N_1416,N_1762);
nor U1805 (N_1805,N_1452,N_1381);
nor U1806 (N_1806,N_1640,N_1241);
and U1807 (N_1807,N_1615,N_1689);
xor U1808 (N_1808,N_1705,N_1623);
nand U1809 (N_1809,N_1318,N_1342);
or U1810 (N_1810,N_1510,N_1584);
nand U1811 (N_1811,N_1287,N_1668);
nand U1812 (N_1812,N_1703,N_1414);
or U1813 (N_1813,N_1290,N_1561);
or U1814 (N_1814,N_1251,N_1530);
nor U1815 (N_1815,N_1574,N_1336);
nand U1816 (N_1816,N_1369,N_1490);
and U1817 (N_1817,N_1701,N_1215);
and U1818 (N_1818,N_1793,N_1432);
and U1819 (N_1819,N_1352,N_1461);
nor U1820 (N_1820,N_1613,N_1564);
and U1821 (N_1821,N_1473,N_1603);
nor U1822 (N_1822,N_1232,N_1317);
or U1823 (N_1823,N_1211,N_1737);
xnor U1824 (N_1824,N_1409,N_1524);
xor U1825 (N_1825,N_1738,N_1570);
or U1826 (N_1826,N_1298,N_1743);
or U1827 (N_1827,N_1760,N_1229);
xnor U1828 (N_1828,N_1258,N_1621);
xor U1829 (N_1829,N_1272,N_1755);
nor U1830 (N_1830,N_1670,N_1253);
xnor U1831 (N_1831,N_1263,N_1501);
and U1832 (N_1832,N_1223,N_1610);
or U1833 (N_1833,N_1388,N_1437);
xor U1834 (N_1834,N_1597,N_1467);
nor U1835 (N_1835,N_1474,N_1338);
and U1836 (N_1836,N_1697,N_1509);
nor U1837 (N_1837,N_1321,N_1683);
nand U1838 (N_1838,N_1325,N_1730);
or U1839 (N_1839,N_1377,N_1658);
or U1840 (N_1840,N_1227,N_1578);
xor U1841 (N_1841,N_1292,N_1442);
xnor U1842 (N_1842,N_1242,N_1711);
or U1843 (N_1843,N_1447,N_1572);
or U1844 (N_1844,N_1669,N_1312);
and U1845 (N_1845,N_1279,N_1596);
nand U1846 (N_1846,N_1780,N_1784);
and U1847 (N_1847,N_1218,N_1727);
nand U1848 (N_1848,N_1357,N_1671);
or U1849 (N_1849,N_1513,N_1492);
or U1850 (N_1850,N_1322,N_1706);
nor U1851 (N_1851,N_1376,N_1568);
xnor U1852 (N_1852,N_1247,N_1580);
or U1853 (N_1853,N_1331,N_1677);
xor U1854 (N_1854,N_1736,N_1694);
nor U1855 (N_1855,N_1546,N_1612);
nand U1856 (N_1856,N_1248,N_1750);
or U1857 (N_1857,N_1332,N_1339);
nand U1858 (N_1858,N_1499,N_1724);
nor U1859 (N_1859,N_1285,N_1310);
or U1860 (N_1860,N_1400,N_1631);
and U1861 (N_1861,N_1739,N_1773);
xnor U1862 (N_1862,N_1265,N_1764);
or U1863 (N_1863,N_1415,N_1240);
nand U1864 (N_1864,N_1632,N_1528);
nor U1865 (N_1865,N_1756,N_1741);
nand U1866 (N_1866,N_1373,N_1446);
xnor U1867 (N_1867,N_1491,N_1257);
and U1868 (N_1868,N_1494,N_1680);
nor U1869 (N_1869,N_1478,N_1255);
nor U1870 (N_1870,N_1348,N_1304);
xor U1871 (N_1871,N_1518,N_1544);
nor U1872 (N_1872,N_1767,N_1319);
or U1873 (N_1873,N_1485,N_1346);
nand U1874 (N_1874,N_1475,N_1709);
xnor U1875 (N_1875,N_1205,N_1606);
or U1876 (N_1876,N_1460,N_1324);
xor U1877 (N_1877,N_1626,N_1763);
nor U1878 (N_1878,N_1252,N_1291);
and U1879 (N_1879,N_1674,N_1207);
xor U1880 (N_1880,N_1673,N_1684);
nor U1881 (N_1881,N_1222,N_1563);
or U1882 (N_1882,N_1722,N_1779);
nand U1883 (N_1883,N_1462,N_1412);
nor U1884 (N_1884,N_1585,N_1430);
nand U1885 (N_1885,N_1386,N_1662);
and U1886 (N_1886,N_1483,N_1591);
nand U1887 (N_1887,N_1515,N_1542);
or U1888 (N_1888,N_1782,N_1519);
nand U1889 (N_1889,N_1387,N_1556);
or U1890 (N_1890,N_1320,N_1573);
xor U1891 (N_1891,N_1394,N_1696);
xor U1892 (N_1892,N_1308,N_1277);
xor U1893 (N_1893,N_1796,N_1487);
xor U1894 (N_1894,N_1708,N_1569);
and U1895 (N_1895,N_1233,N_1602);
or U1896 (N_1896,N_1758,N_1481);
nor U1897 (N_1897,N_1702,N_1350);
nand U1898 (N_1898,N_1629,N_1534);
and U1899 (N_1899,N_1700,N_1309);
nor U1900 (N_1900,N_1249,N_1482);
and U1901 (N_1901,N_1356,N_1374);
and U1902 (N_1902,N_1306,N_1307);
xnor U1903 (N_1903,N_1543,N_1666);
xor U1904 (N_1904,N_1679,N_1398);
xor U1905 (N_1905,N_1234,N_1567);
xnor U1906 (N_1906,N_1557,N_1653);
or U1907 (N_1907,N_1789,N_1450);
xor U1908 (N_1908,N_1728,N_1334);
nor U1909 (N_1909,N_1434,N_1548);
or U1910 (N_1910,N_1648,N_1345);
or U1911 (N_1911,N_1511,N_1766);
and U1912 (N_1912,N_1407,N_1641);
nand U1913 (N_1913,N_1270,N_1443);
nand U1914 (N_1914,N_1571,N_1707);
xnor U1915 (N_1915,N_1713,N_1391);
or U1916 (N_1916,N_1581,N_1379);
or U1917 (N_1917,N_1732,N_1425);
nand U1918 (N_1918,N_1347,N_1261);
and U1919 (N_1919,N_1419,N_1202);
nand U1920 (N_1920,N_1479,N_1370);
nand U1921 (N_1921,N_1704,N_1753);
or U1922 (N_1922,N_1665,N_1281);
nand U1923 (N_1923,N_1588,N_1343);
or U1924 (N_1924,N_1692,N_1436);
xnor U1925 (N_1925,N_1772,N_1271);
and U1926 (N_1926,N_1719,N_1260);
or U1927 (N_1927,N_1206,N_1405);
or U1928 (N_1928,N_1313,N_1403);
nor U1929 (N_1929,N_1533,N_1389);
or U1930 (N_1930,N_1344,N_1385);
nor U1931 (N_1931,N_1477,N_1372);
or U1932 (N_1932,N_1616,N_1231);
nand U1933 (N_1933,N_1451,N_1267);
and U1934 (N_1934,N_1687,N_1219);
nand U1935 (N_1935,N_1681,N_1775);
nand U1936 (N_1936,N_1504,N_1645);
and U1937 (N_1937,N_1341,N_1441);
nand U1938 (N_1938,N_1293,N_1204);
nand U1939 (N_1939,N_1274,N_1607);
and U1940 (N_1940,N_1327,N_1349);
or U1941 (N_1941,N_1362,N_1286);
xnor U1942 (N_1942,N_1250,N_1390);
and U1943 (N_1943,N_1335,N_1208);
nor U1944 (N_1944,N_1678,N_1733);
nor U1945 (N_1945,N_1651,N_1440);
nor U1946 (N_1946,N_1592,N_1686);
xor U1947 (N_1947,N_1470,N_1583);
nor U1948 (N_1948,N_1794,N_1685);
nand U1949 (N_1949,N_1459,N_1627);
xnor U1950 (N_1950,N_1551,N_1495);
nand U1951 (N_1951,N_1464,N_1355);
xnor U1952 (N_1952,N_1582,N_1695);
and U1953 (N_1953,N_1230,N_1224);
nand U1954 (N_1954,N_1471,N_1262);
or U1955 (N_1955,N_1783,N_1545);
and U1956 (N_1956,N_1466,N_1284);
or U1957 (N_1957,N_1295,N_1751);
xor U1958 (N_1958,N_1480,N_1406);
nor U1959 (N_1959,N_1566,N_1525);
nand U1960 (N_1960,N_1213,N_1531);
nand U1961 (N_1961,N_1646,N_1699);
nand U1962 (N_1962,N_1667,N_1489);
xor U1963 (N_1963,N_1595,N_1710);
or U1964 (N_1964,N_1516,N_1535);
nor U1965 (N_1965,N_1555,N_1747);
or U1966 (N_1966,N_1337,N_1484);
xor U1967 (N_1967,N_1601,N_1296);
nor U1968 (N_1968,N_1532,N_1550);
nand U1969 (N_1969,N_1380,N_1236);
xor U1970 (N_1970,N_1663,N_1560);
xnor U1971 (N_1971,N_1647,N_1468);
xnor U1972 (N_1972,N_1418,N_1417);
nand U1973 (N_1973,N_1778,N_1742);
nor U1974 (N_1974,N_1652,N_1774);
xnor U1975 (N_1975,N_1311,N_1426);
xor U1976 (N_1976,N_1365,N_1633);
nor U1977 (N_1977,N_1693,N_1740);
xnor U1978 (N_1978,N_1508,N_1517);
and U1979 (N_1979,N_1644,N_1453);
nor U1980 (N_1980,N_1675,N_1500);
nor U1981 (N_1981,N_1316,N_1383);
or U1982 (N_1982,N_1268,N_1552);
and U1983 (N_1983,N_1547,N_1512);
and U1984 (N_1984,N_1378,N_1619);
and U1985 (N_1985,N_1559,N_1672);
nand U1986 (N_1986,N_1351,N_1752);
nand U1987 (N_1987,N_1422,N_1367);
nor U1988 (N_1988,N_1749,N_1639);
nand U1989 (N_1989,N_1289,N_1521);
and U1990 (N_1990,N_1497,N_1245);
nor U1991 (N_1991,N_1435,N_1396);
xor U1992 (N_1992,N_1201,N_1507);
or U1993 (N_1993,N_1393,N_1235);
nand U1994 (N_1994,N_1527,N_1754);
nor U1995 (N_1995,N_1493,N_1420);
and U1996 (N_1996,N_1448,N_1444);
xor U1997 (N_1997,N_1605,N_1734);
or U1998 (N_1998,N_1203,N_1445);
xnor U1999 (N_1999,N_1593,N_1589);
or U2000 (N_2000,N_1243,N_1770);
xor U2001 (N_2001,N_1590,N_1488);
and U2002 (N_2002,N_1368,N_1776);
and U2003 (N_2003,N_1503,N_1333);
or U2004 (N_2004,N_1294,N_1611);
xnor U2005 (N_2005,N_1329,N_1354);
or U2006 (N_2006,N_1210,N_1617);
nand U2007 (N_2007,N_1522,N_1301);
nand U2008 (N_2008,N_1454,N_1600);
nand U2009 (N_2009,N_1269,N_1785);
and U2010 (N_2010,N_1654,N_1315);
xor U2011 (N_2011,N_1256,N_1326);
or U2012 (N_2012,N_1771,N_1657);
xor U2013 (N_2013,N_1608,N_1792);
nor U2014 (N_2014,N_1220,N_1429);
nor U2015 (N_2015,N_1455,N_1397);
or U2016 (N_2016,N_1664,N_1209);
or U2017 (N_2017,N_1217,N_1577);
xor U2018 (N_2018,N_1638,N_1630);
and U2019 (N_2019,N_1721,N_1275);
or U2020 (N_2020,N_1716,N_1371);
nand U2021 (N_2021,N_1214,N_1659);
xnor U2022 (N_2022,N_1744,N_1323);
nor U2023 (N_2023,N_1463,N_1682);
xnor U2024 (N_2024,N_1714,N_1765);
and U2025 (N_2025,N_1720,N_1384);
or U2026 (N_2026,N_1717,N_1424);
and U2027 (N_2027,N_1302,N_1382);
and U2028 (N_2028,N_1642,N_1458);
or U2029 (N_2029,N_1759,N_1254);
or U2030 (N_2030,N_1498,N_1586);
xor U2031 (N_2031,N_1787,N_1618);
nand U2032 (N_2032,N_1609,N_1239);
xnor U2033 (N_2033,N_1661,N_1748);
nor U2034 (N_2034,N_1637,N_1553);
xnor U2035 (N_2035,N_1283,N_1506);
and U2036 (N_2036,N_1399,N_1541);
or U2037 (N_2037,N_1620,N_1526);
or U2038 (N_2038,N_1433,N_1402);
nand U2039 (N_2039,N_1520,N_1360);
xnor U2040 (N_2040,N_1718,N_1536);
xor U2041 (N_2041,N_1280,N_1200);
xnor U2042 (N_2042,N_1238,N_1729);
nor U2043 (N_2043,N_1226,N_1276);
and U2044 (N_2044,N_1655,N_1575);
xnor U2045 (N_2045,N_1628,N_1363);
nand U2046 (N_2046,N_1438,N_1625);
nor U2047 (N_2047,N_1225,N_1598);
and U2048 (N_2048,N_1410,N_1472);
and U2049 (N_2049,N_1212,N_1392);
nor U2050 (N_2050,N_1735,N_1457);
or U2051 (N_2051,N_1358,N_1624);
or U2052 (N_2052,N_1423,N_1777);
and U2053 (N_2053,N_1636,N_1486);
nand U2054 (N_2054,N_1690,N_1649);
or U2055 (N_2055,N_1340,N_1799);
nor U2056 (N_2056,N_1688,N_1237);
nand U2057 (N_2057,N_1228,N_1216);
xnor U2058 (N_2058,N_1428,N_1788);
and U2059 (N_2059,N_1698,N_1757);
or U2060 (N_2060,N_1330,N_1614);
nor U2061 (N_2061,N_1469,N_1264);
nor U2062 (N_2062,N_1300,N_1634);
xnor U2063 (N_2063,N_1656,N_1421);
and U2064 (N_2064,N_1635,N_1395);
or U2065 (N_2065,N_1244,N_1282);
nor U2066 (N_2066,N_1314,N_1798);
and U2067 (N_2067,N_1562,N_1529);
nor U2068 (N_2068,N_1359,N_1538);
nor U2069 (N_2069,N_1366,N_1576);
nor U2070 (N_2070,N_1514,N_1691);
and U2071 (N_2071,N_1427,N_1715);
and U2072 (N_2072,N_1375,N_1413);
and U2073 (N_2073,N_1643,N_1328);
nand U2074 (N_2074,N_1745,N_1565);
xnor U2075 (N_2075,N_1408,N_1431);
nor U2076 (N_2076,N_1353,N_1790);
or U2077 (N_2077,N_1660,N_1537);
xor U2078 (N_2078,N_1299,N_1795);
nand U2079 (N_2079,N_1791,N_1540);
or U2080 (N_2080,N_1502,N_1558);
xnor U2081 (N_2081,N_1594,N_1305);
nor U2082 (N_2082,N_1712,N_1768);
and U2083 (N_2083,N_1505,N_1676);
or U2084 (N_2084,N_1361,N_1726);
nand U2085 (N_2085,N_1496,N_1599);
nor U2086 (N_2086,N_1725,N_1303);
or U2087 (N_2087,N_1604,N_1650);
xor U2088 (N_2088,N_1781,N_1539);
nor U2089 (N_2089,N_1297,N_1622);
nand U2090 (N_2090,N_1456,N_1554);
nor U2091 (N_2091,N_1476,N_1761);
xnor U2092 (N_2092,N_1587,N_1364);
and U2093 (N_2093,N_1404,N_1797);
nor U2094 (N_2094,N_1439,N_1523);
nor U2095 (N_2095,N_1723,N_1549);
nor U2096 (N_2096,N_1746,N_1449);
nor U2097 (N_2097,N_1246,N_1579);
nand U2098 (N_2098,N_1465,N_1259);
nand U2099 (N_2099,N_1266,N_1786);
xnor U2100 (N_2100,N_1601,N_1332);
or U2101 (N_2101,N_1470,N_1712);
nor U2102 (N_2102,N_1658,N_1201);
nor U2103 (N_2103,N_1652,N_1754);
xnor U2104 (N_2104,N_1369,N_1439);
xor U2105 (N_2105,N_1315,N_1518);
xor U2106 (N_2106,N_1521,N_1767);
and U2107 (N_2107,N_1768,N_1352);
nor U2108 (N_2108,N_1678,N_1247);
and U2109 (N_2109,N_1251,N_1310);
and U2110 (N_2110,N_1262,N_1212);
xor U2111 (N_2111,N_1602,N_1533);
and U2112 (N_2112,N_1246,N_1676);
or U2113 (N_2113,N_1350,N_1779);
nor U2114 (N_2114,N_1287,N_1660);
and U2115 (N_2115,N_1211,N_1363);
and U2116 (N_2116,N_1431,N_1288);
and U2117 (N_2117,N_1529,N_1519);
nor U2118 (N_2118,N_1699,N_1587);
nor U2119 (N_2119,N_1404,N_1556);
xor U2120 (N_2120,N_1771,N_1404);
and U2121 (N_2121,N_1348,N_1691);
and U2122 (N_2122,N_1350,N_1318);
nor U2123 (N_2123,N_1459,N_1625);
xnor U2124 (N_2124,N_1429,N_1371);
or U2125 (N_2125,N_1313,N_1295);
or U2126 (N_2126,N_1217,N_1239);
xnor U2127 (N_2127,N_1526,N_1668);
xnor U2128 (N_2128,N_1607,N_1640);
or U2129 (N_2129,N_1541,N_1606);
nor U2130 (N_2130,N_1585,N_1641);
nand U2131 (N_2131,N_1224,N_1719);
nor U2132 (N_2132,N_1714,N_1436);
and U2133 (N_2133,N_1772,N_1553);
and U2134 (N_2134,N_1325,N_1337);
nand U2135 (N_2135,N_1446,N_1693);
xnor U2136 (N_2136,N_1336,N_1248);
xnor U2137 (N_2137,N_1363,N_1751);
and U2138 (N_2138,N_1319,N_1211);
nand U2139 (N_2139,N_1454,N_1789);
nand U2140 (N_2140,N_1746,N_1344);
and U2141 (N_2141,N_1518,N_1618);
and U2142 (N_2142,N_1544,N_1337);
nand U2143 (N_2143,N_1460,N_1368);
or U2144 (N_2144,N_1492,N_1363);
or U2145 (N_2145,N_1367,N_1704);
xor U2146 (N_2146,N_1342,N_1579);
xnor U2147 (N_2147,N_1219,N_1474);
xnor U2148 (N_2148,N_1398,N_1430);
nand U2149 (N_2149,N_1798,N_1369);
xnor U2150 (N_2150,N_1520,N_1705);
nand U2151 (N_2151,N_1695,N_1215);
or U2152 (N_2152,N_1507,N_1291);
or U2153 (N_2153,N_1401,N_1226);
xnor U2154 (N_2154,N_1374,N_1592);
or U2155 (N_2155,N_1578,N_1434);
xnor U2156 (N_2156,N_1450,N_1651);
and U2157 (N_2157,N_1747,N_1427);
xnor U2158 (N_2158,N_1351,N_1781);
or U2159 (N_2159,N_1560,N_1266);
or U2160 (N_2160,N_1761,N_1401);
nor U2161 (N_2161,N_1523,N_1641);
or U2162 (N_2162,N_1279,N_1387);
xnor U2163 (N_2163,N_1534,N_1208);
and U2164 (N_2164,N_1565,N_1210);
nor U2165 (N_2165,N_1251,N_1212);
and U2166 (N_2166,N_1563,N_1219);
and U2167 (N_2167,N_1535,N_1515);
nor U2168 (N_2168,N_1448,N_1295);
xnor U2169 (N_2169,N_1263,N_1495);
or U2170 (N_2170,N_1679,N_1240);
xnor U2171 (N_2171,N_1419,N_1474);
or U2172 (N_2172,N_1394,N_1211);
and U2173 (N_2173,N_1489,N_1684);
or U2174 (N_2174,N_1770,N_1705);
xnor U2175 (N_2175,N_1764,N_1628);
and U2176 (N_2176,N_1598,N_1449);
and U2177 (N_2177,N_1754,N_1410);
nand U2178 (N_2178,N_1597,N_1344);
and U2179 (N_2179,N_1249,N_1429);
nor U2180 (N_2180,N_1767,N_1225);
xor U2181 (N_2181,N_1662,N_1253);
xnor U2182 (N_2182,N_1317,N_1551);
xnor U2183 (N_2183,N_1408,N_1436);
nand U2184 (N_2184,N_1565,N_1555);
and U2185 (N_2185,N_1578,N_1629);
xor U2186 (N_2186,N_1484,N_1446);
or U2187 (N_2187,N_1648,N_1674);
nor U2188 (N_2188,N_1476,N_1456);
and U2189 (N_2189,N_1291,N_1499);
and U2190 (N_2190,N_1389,N_1514);
nor U2191 (N_2191,N_1310,N_1274);
xor U2192 (N_2192,N_1602,N_1727);
nand U2193 (N_2193,N_1791,N_1298);
nor U2194 (N_2194,N_1626,N_1549);
xor U2195 (N_2195,N_1280,N_1299);
xnor U2196 (N_2196,N_1445,N_1609);
and U2197 (N_2197,N_1228,N_1471);
or U2198 (N_2198,N_1301,N_1514);
xor U2199 (N_2199,N_1774,N_1561);
xnor U2200 (N_2200,N_1630,N_1297);
nor U2201 (N_2201,N_1223,N_1601);
xnor U2202 (N_2202,N_1651,N_1407);
xnor U2203 (N_2203,N_1564,N_1736);
nand U2204 (N_2204,N_1562,N_1281);
xor U2205 (N_2205,N_1251,N_1688);
and U2206 (N_2206,N_1267,N_1676);
and U2207 (N_2207,N_1735,N_1553);
nand U2208 (N_2208,N_1774,N_1410);
and U2209 (N_2209,N_1422,N_1303);
xor U2210 (N_2210,N_1370,N_1358);
xor U2211 (N_2211,N_1445,N_1260);
or U2212 (N_2212,N_1530,N_1230);
and U2213 (N_2213,N_1760,N_1597);
or U2214 (N_2214,N_1539,N_1321);
nor U2215 (N_2215,N_1675,N_1699);
nand U2216 (N_2216,N_1295,N_1255);
and U2217 (N_2217,N_1298,N_1212);
nor U2218 (N_2218,N_1481,N_1666);
and U2219 (N_2219,N_1639,N_1755);
nand U2220 (N_2220,N_1718,N_1646);
or U2221 (N_2221,N_1732,N_1655);
xnor U2222 (N_2222,N_1294,N_1600);
nor U2223 (N_2223,N_1302,N_1694);
nor U2224 (N_2224,N_1606,N_1495);
nor U2225 (N_2225,N_1229,N_1434);
nand U2226 (N_2226,N_1306,N_1717);
and U2227 (N_2227,N_1453,N_1740);
or U2228 (N_2228,N_1533,N_1406);
xnor U2229 (N_2229,N_1525,N_1222);
nand U2230 (N_2230,N_1631,N_1360);
or U2231 (N_2231,N_1344,N_1427);
or U2232 (N_2232,N_1684,N_1349);
or U2233 (N_2233,N_1544,N_1776);
and U2234 (N_2234,N_1586,N_1529);
nor U2235 (N_2235,N_1230,N_1692);
nor U2236 (N_2236,N_1409,N_1254);
or U2237 (N_2237,N_1412,N_1762);
nand U2238 (N_2238,N_1428,N_1559);
nor U2239 (N_2239,N_1643,N_1293);
nor U2240 (N_2240,N_1471,N_1248);
nand U2241 (N_2241,N_1389,N_1607);
and U2242 (N_2242,N_1683,N_1414);
or U2243 (N_2243,N_1769,N_1348);
nand U2244 (N_2244,N_1200,N_1403);
or U2245 (N_2245,N_1370,N_1285);
nor U2246 (N_2246,N_1726,N_1374);
and U2247 (N_2247,N_1303,N_1765);
or U2248 (N_2248,N_1479,N_1526);
nor U2249 (N_2249,N_1322,N_1719);
and U2250 (N_2250,N_1296,N_1636);
xnor U2251 (N_2251,N_1588,N_1489);
nor U2252 (N_2252,N_1339,N_1745);
or U2253 (N_2253,N_1544,N_1233);
or U2254 (N_2254,N_1242,N_1707);
xor U2255 (N_2255,N_1773,N_1788);
or U2256 (N_2256,N_1616,N_1534);
xnor U2257 (N_2257,N_1287,N_1740);
xnor U2258 (N_2258,N_1727,N_1452);
xor U2259 (N_2259,N_1692,N_1470);
or U2260 (N_2260,N_1693,N_1645);
nor U2261 (N_2261,N_1427,N_1393);
nand U2262 (N_2262,N_1775,N_1629);
xnor U2263 (N_2263,N_1411,N_1563);
and U2264 (N_2264,N_1594,N_1519);
and U2265 (N_2265,N_1500,N_1532);
nor U2266 (N_2266,N_1471,N_1491);
nand U2267 (N_2267,N_1645,N_1636);
or U2268 (N_2268,N_1455,N_1370);
and U2269 (N_2269,N_1470,N_1321);
xor U2270 (N_2270,N_1595,N_1233);
or U2271 (N_2271,N_1705,N_1784);
or U2272 (N_2272,N_1573,N_1360);
xnor U2273 (N_2273,N_1590,N_1311);
nand U2274 (N_2274,N_1604,N_1386);
or U2275 (N_2275,N_1529,N_1398);
nor U2276 (N_2276,N_1664,N_1451);
nand U2277 (N_2277,N_1590,N_1293);
nor U2278 (N_2278,N_1475,N_1240);
or U2279 (N_2279,N_1235,N_1629);
xor U2280 (N_2280,N_1590,N_1443);
nand U2281 (N_2281,N_1599,N_1598);
nor U2282 (N_2282,N_1731,N_1502);
or U2283 (N_2283,N_1593,N_1319);
or U2284 (N_2284,N_1347,N_1472);
and U2285 (N_2285,N_1623,N_1723);
nor U2286 (N_2286,N_1256,N_1787);
xor U2287 (N_2287,N_1230,N_1404);
nor U2288 (N_2288,N_1391,N_1220);
xor U2289 (N_2289,N_1680,N_1258);
and U2290 (N_2290,N_1445,N_1254);
xnor U2291 (N_2291,N_1412,N_1245);
or U2292 (N_2292,N_1434,N_1765);
and U2293 (N_2293,N_1689,N_1726);
and U2294 (N_2294,N_1364,N_1794);
nand U2295 (N_2295,N_1584,N_1250);
nand U2296 (N_2296,N_1279,N_1218);
xor U2297 (N_2297,N_1462,N_1714);
or U2298 (N_2298,N_1419,N_1304);
nor U2299 (N_2299,N_1583,N_1236);
or U2300 (N_2300,N_1277,N_1552);
or U2301 (N_2301,N_1375,N_1607);
nor U2302 (N_2302,N_1691,N_1550);
or U2303 (N_2303,N_1653,N_1402);
nand U2304 (N_2304,N_1458,N_1607);
xnor U2305 (N_2305,N_1690,N_1203);
xor U2306 (N_2306,N_1305,N_1539);
or U2307 (N_2307,N_1443,N_1727);
or U2308 (N_2308,N_1705,N_1455);
or U2309 (N_2309,N_1369,N_1241);
or U2310 (N_2310,N_1586,N_1346);
xor U2311 (N_2311,N_1549,N_1322);
nand U2312 (N_2312,N_1295,N_1423);
nor U2313 (N_2313,N_1283,N_1640);
and U2314 (N_2314,N_1682,N_1518);
and U2315 (N_2315,N_1697,N_1470);
nand U2316 (N_2316,N_1663,N_1368);
or U2317 (N_2317,N_1205,N_1213);
and U2318 (N_2318,N_1549,N_1657);
nor U2319 (N_2319,N_1296,N_1734);
xnor U2320 (N_2320,N_1645,N_1245);
nor U2321 (N_2321,N_1241,N_1361);
or U2322 (N_2322,N_1519,N_1729);
and U2323 (N_2323,N_1687,N_1459);
nor U2324 (N_2324,N_1458,N_1368);
nand U2325 (N_2325,N_1289,N_1613);
and U2326 (N_2326,N_1774,N_1316);
nand U2327 (N_2327,N_1472,N_1601);
or U2328 (N_2328,N_1275,N_1636);
or U2329 (N_2329,N_1425,N_1213);
nand U2330 (N_2330,N_1728,N_1281);
nor U2331 (N_2331,N_1753,N_1638);
and U2332 (N_2332,N_1467,N_1335);
and U2333 (N_2333,N_1788,N_1423);
and U2334 (N_2334,N_1673,N_1600);
nand U2335 (N_2335,N_1692,N_1410);
and U2336 (N_2336,N_1306,N_1586);
or U2337 (N_2337,N_1312,N_1516);
xor U2338 (N_2338,N_1354,N_1705);
or U2339 (N_2339,N_1313,N_1234);
xor U2340 (N_2340,N_1710,N_1589);
xor U2341 (N_2341,N_1692,N_1634);
nor U2342 (N_2342,N_1768,N_1628);
nand U2343 (N_2343,N_1446,N_1513);
xor U2344 (N_2344,N_1276,N_1519);
nand U2345 (N_2345,N_1286,N_1445);
and U2346 (N_2346,N_1470,N_1772);
nor U2347 (N_2347,N_1332,N_1692);
and U2348 (N_2348,N_1451,N_1719);
and U2349 (N_2349,N_1672,N_1353);
or U2350 (N_2350,N_1692,N_1493);
or U2351 (N_2351,N_1516,N_1266);
xnor U2352 (N_2352,N_1392,N_1349);
nand U2353 (N_2353,N_1647,N_1657);
or U2354 (N_2354,N_1798,N_1609);
or U2355 (N_2355,N_1285,N_1735);
nor U2356 (N_2356,N_1236,N_1535);
or U2357 (N_2357,N_1649,N_1367);
or U2358 (N_2358,N_1556,N_1428);
or U2359 (N_2359,N_1645,N_1524);
and U2360 (N_2360,N_1798,N_1243);
or U2361 (N_2361,N_1589,N_1576);
nor U2362 (N_2362,N_1748,N_1603);
or U2363 (N_2363,N_1697,N_1211);
nor U2364 (N_2364,N_1618,N_1464);
nor U2365 (N_2365,N_1716,N_1504);
nand U2366 (N_2366,N_1460,N_1705);
nor U2367 (N_2367,N_1438,N_1751);
or U2368 (N_2368,N_1723,N_1379);
nor U2369 (N_2369,N_1490,N_1633);
xor U2370 (N_2370,N_1214,N_1666);
nor U2371 (N_2371,N_1404,N_1626);
xnor U2372 (N_2372,N_1599,N_1423);
xnor U2373 (N_2373,N_1608,N_1263);
nor U2374 (N_2374,N_1787,N_1497);
nor U2375 (N_2375,N_1593,N_1490);
nand U2376 (N_2376,N_1433,N_1791);
and U2377 (N_2377,N_1683,N_1344);
nand U2378 (N_2378,N_1592,N_1767);
and U2379 (N_2379,N_1609,N_1617);
or U2380 (N_2380,N_1281,N_1452);
or U2381 (N_2381,N_1682,N_1768);
nand U2382 (N_2382,N_1626,N_1449);
and U2383 (N_2383,N_1529,N_1492);
and U2384 (N_2384,N_1603,N_1394);
nand U2385 (N_2385,N_1717,N_1761);
nor U2386 (N_2386,N_1758,N_1309);
and U2387 (N_2387,N_1328,N_1314);
or U2388 (N_2388,N_1766,N_1695);
nand U2389 (N_2389,N_1628,N_1562);
xor U2390 (N_2390,N_1320,N_1327);
and U2391 (N_2391,N_1644,N_1260);
nand U2392 (N_2392,N_1381,N_1744);
nand U2393 (N_2393,N_1422,N_1773);
xor U2394 (N_2394,N_1266,N_1222);
nand U2395 (N_2395,N_1346,N_1456);
xor U2396 (N_2396,N_1476,N_1450);
and U2397 (N_2397,N_1734,N_1645);
or U2398 (N_2398,N_1498,N_1786);
xnor U2399 (N_2399,N_1633,N_1247);
nand U2400 (N_2400,N_2119,N_1980);
nand U2401 (N_2401,N_2391,N_2041);
xor U2402 (N_2402,N_2355,N_2397);
nor U2403 (N_2403,N_1918,N_1976);
nor U2404 (N_2404,N_1868,N_2225);
xnor U2405 (N_2405,N_2271,N_2223);
nor U2406 (N_2406,N_1981,N_2348);
nand U2407 (N_2407,N_1869,N_2115);
nand U2408 (N_2408,N_2054,N_2024);
xor U2409 (N_2409,N_1867,N_1933);
or U2410 (N_2410,N_2079,N_2237);
nand U2411 (N_2411,N_1952,N_2318);
xnor U2412 (N_2412,N_2309,N_1833);
or U2413 (N_2413,N_2205,N_2058);
and U2414 (N_2414,N_1916,N_2300);
nand U2415 (N_2415,N_2067,N_1817);
nand U2416 (N_2416,N_2181,N_1970);
xor U2417 (N_2417,N_2099,N_1820);
or U2418 (N_2418,N_2062,N_2144);
nand U2419 (N_2419,N_2023,N_2284);
nor U2420 (N_2420,N_2342,N_2037);
and U2421 (N_2421,N_2055,N_2220);
and U2422 (N_2422,N_1897,N_2343);
nor U2423 (N_2423,N_2094,N_1965);
nor U2424 (N_2424,N_1842,N_2340);
or U2425 (N_2425,N_2042,N_2235);
xnor U2426 (N_2426,N_2307,N_2159);
and U2427 (N_2427,N_1816,N_2392);
xnor U2428 (N_2428,N_2087,N_1846);
or U2429 (N_2429,N_2283,N_1852);
nand U2430 (N_2430,N_2113,N_2222);
nand U2431 (N_2431,N_2035,N_1861);
xnor U2432 (N_2432,N_2239,N_2091);
nand U2433 (N_2433,N_2388,N_1804);
nor U2434 (N_2434,N_2289,N_2395);
xor U2435 (N_2435,N_2232,N_1908);
nand U2436 (N_2436,N_1988,N_2206);
xnor U2437 (N_2437,N_2294,N_2290);
or U2438 (N_2438,N_2036,N_2350);
or U2439 (N_2439,N_2191,N_2049);
nand U2440 (N_2440,N_2163,N_1932);
nor U2441 (N_2441,N_1931,N_2269);
and U2442 (N_2442,N_1955,N_1996);
and U2443 (N_2443,N_2304,N_2168);
nor U2444 (N_2444,N_2227,N_2393);
or U2445 (N_2445,N_2177,N_2344);
and U2446 (N_2446,N_2129,N_1824);
or U2447 (N_2447,N_2215,N_1802);
and U2448 (N_2448,N_2174,N_2110);
nor U2449 (N_2449,N_2061,N_1902);
nor U2450 (N_2450,N_1888,N_1963);
nand U2451 (N_2451,N_2371,N_2127);
xnor U2452 (N_2452,N_1972,N_2019);
xor U2453 (N_2453,N_1989,N_2018);
xor U2454 (N_2454,N_1940,N_2199);
or U2455 (N_2455,N_1911,N_1862);
nor U2456 (N_2456,N_1878,N_2333);
and U2457 (N_2457,N_1815,N_1929);
nand U2458 (N_2458,N_2243,N_2245);
and U2459 (N_2459,N_1812,N_2224);
nand U2460 (N_2460,N_1857,N_1999);
nand U2461 (N_2461,N_1900,N_1984);
and U2462 (N_2462,N_1991,N_2085);
or U2463 (N_2463,N_2172,N_1847);
nor U2464 (N_2464,N_2069,N_2108);
xor U2465 (N_2465,N_2211,N_1905);
nand U2466 (N_2466,N_2261,N_2381);
or U2467 (N_2467,N_2286,N_2010);
and U2468 (N_2468,N_2250,N_2167);
nand U2469 (N_2469,N_2276,N_1865);
nand U2470 (N_2470,N_2007,N_1977);
or U2471 (N_2471,N_2095,N_2123);
and U2472 (N_2472,N_2154,N_1953);
or U2473 (N_2473,N_2260,N_1926);
and U2474 (N_2474,N_1913,N_2143);
or U2475 (N_2475,N_2238,N_2270);
and U2476 (N_2476,N_1990,N_2236);
and U2477 (N_2477,N_2396,N_1998);
nand U2478 (N_2478,N_1901,N_1956);
or U2479 (N_2479,N_2002,N_2106);
nor U2480 (N_2480,N_2394,N_1938);
nor U2481 (N_2481,N_2358,N_1946);
nor U2482 (N_2482,N_2248,N_2114);
nand U2483 (N_2483,N_1964,N_2162);
nand U2484 (N_2484,N_1805,N_2189);
nand U2485 (N_2485,N_2210,N_1822);
or U2486 (N_2486,N_1962,N_2370);
nand U2487 (N_2487,N_1966,N_2226);
nand U2488 (N_2488,N_2230,N_1982);
nand U2489 (N_2489,N_2029,N_2313);
nor U2490 (N_2490,N_2016,N_1967);
nand U2491 (N_2491,N_2126,N_2298);
nor U2492 (N_2492,N_1873,N_2130);
nand U2493 (N_2493,N_2098,N_2198);
or U2494 (N_2494,N_2213,N_1829);
nor U2495 (N_2495,N_2075,N_2074);
xor U2496 (N_2496,N_2195,N_2066);
xnor U2497 (N_2497,N_2332,N_1985);
or U2498 (N_2498,N_2012,N_2048);
xnor U2499 (N_2499,N_2202,N_1885);
and U2500 (N_2500,N_1922,N_1809);
or U2501 (N_2501,N_2273,N_1870);
and U2502 (N_2502,N_2229,N_1856);
and U2503 (N_2503,N_2104,N_2182);
and U2504 (N_2504,N_1854,N_1928);
or U2505 (N_2505,N_2386,N_2352);
nand U2506 (N_2506,N_1903,N_2112);
xnor U2507 (N_2507,N_2021,N_2297);
xor U2508 (N_2508,N_2073,N_1979);
and U2509 (N_2509,N_1887,N_2032);
nor U2510 (N_2510,N_2088,N_1904);
and U2511 (N_2511,N_2315,N_2004);
xor U2512 (N_2512,N_1808,N_2080);
or U2513 (N_2513,N_2389,N_2345);
xnor U2514 (N_2514,N_1961,N_1934);
or U2515 (N_2515,N_2338,N_2192);
or U2516 (N_2516,N_2096,N_2111);
or U2517 (N_2517,N_2179,N_1975);
or U2518 (N_2518,N_2217,N_2193);
and U2519 (N_2519,N_1923,N_1880);
nand U2520 (N_2520,N_1813,N_2285);
nand U2521 (N_2521,N_2322,N_2363);
and U2522 (N_2522,N_2169,N_1921);
nor U2523 (N_2523,N_1917,N_2158);
and U2524 (N_2524,N_2252,N_2266);
xnor U2525 (N_2525,N_2367,N_2103);
xnor U2526 (N_2526,N_1850,N_2118);
nand U2527 (N_2527,N_1872,N_2006);
or U2528 (N_2528,N_2296,N_1924);
and U2529 (N_2529,N_2038,N_2337);
nand U2530 (N_2530,N_2278,N_2040);
xnor U2531 (N_2531,N_1874,N_1910);
nor U2532 (N_2532,N_2317,N_2244);
and U2533 (N_2533,N_2207,N_1915);
or U2534 (N_2534,N_1927,N_2214);
or U2535 (N_2535,N_1866,N_2197);
nand U2536 (N_2536,N_2008,N_2184);
nand U2537 (N_2537,N_1837,N_1987);
nand U2538 (N_2538,N_1899,N_2282);
and U2539 (N_2539,N_2161,N_2334);
and U2540 (N_2540,N_2323,N_2131);
and U2541 (N_2541,N_1947,N_2288);
and U2542 (N_2542,N_2052,N_2132);
or U2543 (N_2543,N_1801,N_2009);
and U2544 (N_2544,N_2241,N_2152);
and U2545 (N_2545,N_1864,N_2145);
xnor U2546 (N_2546,N_2256,N_2136);
nand U2547 (N_2547,N_1830,N_2274);
and U2548 (N_2548,N_1906,N_1823);
xor U2549 (N_2549,N_2212,N_1859);
and U2550 (N_2550,N_2180,N_2135);
and U2551 (N_2551,N_2385,N_2233);
and U2552 (N_2552,N_2291,N_1858);
nor U2553 (N_2553,N_2240,N_1958);
xnor U2554 (N_2554,N_1919,N_2287);
xnor U2555 (N_2555,N_2321,N_2142);
and U2556 (N_2556,N_2133,N_2204);
or U2557 (N_2557,N_1914,N_2022);
and U2558 (N_2558,N_2308,N_2025);
xor U2559 (N_2559,N_1879,N_2272);
or U2560 (N_2560,N_1960,N_2076);
and U2561 (N_2561,N_2357,N_2314);
or U2562 (N_2562,N_1936,N_2183);
xnor U2563 (N_2563,N_1909,N_2335);
and U2564 (N_2564,N_1951,N_2319);
nor U2565 (N_2565,N_1945,N_2380);
nand U2566 (N_2566,N_2003,N_2302);
and U2567 (N_2567,N_2378,N_2125);
nor U2568 (N_2568,N_2147,N_2330);
or U2569 (N_2569,N_2387,N_2398);
or U2570 (N_2570,N_2100,N_2293);
xnor U2571 (N_2571,N_1810,N_2090);
or U2572 (N_2572,N_2082,N_2165);
xor U2573 (N_2573,N_1886,N_2228);
and U2574 (N_2574,N_2185,N_2219);
nand U2575 (N_2575,N_2155,N_2324);
nor U2576 (N_2576,N_2063,N_2031);
or U2577 (N_2577,N_1944,N_2186);
nand U2578 (N_2578,N_1968,N_2362);
nand U2579 (N_2579,N_2268,N_2005);
nand U2580 (N_2580,N_2316,N_2331);
nor U2581 (N_2581,N_2249,N_2234);
or U2582 (N_2582,N_2175,N_2336);
or U2583 (N_2583,N_1884,N_1844);
nand U2584 (N_2584,N_2017,N_2045);
xnor U2585 (N_2585,N_2320,N_1819);
nor U2586 (N_2586,N_2341,N_1821);
or U2587 (N_2587,N_1950,N_2188);
and U2588 (N_2588,N_1920,N_2015);
nor U2589 (N_2589,N_2001,N_2146);
or U2590 (N_2590,N_1832,N_1978);
nand U2591 (N_2591,N_2280,N_1840);
nand U2592 (N_2592,N_2301,N_2277);
nand U2593 (N_2593,N_2360,N_2097);
nand U2594 (N_2594,N_2384,N_2379);
xnor U2595 (N_2595,N_2328,N_2347);
xor U2596 (N_2596,N_1806,N_1892);
nand U2597 (N_2597,N_2390,N_2077);
nand U2598 (N_2598,N_1890,N_1834);
xnor U2599 (N_2599,N_2121,N_1848);
and U2600 (N_2600,N_2216,N_2372);
or U2601 (N_2601,N_2327,N_1893);
nor U2602 (N_2602,N_2072,N_2329);
and U2603 (N_2603,N_1853,N_2070);
xnor U2604 (N_2604,N_1925,N_2275);
and U2605 (N_2605,N_2050,N_1896);
and U2606 (N_2606,N_2039,N_2011);
or U2607 (N_2607,N_2306,N_1845);
xor U2608 (N_2608,N_2034,N_1891);
or U2609 (N_2609,N_1828,N_2056);
or U2610 (N_2610,N_1803,N_2218);
xor U2611 (N_2611,N_2014,N_2346);
nor U2612 (N_2612,N_2376,N_2164);
or U2613 (N_2613,N_1941,N_2292);
nor U2614 (N_2614,N_2148,N_1954);
nand U2615 (N_2615,N_2200,N_2265);
and U2616 (N_2616,N_1993,N_2255);
nand U2617 (N_2617,N_2065,N_1889);
nand U2618 (N_2618,N_2043,N_2305);
nand U2619 (N_2619,N_1969,N_2013);
nor U2620 (N_2620,N_1907,N_2083);
xor U2621 (N_2621,N_1992,N_1937);
nor U2622 (N_2622,N_2382,N_1836);
and U2623 (N_2623,N_2120,N_2101);
or U2624 (N_2624,N_2368,N_2377);
xnor U2625 (N_2625,N_2093,N_1943);
or U2626 (N_2626,N_2047,N_1959);
or U2627 (N_2627,N_1949,N_2089);
or U2628 (N_2628,N_2109,N_2369);
nor U2629 (N_2629,N_2176,N_1838);
nor U2630 (N_2630,N_2160,N_2326);
or U2631 (N_2631,N_2262,N_1826);
and U2632 (N_2632,N_1895,N_2353);
nand U2633 (N_2633,N_1841,N_1855);
nand U2634 (N_2634,N_2311,N_2020);
nor U2635 (N_2635,N_2151,N_2267);
xnor U2636 (N_2636,N_2122,N_2257);
xor U2637 (N_2637,N_2231,N_1882);
nand U2638 (N_2638,N_1811,N_2263);
and U2639 (N_2639,N_2383,N_2156);
or U2640 (N_2640,N_2196,N_1983);
nand U2641 (N_2641,N_1839,N_1912);
xor U2642 (N_2642,N_1994,N_2139);
and U2643 (N_2643,N_2351,N_2086);
xor U2644 (N_2644,N_2312,N_2359);
and U2645 (N_2645,N_2325,N_2399);
nor U2646 (N_2646,N_1863,N_2057);
xnor U2647 (N_2647,N_2201,N_2373);
xor U2648 (N_2648,N_2365,N_2246);
nand U2649 (N_2649,N_1827,N_2128);
nor U2650 (N_2650,N_2000,N_1800);
nand U2651 (N_2651,N_2242,N_2064);
nor U2652 (N_2652,N_2364,N_2279);
nand U2653 (N_2653,N_1898,N_1871);
and U2654 (N_2654,N_2060,N_2026);
nor U2655 (N_2655,N_2166,N_2157);
nand U2656 (N_2656,N_2051,N_2253);
nor U2657 (N_2657,N_2310,N_2354);
nand U2658 (N_2658,N_1849,N_2194);
xnor U2659 (N_2659,N_2059,N_1957);
and U2660 (N_2660,N_2366,N_1971);
or U2661 (N_2661,N_1948,N_2078);
nand U2662 (N_2662,N_2150,N_2361);
nor U2663 (N_2663,N_1939,N_2187);
nor U2664 (N_2664,N_1930,N_2190);
nor U2665 (N_2665,N_2171,N_2281);
nand U2666 (N_2666,N_2030,N_2138);
and U2667 (N_2667,N_1881,N_1876);
nand U2668 (N_2668,N_2251,N_1877);
xor U2669 (N_2669,N_1935,N_2081);
nand U2670 (N_2670,N_1814,N_1883);
or U2671 (N_2671,N_2084,N_2303);
or U2672 (N_2672,N_1843,N_2356);
and U2673 (N_2673,N_1894,N_1807);
or U2674 (N_2674,N_2105,N_2068);
nand U2675 (N_2675,N_2375,N_2254);
nor U2676 (N_2676,N_2027,N_2046);
or U2677 (N_2677,N_2140,N_2044);
xor U2678 (N_2678,N_1818,N_1974);
or U2679 (N_2679,N_2209,N_2173);
or U2680 (N_2680,N_2107,N_2117);
nor U2681 (N_2681,N_1973,N_2092);
or U2682 (N_2682,N_2299,N_1997);
nor U2683 (N_2683,N_2102,N_2033);
or U2684 (N_2684,N_1851,N_1860);
nand U2685 (N_2685,N_2374,N_1942);
nor U2686 (N_2686,N_2124,N_2141);
nor U2687 (N_2687,N_1986,N_2339);
or U2688 (N_2688,N_2208,N_2028);
and U2689 (N_2689,N_2295,N_2071);
and U2690 (N_2690,N_1825,N_2203);
nand U2691 (N_2691,N_2221,N_2153);
or U2692 (N_2692,N_2134,N_2170);
nor U2693 (N_2693,N_2053,N_2247);
xor U2694 (N_2694,N_1995,N_2349);
nand U2695 (N_2695,N_2137,N_2149);
nor U2696 (N_2696,N_1835,N_2258);
nand U2697 (N_2697,N_2116,N_1831);
or U2698 (N_2698,N_2259,N_2264);
or U2699 (N_2699,N_2178,N_1875);
and U2700 (N_2700,N_2121,N_1996);
or U2701 (N_2701,N_2308,N_2109);
nor U2702 (N_2702,N_2009,N_2331);
and U2703 (N_2703,N_2206,N_2074);
nand U2704 (N_2704,N_1982,N_2292);
nand U2705 (N_2705,N_1807,N_2200);
nor U2706 (N_2706,N_1968,N_2172);
and U2707 (N_2707,N_2066,N_1890);
nor U2708 (N_2708,N_2346,N_2138);
and U2709 (N_2709,N_1913,N_2053);
nand U2710 (N_2710,N_2178,N_2265);
and U2711 (N_2711,N_2148,N_2001);
nor U2712 (N_2712,N_2114,N_2023);
or U2713 (N_2713,N_1804,N_2206);
nand U2714 (N_2714,N_2259,N_1874);
nor U2715 (N_2715,N_1992,N_1950);
and U2716 (N_2716,N_2206,N_2063);
nand U2717 (N_2717,N_1804,N_1815);
nand U2718 (N_2718,N_2089,N_2356);
nand U2719 (N_2719,N_2246,N_2216);
nor U2720 (N_2720,N_2160,N_2081);
nor U2721 (N_2721,N_2213,N_2313);
nor U2722 (N_2722,N_1843,N_2003);
nand U2723 (N_2723,N_2102,N_2332);
or U2724 (N_2724,N_2253,N_2110);
and U2725 (N_2725,N_2249,N_2354);
or U2726 (N_2726,N_2323,N_2012);
xor U2727 (N_2727,N_2027,N_2116);
or U2728 (N_2728,N_2324,N_2379);
xor U2729 (N_2729,N_2091,N_2013);
nand U2730 (N_2730,N_2392,N_2017);
and U2731 (N_2731,N_1806,N_2139);
and U2732 (N_2732,N_2081,N_2032);
nor U2733 (N_2733,N_2060,N_1899);
nor U2734 (N_2734,N_1838,N_2310);
or U2735 (N_2735,N_2040,N_2048);
and U2736 (N_2736,N_1923,N_2080);
xnor U2737 (N_2737,N_1935,N_1946);
xor U2738 (N_2738,N_1846,N_1979);
and U2739 (N_2739,N_1823,N_2173);
nand U2740 (N_2740,N_1945,N_2361);
xor U2741 (N_2741,N_1814,N_1911);
or U2742 (N_2742,N_2026,N_2086);
nor U2743 (N_2743,N_1868,N_2350);
nor U2744 (N_2744,N_1974,N_2008);
nand U2745 (N_2745,N_2154,N_1959);
xnor U2746 (N_2746,N_2290,N_1906);
nand U2747 (N_2747,N_2331,N_1969);
nand U2748 (N_2748,N_1850,N_2177);
xor U2749 (N_2749,N_2189,N_1826);
xor U2750 (N_2750,N_2088,N_1826);
and U2751 (N_2751,N_1888,N_2284);
nor U2752 (N_2752,N_2135,N_2290);
nand U2753 (N_2753,N_2387,N_2339);
xnor U2754 (N_2754,N_1970,N_1887);
and U2755 (N_2755,N_2262,N_2344);
nor U2756 (N_2756,N_1971,N_1874);
or U2757 (N_2757,N_1951,N_2348);
or U2758 (N_2758,N_2011,N_1809);
and U2759 (N_2759,N_2217,N_1848);
and U2760 (N_2760,N_1943,N_2199);
xnor U2761 (N_2761,N_2254,N_2336);
nand U2762 (N_2762,N_1971,N_2086);
and U2763 (N_2763,N_1898,N_2371);
and U2764 (N_2764,N_1909,N_2097);
xor U2765 (N_2765,N_2273,N_2009);
xnor U2766 (N_2766,N_2267,N_2075);
nor U2767 (N_2767,N_2225,N_2145);
and U2768 (N_2768,N_2323,N_2080);
or U2769 (N_2769,N_2347,N_1851);
nor U2770 (N_2770,N_2373,N_2005);
nand U2771 (N_2771,N_2263,N_2090);
or U2772 (N_2772,N_1856,N_1879);
and U2773 (N_2773,N_1889,N_2267);
nand U2774 (N_2774,N_1874,N_2363);
nor U2775 (N_2775,N_2385,N_1831);
nand U2776 (N_2776,N_1984,N_2014);
or U2777 (N_2777,N_1979,N_1917);
nand U2778 (N_2778,N_2317,N_2376);
nand U2779 (N_2779,N_1875,N_2222);
xor U2780 (N_2780,N_2081,N_2370);
xnor U2781 (N_2781,N_2002,N_2316);
nand U2782 (N_2782,N_2221,N_2217);
or U2783 (N_2783,N_1819,N_1947);
and U2784 (N_2784,N_2375,N_2237);
nand U2785 (N_2785,N_1880,N_2344);
or U2786 (N_2786,N_1970,N_1899);
xnor U2787 (N_2787,N_2154,N_2061);
and U2788 (N_2788,N_2063,N_2114);
nand U2789 (N_2789,N_2148,N_2223);
or U2790 (N_2790,N_2112,N_2173);
or U2791 (N_2791,N_2189,N_1996);
nand U2792 (N_2792,N_2275,N_1816);
xor U2793 (N_2793,N_2305,N_1909);
and U2794 (N_2794,N_2245,N_2099);
xnor U2795 (N_2795,N_1850,N_2114);
nor U2796 (N_2796,N_2234,N_2012);
or U2797 (N_2797,N_1982,N_2032);
nor U2798 (N_2798,N_1893,N_2023);
and U2799 (N_2799,N_2260,N_2199);
xor U2800 (N_2800,N_2259,N_2101);
or U2801 (N_2801,N_2222,N_2109);
or U2802 (N_2802,N_1926,N_2377);
xnor U2803 (N_2803,N_2174,N_2226);
nand U2804 (N_2804,N_2067,N_1858);
and U2805 (N_2805,N_2276,N_2252);
xor U2806 (N_2806,N_1926,N_2045);
nor U2807 (N_2807,N_1977,N_2367);
xor U2808 (N_2808,N_2272,N_1850);
nor U2809 (N_2809,N_1903,N_2306);
xor U2810 (N_2810,N_2234,N_2280);
and U2811 (N_2811,N_1919,N_2205);
or U2812 (N_2812,N_2226,N_2294);
or U2813 (N_2813,N_1970,N_1815);
xor U2814 (N_2814,N_1878,N_2062);
or U2815 (N_2815,N_2289,N_2092);
xor U2816 (N_2816,N_1994,N_1852);
xor U2817 (N_2817,N_2078,N_2342);
xnor U2818 (N_2818,N_2012,N_1800);
xor U2819 (N_2819,N_1948,N_1838);
xor U2820 (N_2820,N_2191,N_2137);
or U2821 (N_2821,N_1909,N_2373);
xor U2822 (N_2822,N_2236,N_2367);
nor U2823 (N_2823,N_1995,N_2111);
or U2824 (N_2824,N_2210,N_2270);
or U2825 (N_2825,N_2386,N_2164);
nor U2826 (N_2826,N_1929,N_2331);
xnor U2827 (N_2827,N_1838,N_2104);
or U2828 (N_2828,N_2043,N_1986);
nor U2829 (N_2829,N_2026,N_2291);
nor U2830 (N_2830,N_2290,N_2065);
nor U2831 (N_2831,N_1873,N_2254);
xnor U2832 (N_2832,N_2078,N_2244);
nor U2833 (N_2833,N_1958,N_2383);
or U2834 (N_2834,N_1850,N_1863);
and U2835 (N_2835,N_2288,N_1996);
and U2836 (N_2836,N_2316,N_2311);
xor U2837 (N_2837,N_2319,N_1900);
and U2838 (N_2838,N_1998,N_2170);
xor U2839 (N_2839,N_1878,N_2262);
nand U2840 (N_2840,N_1925,N_2170);
xor U2841 (N_2841,N_2339,N_2185);
or U2842 (N_2842,N_1820,N_2176);
nand U2843 (N_2843,N_1896,N_2151);
xor U2844 (N_2844,N_2152,N_2169);
nand U2845 (N_2845,N_1987,N_1978);
and U2846 (N_2846,N_2134,N_1850);
or U2847 (N_2847,N_1868,N_2064);
and U2848 (N_2848,N_2191,N_2163);
nor U2849 (N_2849,N_2005,N_1819);
xor U2850 (N_2850,N_2345,N_2000);
or U2851 (N_2851,N_2195,N_1921);
nand U2852 (N_2852,N_2043,N_2267);
and U2853 (N_2853,N_2100,N_2294);
or U2854 (N_2854,N_1943,N_2372);
xnor U2855 (N_2855,N_2202,N_2333);
nor U2856 (N_2856,N_1919,N_2273);
and U2857 (N_2857,N_1990,N_2121);
nor U2858 (N_2858,N_2176,N_2018);
xnor U2859 (N_2859,N_2236,N_1858);
nand U2860 (N_2860,N_2364,N_2192);
nor U2861 (N_2861,N_2032,N_1990);
xnor U2862 (N_2862,N_2375,N_1983);
nor U2863 (N_2863,N_2323,N_1853);
or U2864 (N_2864,N_1988,N_2136);
xor U2865 (N_2865,N_2206,N_1817);
or U2866 (N_2866,N_2313,N_2109);
xnor U2867 (N_2867,N_2230,N_1803);
nand U2868 (N_2868,N_2164,N_2372);
and U2869 (N_2869,N_2220,N_1817);
nand U2870 (N_2870,N_2190,N_2192);
and U2871 (N_2871,N_2145,N_2215);
or U2872 (N_2872,N_1920,N_2156);
xnor U2873 (N_2873,N_1857,N_2133);
and U2874 (N_2874,N_2053,N_2243);
nand U2875 (N_2875,N_1832,N_2283);
nand U2876 (N_2876,N_2259,N_1867);
nor U2877 (N_2877,N_2331,N_2195);
or U2878 (N_2878,N_1889,N_2163);
nand U2879 (N_2879,N_1966,N_1997);
xor U2880 (N_2880,N_1872,N_2113);
and U2881 (N_2881,N_2173,N_2087);
xnor U2882 (N_2882,N_1940,N_2015);
xnor U2883 (N_2883,N_2235,N_2212);
xor U2884 (N_2884,N_2230,N_2379);
or U2885 (N_2885,N_2282,N_2370);
or U2886 (N_2886,N_1883,N_1831);
xnor U2887 (N_2887,N_2014,N_2301);
nor U2888 (N_2888,N_2076,N_2087);
and U2889 (N_2889,N_1913,N_2115);
and U2890 (N_2890,N_2174,N_1869);
nand U2891 (N_2891,N_1850,N_1807);
and U2892 (N_2892,N_2298,N_1972);
nor U2893 (N_2893,N_2283,N_1827);
and U2894 (N_2894,N_2335,N_2112);
or U2895 (N_2895,N_1863,N_2079);
or U2896 (N_2896,N_1872,N_2356);
or U2897 (N_2897,N_2216,N_2393);
xnor U2898 (N_2898,N_2263,N_1958);
nand U2899 (N_2899,N_2337,N_1954);
or U2900 (N_2900,N_1846,N_1827);
and U2901 (N_2901,N_2150,N_1841);
or U2902 (N_2902,N_2258,N_2344);
nand U2903 (N_2903,N_1842,N_2302);
or U2904 (N_2904,N_1841,N_2263);
nor U2905 (N_2905,N_2117,N_2271);
nor U2906 (N_2906,N_2354,N_2243);
and U2907 (N_2907,N_2220,N_1849);
nor U2908 (N_2908,N_2227,N_1920);
or U2909 (N_2909,N_1978,N_2101);
or U2910 (N_2910,N_2309,N_2307);
or U2911 (N_2911,N_1922,N_2093);
nand U2912 (N_2912,N_2090,N_1864);
xor U2913 (N_2913,N_2145,N_1948);
nor U2914 (N_2914,N_2013,N_2140);
and U2915 (N_2915,N_1929,N_1956);
xnor U2916 (N_2916,N_1859,N_2177);
nor U2917 (N_2917,N_2008,N_2090);
or U2918 (N_2918,N_1858,N_2351);
and U2919 (N_2919,N_1842,N_2059);
nand U2920 (N_2920,N_2344,N_2066);
or U2921 (N_2921,N_2002,N_2184);
xor U2922 (N_2922,N_2223,N_2345);
and U2923 (N_2923,N_2222,N_2117);
and U2924 (N_2924,N_2174,N_2044);
nand U2925 (N_2925,N_2291,N_2199);
or U2926 (N_2926,N_2358,N_2154);
xor U2927 (N_2927,N_1852,N_2061);
nand U2928 (N_2928,N_2382,N_2098);
and U2929 (N_2929,N_2022,N_1941);
nand U2930 (N_2930,N_2193,N_1874);
nor U2931 (N_2931,N_2042,N_1898);
xor U2932 (N_2932,N_2039,N_1956);
xor U2933 (N_2933,N_2345,N_1901);
nand U2934 (N_2934,N_2227,N_1946);
nand U2935 (N_2935,N_2157,N_2036);
and U2936 (N_2936,N_1918,N_1926);
nand U2937 (N_2937,N_2162,N_1967);
or U2938 (N_2938,N_2114,N_1978);
or U2939 (N_2939,N_2232,N_2219);
nor U2940 (N_2940,N_2378,N_1827);
and U2941 (N_2941,N_2177,N_2377);
nor U2942 (N_2942,N_2132,N_2242);
nor U2943 (N_2943,N_2068,N_2032);
or U2944 (N_2944,N_2345,N_2246);
xor U2945 (N_2945,N_2120,N_2018);
nor U2946 (N_2946,N_1902,N_2384);
or U2947 (N_2947,N_2214,N_1923);
xor U2948 (N_2948,N_1804,N_2017);
nor U2949 (N_2949,N_1961,N_2245);
nor U2950 (N_2950,N_2105,N_2000);
xor U2951 (N_2951,N_2107,N_2277);
nand U2952 (N_2952,N_2076,N_2394);
or U2953 (N_2953,N_1915,N_2223);
and U2954 (N_2954,N_1985,N_1819);
and U2955 (N_2955,N_1830,N_2168);
or U2956 (N_2956,N_2210,N_2212);
nand U2957 (N_2957,N_2158,N_1925);
and U2958 (N_2958,N_2358,N_2290);
nor U2959 (N_2959,N_2018,N_2285);
or U2960 (N_2960,N_2107,N_1922);
nor U2961 (N_2961,N_2301,N_2229);
nand U2962 (N_2962,N_2189,N_2135);
or U2963 (N_2963,N_1948,N_2022);
nor U2964 (N_2964,N_2106,N_2056);
and U2965 (N_2965,N_2069,N_1988);
xnor U2966 (N_2966,N_2231,N_2352);
xnor U2967 (N_2967,N_2070,N_2162);
nand U2968 (N_2968,N_2389,N_2102);
xnor U2969 (N_2969,N_1958,N_2026);
xor U2970 (N_2970,N_2374,N_2263);
and U2971 (N_2971,N_2166,N_2151);
or U2972 (N_2972,N_1843,N_2342);
and U2973 (N_2973,N_2044,N_1959);
nor U2974 (N_2974,N_2134,N_1958);
nand U2975 (N_2975,N_1933,N_1843);
xnor U2976 (N_2976,N_2324,N_2253);
nor U2977 (N_2977,N_2048,N_2238);
or U2978 (N_2978,N_2080,N_1872);
nand U2979 (N_2979,N_2307,N_2230);
nor U2980 (N_2980,N_1909,N_2164);
nand U2981 (N_2981,N_2350,N_2207);
xor U2982 (N_2982,N_2050,N_2195);
nor U2983 (N_2983,N_2067,N_1844);
or U2984 (N_2984,N_2076,N_2071);
and U2985 (N_2985,N_1831,N_2133);
xor U2986 (N_2986,N_2212,N_2010);
nand U2987 (N_2987,N_1893,N_2132);
nand U2988 (N_2988,N_2364,N_2328);
nor U2989 (N_2989,N_2043,N_2364);
nand U2990 (N_2990,N_1968,N_2278);
nor U2991 (N_2991,N_2175,N_2065);
and U2992 (N_2992,N_1833,N_1926);
or U2993 (N_2993,N_2033,N_1923);
xor U2994 (N_2994,N_2093,N_1927);
nor U2995 (N_2995,N_1832,N_2178);
nor U2996 (N_2996,N_2032,N_2106);
nand U2997 (N_2997,N_1926,N_2012);
xnor U2998 (N_2998,N_2004,N_1941);
nor U2999 (N_2999,N_2149,N_1885);
xor UO_0 (O_0,N_2620,N_2722);
or UO_1 (O_1,N_2436,N_2460);
or UO_2 (O_2,N_2601,N_2516);
or UO_3 (O_3,N_2437,N_2865);
xor UO_4 (O_4,N_2679,N_2962);
or UO_5 (O_5,N_2806,N_2606);
and UO_6 (O_6,N_2415,N_2653);
or UO_7 (O_7,N_2639,N_2476);
and UO_8 (O_8,N_2830,N_2974);
xnor UO_9 (O_9,N_2984,N_2633);
and UO_10 (O_10,N_2877,N_2645);
nand UO_11 (O_11,N_2610,N_2863);
or UO_12 (O_12,N_2473,N_2424);
and UO_13 (O_13,N_2650,N_2920);
xnor UO_14 (O_14,N_2922,N_2836);
xor UO_15 (O_15,N_2578,N_2738);
nor UO_16 (O_16,N_2958,N_2894);
nand UO_17 (O_17,N_2717,N_2915);
xnor UO_18 (O_18,N_2659,N_2888);
and UO_19 (O_19,N_2911,N_2528);
and UO_20 (O_20,N_2994,N_2826);
nor UO_21 (O_21,N_2847,N_2440);
nand UO_22 (O_22,N_2411,N_2693);
or UO_23 (O_23,N_2593,N_2490);
nor UO_24 (O_24,N_2913,N_2672);
nand UO_25 (O_25,N_2742,N_2663);
and UO_26 (O_26,N_2542,N_2741);
and UO_27 (O_27,N_2932,N_2782);
nor UO_28 (O_28,N_2892,N_2952);
and UO_29 (O_29,N_2852,N_2868);
xor UO_30 (O_30,N_2749,N_2454);
nand UO_31 (O_31,N_2690,N_2858);
or UO_32 (O_32,N_2548,N_2446);
nor UO_33 (O_33,N_2763,N_2621);
and UO_34 (O_34,N_2678,N_2756);
nor UO_35 (O_35,N_2552,N_2919);
xor UO_36 (O_36,N_2687,N_2872);
nand UO_37 (O_37,N_2546,N_2670);
nor UO_38 (O_38,N_2455,N_2889);
nor UO_39 (O_39,N_2870,N_2481);
nor UO_40 (O_40,N_2615,N_2416);
nand UO_41 (O_41,N_2864,N_2898);
nand UO_42 (O_42,N_2776,N_2676);
and UO_43 (O_43,N_2406,N_2684);
and UO_44 (O_44,N_2703,N_2423);
and UO_45 (O_45,N_2926,N_2708);
and UO_46 (O_46,N_2401,N_2602);
or UO_47 (O_47,N_2982,N_2853);
nand UO_48 (O_48,N_2517,N_2686);
or UO_49 (O_49,N_2873,N_2859);
nor UO_50 (O_50,N_2583,N_2652);
xor UO_51 (O_51,N_2488,N_2584);
xnor UO_52 (O_52,N_2587,N_2456);
or UO_53 (O_53,N_2808,N_2486);
nand UO_54 (O_54,N_2443,N_2472);
and UO_55 (O_55,N_2657,N_2532);
or UO_56 (O_56,N_2519,N_2407);
or UO_57 (O_57,N_2524,N_2483);
nor UO_58 (O_58,N_2910,N_2726);
xor UO_59 (O_59,N_2414,N_2500);
xnor UO_60 (O_60,N_2625,N_2945);
nor UO_61 (O_61,N_2995,N_2970);
nor UO_62 (O_62,N_2997,N_2783);
nand UO_63 (O_63,N_2513,N_2885);
xor UO_64 (O_64,N_2908,N_2711);
xor UO_65 (O_65,N_2560,N_2784);
or UO_66 (O_66,N_2824,N_2507);
and UO_67 (O_67,N_2939,N_2940);
or UO_68 (O_68,N_2555,N_2655);
xor UO_69 (O_69,N_2767,N_2421);
or UO_70 (O_70,N_2732,N_2575);
xor UO_71 (O_71,N_2981,N_2953);
nor UO_72 (O_72,N_2880,N_2760);
nand UO_73 (O_73,N_2505,N_2478);
and UO_74 (O_74,N_2835,N_2701);
or UO_75 (O_75,N_2903,N_2842);
and UO_76 (O_76,N_2772,N_2420);
xor UO_77 (O_77,N_2720,N_2599);
or UO_78 (O_78,N_2462,N_2484);
or UO_79 (O_79,N_2739,N_2860);
or UO_80 (O_80,N_2967,N_2807);
and UO_81 (O_81,N_2805,N_2809);
nor UO_82 (O_82,N_2937,N_2656);
nand UO_83 (O_83,N_2669,N_2603);
and UO_84 (O_84,N_2475,N_2530);
and UO_85 (O_85,N_2408,N_2631);
xnor UO_86 (O_86,N_2534,N_2660);
xnor UO_87 (O_87,N_2719,N_2707);
or UO_88 (O_88,N_2907,N_2536);
xor UO_89 (O_89,N_2512,N_2777);
or UO_90 (O_90,N_2674,N_2518);
or UO_91 (O_91,N_2886,N_2727);
nor UO_92 (O_92,N_2794,N_2677);
and UO_93 (O_93,N_2554,N_2773);
or UO_94 (O_94,N_2551,N_2789);
and UO_95 (O_95,N_2923,N_2626);
and UO_96 (O_96,N_2980,N_2457);
nor UO_97 (O_97,N_2831,N_2662);
nor UO_98 (O_98,N_2430,N_2881);
and UO_99 (O_99,N_2856,N_2649);
or UO_100 (O_100,N_2562,N_2931);
xor UO_101 (O_101,N_2751,N_2503);
and UO_102 (O_102,N_2628,N_2692);
nand UO_103 (O_103,N_2410,N_2422);
or UO_104 (O_104,N_2441,N_2569);
and UO_105 (O_105,N_2497,N_2594);
or UO_106 (O_106,N_2567,N_2957);
or UO_107 (O_107,N_2468,N_2874);
nor UO_108 (O_108,N_2774,N_2718);
nand UO_109 (O_109,N_2523,N_2447);
and UO_110 (O_110,N_2985,N_2816);
nor UO_111 (O_111,N_2986,N_2458);
and UO_112 (O_112,N_2916,N_2812);
and UO_113 (O_113,N_2613,N_2696);
nor UO_114 (O_114,N_2418,N_2752);
xnor UO_115 (O_115,N_2938,N_2492);
xor UO_116 (O_116,N_2733,N_2721);
nand UO_117 (O_117,N_2566,N_2788);
nand UO_118 (O_118,N_2884,N_2522);
nand UO_119 (O_119,N_2704,N_2493);
nor UO_120 (O_120,N_2851,N_2553);
nand UO_121 (O_121,N_2409,N_2637);
and UO_122 (O_122,N_2956,N_2453);
nand UO_123 (O_123,N_2841,N_2582);
nor UO_124 (O_124,N_2768,N_2736);
nor UO_125 (O_125,N_2491,N_2833);
or UO_126 (O_126,N_2878,N_2658);
nand UO_127 (O_127,N_2747,N_2438);
nor UO_128 (O_128,N_2502,N_2654);
xor UO_129 (O_129,N_2465,N_2682);
nor UO_130 (O_130,N_2861,N_2999);
nand UO_131 (O_131,N_2461,N_2731);
nor UO_132 (O_132,N_2564,N_2758);
or UO_133 (O_133,N_2675,N_2963);
nand UO_134 (O_134,N_2769,N_2558);
nor UO_135 (O_135,N_2821,N_2787);
nand UO_136 (O_136,N_2790,N_2728);
nor UO_137 (O_137,N_2681,N_2539);
nand UO_138 (O_138,N_2799,N_2664);
nor UO_139 (O_139,N_2622,N_2757);
nor UO_140 (O_140,N_2434,N_2730);
or UO_141 (O_141,N_2604,N_2734);
nor UO_142 (O_142,N_2705,N_2725);
or UO_143 (O_143,N_2404,N_2469);
xnor UO_144 (O_144,N_2815,N_2494);
nor UO_145 (O_145,N_2972,N_2452);
and UO_146 (O_146,N_2825,N_2811);
nand UO_147 (O_147,N_2869,N_2629);
and UO_148 (O_148,N_2557,N_2897);
nor UO_149 (O_149,N_2533,N_2618);
nor UO_150 (O_150,N_2527,N_2998);
nor UO_151 (O_151,N_2688,N_2561);
and UO_152 (O_152,N_2433,N_2771);
or UO_153 (O_153,N_2803,N_2798);
nand UO_154 (O_154,N_2425,N_2685);
or UO_155 (O_155,N_2862,N_2918);
nor UO_156 (O_156,N_2796,N_2933);
and UO_157 (O_157,N_2431,N_2780);
xnor UO_158 (O_158,N_2598,N_2909);
and UO_159 (O_159,N_2944,N_2680);
and UO_160 (O_160,N_2827,N_2753);
nand UO_161 (O_161,N_2540,N_2586);
nand UO_162 (O_162,N_2417,N_2463);
and UO_163 (O_163,N_2448,N_2973);
or UO_164 (O_164,N_2579,N_2596);
and UO_165 (O_165,N_2700,N_2979);
xnor UO_166 (O_166,N_2935,N_2451);
nor UO_167 (O_167,N_2668,N_2729);
nand UO_168 (O_168,N_2744,N_2781);
nand UO_169 (O_169,N_2951,N_2934);
and UO_170 (O_170,N_2823,N_2444);
nor UO_171 (O_171,N_2499,N_2574);
nor UO_172 (O_172,N_2890,N_2403);
nand UO_173 (O_173,N_2627,N_2432);
nand UO_174 (O_174,N_2996,N_2459);
and UO_175 (O_175,N_2571,N_2900);
or UO_176 (O_176,N_2445,N_2636);
or UO_177 (O_177,N_2541,N_2959);
or UO_178 (O_178,N_2971,N_2930);
and UO_179 (O_179,N_2644,N_2565);
or UO_180 (O_180,N_2817,N_2891);
nor UO_181 (O_181,N_2577,N_2611);
or UO_182 (O_182,N_2419,N_2702);
or UO_183 (O_183,N_2845,N_2683);
nand UO_184 (O_184,N_2792,N_2485);
nor UO_185 (O_185,N_2810,N_2665);
nand UO_186 (O_186,N_2914,N_2715);
nand UO_187 (O_187,N_2879,N_2474);
and UO_188 (O_188,N_2800,N_2901);
or UO_189 (O_189,N_2521,N_2829);
xor UO_190 (O_190,N_2837,N_2820);
nand UO_191 (O_191,N_2543,N_2537);
xor UO_192 (O_192,N_2866,N_2902);
xor UO_193 (O_193,N_2617,N_2412);
or UO_194 (O_194,N_2716,N_2887);
nand UO_195 (O_195,N_2813,N_2843);
xnor UO_196 (O_196,N_2960,N_2619);
nor UO_197 (O_197,N_2975,N_2871);
xnor UO_198 (O_198,N_2651,N_2466);
nor UO_199 (O_199,N_2941,N_2762);
or UO_200 (O_200,N_2710,N_2882);
and UO_201 (O_201,N_2426,N_2802);
and UO_202 (O_202,N_2612,N_2470);
or UO_203 (O_203,N_2589,N_2641);
nand UO_204 (O_204,N_2899,N_2508);
or UO_205 (O_205,N_2495,N_2597);
and UO_206 (O_206,N_2814,N_2917);
xnor UO_207 (O_207,N_2405,N_2605);
nor UO_208 (O_208,N_2969,N_2576);
xnor UO_209 (O_209,N_2713,N_2992);
and UO_210 (O_210,N_2989,N_2514);
and UO_211 (O_211,N_2666,N_2695);
nor UO_212 (O_212,N_2976,N_2766);
or UO_213 (O_213,N_2801,N_2489);
and UO_214 (O_214,N_2950,N_2895);
nand UO_215 (O_215,N_2667,N_2550);
nand UO_216 (O_216,N_2797,N_2966);
and UO_217 (O_217,N_2954,N_2531);
and UO_218 (O_218,N_2600,N_2661);
nand UO_219 (O_219,N_2961,N_2990);
nand UO_220 (O_220,N_2750,N_2487);
xor UO_221 (O_221,N_2924,N_2712);
nor UO_222 (O_222,N_2544,N_2526);
or UO_223 (O_223,N_2623,N_2689);
nor UO_224 (O_224,N_2977,N_2697);
xor UO_225 (O_225,N_2640,N_2844);
and UO_226 (O_226,N_2785,N_2743);
or UO_227 (O_227,N_2987,N_2883);
or UO_228 (O_228,N_2840,N_2624);
or UO_229 (O_229,N_2754,N_2525);
xnor UO_230 (O_230,N_2607,N_2504);
xnor UO_231 (O_231,N_2714,N_2838);
and UO_232 (O_232,N_2988,N_2983);
and UO_233 (O_233,N_2706,N_2949);
nand UO_234 (O_234,N_2450,N_2634);
or UO_235 (O_235,N_2616,N_2556);
nand UO_236 (O_236,N_2647,N_2608);
nand UO_237 (O_237,N_2896,N_2875);
xnor UO_238 (O_238,N_2671,N_2828);
or UO_239 (O_239,N_2804,N_2955);
xor UO_240 (O_240,N_2740,N_2635);
or UO_241 (O_241,N_2609,N_2529);
xnor UO_242 (O_242,N_2942,N_2427);
nand UO_243 (O_243,N_2435,N_2822);
nor UO_244 (O_244,N_2779,N_2642);
or UO_245 (O_245,N_2964,N_2832);
nand UO_246 (O_246,N_2993,N_2413);
nand UO_247 (O_247,N_2849,N_2948);
xor UO_248 (O_248,N_2819,N_2638);
and UO_249 (O_249,N_2778,N_2588);
nand UO_250 (O_250,N_2595,N_2632);
nand UO_251 (O_251,N_2538,N_2936);
and UO_252 (O_252,N_2921,N_2428);
nand UO_253 (O_253,N_2510,N_2723);
and UO_254 (O_254,N_2737,N_2429);
or UO_255 (O_255,N_2943,N_2709);
and UO_256 (O_256,N_2786,N_2929);
nand UO_257 (O_257,N_2991,N_2496);
nor UO_258 (O_258,N_2912,N_2834);
nor UO_259 (O_259,N_2482,N_2906);
or UO_260 (O_260,N_2775,N_2839);
or UO_261 (O_261,N_2442,N_2947);
or UO_262 (O_262,N_2846,N_2698);
or UO_263 (O_263,N_2439,N_2904);
nand UO_264 (O_264,N_2559,N_2547);
xor UO_265 (O_265,N_2568,N_2854);
nor UO_266 (O_266,N_2467,N_2570);
or UO_267 (O_267,N_2673,N_2759);
xnor UO_268 (O_268,N_2876,N_2791);
nand UO_269 (O_269,N_2761,N_2848);
nand UO_270 (O_270,N_2400,N_2580);
nor UO_271 (O_271,N_2480,N_2946);
xnor UO_272 (O_272,N_2764,N_2867);
xnor UO_273 (O_273,N_2818,N_2572);
and UO_274 (O_274,N_2477,N_2968);
and UO_275 (O_275,N_2581,N_2509);
nand UO_276 (O_276,N_2855,N_2402);
nor UO_277 (O_277,N_2927,N_2590);
nor UO_278 (O_278,N_2893,N_2965);
and UO_279 (O_279,N_2520,N_2498);
xnor UO_280 (O_280,N_2585,N_2563);
or UO_281 (O_281,N_2535,N_2755);
nor UO_282 (O_282,N_2748,N_2549);
nor UO_283 (O_283,N_2545,N_2795);
nand UO_284 (O_284,N_2592,N_2471);
xor UO_285 (O_285,N_2928,N_2746);
nor UO_286 (O_286,N_2573,N_2745);
xor UO_287 (O_287,N_2735,N_2694);
xnor UO_288 (O_288,N_2511,N_2850);
and UO_289 (O_289,N_2515,N_2793);
nor UO_290 (O_290,N_2449,N_2770);
nand UO_291 (O_291,N_2724,N_2643);
xor UO_292 (O_292,N_2464,N_2614);
or UO_293 (O_293,N_2905,N_2479);
nor UO_294 (O_294,N_2501,N_2978);
xnor UO_295 (O_295,N_2925,N_2857);
and UO_296 (O_296,N_2506,N_2691);
nor UO_297 (O_297,N_2591,N_2648);
nor UO_298 (O_298,N_2699,N_2765);
nand UO_299 (O_299,N_2646,N_2630);
xnor UO_300 (O_300,N_2410,N_2865);
or UO_301 (O_301,N_2756,N_2905);
xnor UO_302 (O_302,N_2722,N_2416);
and UO_303 (O_303,N_2931,N_2975);
or UO_304 (O_304,N_2919,N_2877);
xor UO_305 (O_305,N_2712,N_2478);
nor UO_306 (O_306,N_2681,N_2716);
nor UO_307 (O_307,N_2865,N_2779);
nor UO_308 (O_308,N_2560,N_2724);
xor UO_309 (O_309,N_2870,N_2499);
nand UO_310 (O_310,N_2855,N_2535);
and UO_311 (O_311,N_2655,N_2408);
nand UO_312 (O_312,N_2767,N_2668);
xor UO_313 (O_313,N_2492,N_2595);
and UO_314 (O_314,N_2587,N_2612);
nand UO_315 (O_315,N_2811,N_2407);
nor UO_316 (O_316,N_2719,N_2949);
nand UO_317 (O_317,N_2529,N_2433);
nand UO_318 (O_318,N_2420,N_2952);
nor UO_319 (O_319,N_2876,N_2589);
and UO_320 (O_320,N_2613,N_2849);
xor UO_321 (O_321,N_2979,N_2448);
nand UO_322 (O_322,N_2775,N_2776);
and UO_323 (O_323,N_2446,N_2723);
nor UO_324 (O_324,N_2501,N_2744);
xor UO_325 (O_325,N_2688,N_2899);
or UO_326 (O_326,N_2867,N_2993);
nor UO_327 (O_327,N_2971,N_2552);
nand UO_328 (O_328,N_2856,N_2655);
nor UO_329 (O_329,N_2460,N_2766);
nand UO_330 (O_330,N_2781,N_2480);
nand UO_331 (O_331,N_2785,N_2544);
and UO_332 (O_332,N_2499,N_2628);
xor UO_333 (O_333,N_2667,N_2694);
and UO_334 (O_334,N_2948,N_2800);
and UO_335 (O_335,N_2880,N_2759);
xnor UO_336 (O_336,N_2483,N_2843);
nand UO_337 (O_337,N_2427,N_2912);
nand UO_338 (O_338,N_2661,N_2732);
nor UO_339 (O_339,N_2885,N_2659);
or UO_340 (O_340,N_2534,N_2648);
and UO_341 (O_341,N_2546,N_2978);
nor UO_342 (O_342,N_2956,N_2649);
nand UO_343 (O_343,N_2969,N_2785);
nand UO_344 (O_344,N_2918,N_2785);
nor UO_345 (O_345,N_2484,N_2946);
xnor UO_346 (O_346,N_2743,N_2642);
nor UO_347 (O_347,N_2940,N_2562);
nand UO_348 (O_348,N_2972,N_2446);
and UO_349 (O_349,N_2788,N_2980);
nor UO_350 (O_350,N_2968,N_2995);
xor UO_351 (O_351,N_2536,N_2551);
nor UO_352 (O_352,N_2827,N_2698);
nor UO_353 (O_353,N_2476,N_2847);
xor UO_354 (O_354,N_2538,N_2482);
and UO_355 (O_355,N_2570,N_2545);
and UO_356 (O_356,N_2880,N_2489);
nor UO_357 (O_357,N_2762,N_2604);
or UO_358 (O_358,N_2422,N_2675);
xor UO_359 (O_359,N_2518,N_2797);
or UO_360 (O_360,N_2471,N_2527);
xor UO_361 (O_361,N_2736,N_2548);
nor UO_362 (O_362,N_2760,N_2489);
nor UO_363 (O_363,N_2623,N_2872);
nand UO_364 (O_364,N_2426,N_2611);
nor UO_365 (O_365,N_2679,N_2909);
nand UO_366 (O_366,N_2541,N_2765);
xor UO_367 (O_367,N_2907,N_2744);
xor UO_368 (O_368,N_2897,N_2999);
xor UO_369 (O_369,N_2973,N_2972);
xnor UO_370 (O_370,N_2813,N_2581);
xnor UO_371 (O_371,N_2831,N_2429);
xor UO_372 (O_372,N_2746,N_2899);
nand UO_373 (O_373,N_2929,N_2965);
nor UO_374 (O_374,N_2822,N_2447);
and UO_375 (O_375,N_2768,N_2996);
nand UO_376 (O_376,N_2478,N_2921);
and UO_377 (O_377,N_2815,N_2433);
or UO_378 (O_378,N_2647,N_2929);
and UO_379 (O_379,N_2736,N_2549);
nand UO_380 (O_380,N_2457,N_2523);
nor UO_381 (O_381,N_2810,N_2747);
or UO_382 (O_382,N_2978,N_2439);
nor UO_383 (O_383,N_2479,N_2759);
nor UO_384 (O_384,N_2495,N_2550);
nand UO_385 (O_385,N_2882,N_2877);
nor UO_386 (O_386,N_2723,N_2501);
nand UO_387 (O_387,N_2595,N_2941);
and UO_388 (O_388,N_2657,N_2949);
xor UO_389 (O_389,N_2866,N_2915);
and UO_390 (O_390,N_2589,N_2403);
nand UO_391 (O_391,N_2940,N_2457);
xor UO_392 (O_392,N_2609,N_2521);
and UO_393 (O_393,N_2442,N_2669);
xnor UO_394 (O_394,N_2825,N_2580);
xor UO_395 (O_395,N_2991,N_2721);
or UO_396 (O_396,N_2621,N_2505);
nand UO_397 (O_397,N_2659,N_2714);
nand UO_398 (O_398,N_2435,N_2685);
nor UO_399 (O_399,N_2469,N_2535);
nor UO_400 (O_400,N_2758,N_2914);
and UO_401 (O_401,N_2511,N_2891);
xor UO_402 (O_402,N_2500,N_2762);
or UO_403 (O_403,N_2698,N_2896);
or UO_404 (O_404,N_2402,N_2955);
nor UO_405 (O_405,N_2851,N_2806);
nor UO_406 (O_406,N_2661,N_2647);
xnor UO_407 (O_407,N_2752,N_2793);
nor UO_408 (O_408,N_2732,N_2829);
nor UO_409 (O_409,N_2494,N_2941);
xnor UO_410 (O_410,N_2558,N_2814);
or UO_411 (O_411,N_2714,N_2972);
nand UO_412 (O_412,N_2588,N_2965);
xor UO_413 (O_413,N_2953,N_2697);
nand UO_414 (O_414,N_2640,N_2418);
xnor UO_415 (O_415,N_2823,N_2439);
or UO_416 (O_416,N_2445,N_2408);
nor UO_417 (O_417,N_2745,N_2864);
or UO_418 (O_418,N_2644,N_2774);
nor UO_419 (O_419,N_2728,N_2850);
xnor UO_420 (O_420,N_2990,N_2672);
nor UO_421 (O_421,N_2424,N_2737);
xnor UO_422 (O_422,N_2440,N_2548);
or UO_423 (O_423,N_2635,N_2417);
and UO_424 (O_424,N_2503,N_2577);
nand UO_425 (O_425,N_2621,N_2415);
nor UO_426 (O_426,N_2684,N_2707);
nor UO_427 (O_427,N_2641,N_2961);
xnor UO_428 (O_428,N_2684,N_2681);
nand UO_429 (O_429,N_2935,N_2811);
or UO_430 (O_430,N_2676,N_2860);
nand UO_431 (O_431,N_2488,N_2772);
or UO_432 (O_432,N_2802,N_2782);
nor UO_433 (O_433,N_2637,N_2425);
nor UO_434 (O_434,N_2868,N_2808);
or UO_435 (O_435,N_2540,N_2429);
nand UO_436 (O_436,N_2701,N_2652);
and UO_437 (O_437,N_2971,N_2540);
xnor UO_438 (O_438,N_2412,N_2802);
and UO_439 (O_439,N_2770,N_2672);
nand UO_440 (O_440,N_2761,N_2552);
or UO_441 (O_441,N_2696,N_2524);
or UO_442 (O_442,N_2799,N_2818);
or UO_443 (O_443,N_2409,N_2670);
nor UO_444 (O_444,N_2908,N_2631);
xor UO_445 (O_445,N_2656,N_2497);
nand UO_446 (O_446,N_2430,N_2882);
xnor UO_447 (O_447,N_2799,N_2524);
nand UO_448 (O_448,N_2845,N_2994);
nor UO_449 (O_449,N_2680,N_2437);
or UO_450 (O_450,N_2937,N_2843);
nor UO_451 (O_451,N_2486,N_2715);
and UO_452 (O_452,N_2848,N_2638);
xor UO_453 (O_453,N_2762,N_2468);
and UO_454 (O_454,N_2920,N_2769);
nor UO_455 (O_455,N_2586,N_2769);
and UO_456 (O_456,N_2583,N_2730);
or UO_457 (O_457,N_2537,N_2430);
nor UO_458 (O_458,N_2847,N_2415);
nor UO_459 (O_459,N_2952,N_2715);
nor UO_460 (O_460,N_2530,N_2961);
nand UO_461 (O_461,N_2446,N_2601);
and UO_462 (O_462,N_2474,N_2747);
and UO_463 (O_463,N_2519,N_2781);
nor UO_464 (O_464,N_2810,N_2775);
nor UO_465 (O_465,N_2665,N_2925);
or UO_466 (O_466,N_2883,N_2783);
nor UO_467 (O_467,N_2526,N_2688);
and UO_468 (O_468,N_2948,N_2600);
and UO_469 (O_469,N_2614,N_2554);
and UO_470 (O_470,N_2435,N_2432);
or UO_471 (O_471,N_2543,N_2754);
nand UO_472 (O_472,N_2849,N_2431);
nor UO_473 (O_473,N_2861,N_2906);
nand UO_474 (O_474,N_2859,N_2402);
xnor UO_475 (O_475,N_2670,N_2845);
or UO_476 (O_476,N_2765,N_2534);
nor UO_477 (O_477,N_2421,N_2808);
and UO_478 (O_478,N_2971,N_2958);
or UO_479 (O_479,N_2912,N_2751);
xnor UO_480 (O_480,N_2831,N_2631);
nor UO_481 (O_481,N_2872,N_2856);
xnor UO_482 (O_482,N_2948,N_2871);
nand UO_483 (O_483,N_2950,N_2876);
nor UO_484 (O_484,N_2675,N_2830);
nor UO_485 (O_485,N_2489,N_2948);
and UO_486 (O_486,N_2615,N_2535);
nor UO_487 (O_487,N_2930,N_2966);
and UO_488 (O_488,N_2714,N_2860);
nand UO_489 (O_489,N_2972,N_2418);
xor UO_490 (O_490,N_2416,N_2766);
xor UO_491 (O_491,N_2549,N_2891);
and UO_492 (O_492,N_2789,N_2685);
nand UO_493 (O_493,N_2647,N_2463);
xnor UO_494 (O_494,N_2633,N_2611);
xor UO_495 (O_495,N_2583,N_2846);
nand UO_496 (O_496,N_2744,N_2608);
nand UO_497 (O_497,N_2646,N_2966);
or UO_498 (O_498,N_2881,N_2716);
or UO_499 (O_499,N_2903,N_2716);
endmodule